
module aes ( clk, rst, ld, done, \key[127] , \key[126] , \key[125] , 
        \key[124] , \key[123] , \key[122] , \key[121] , \key[120] , \key[119] , 
        \key[118] , \key[117] , \key[116] , \key[115] , \key[114] , \key[113] , 
        \key[112] , \key[111] , \key[110] , \key[109] , \key[108] , \key[107] , 
        \key[106] , \key[105] , \key[104] , \key[103] , \key[102] , \key[101] , 
        \key[100] , \key[99] , \key[98] , \key[97] , \key[96] , \key[95] , 
        \key[94] , \key[93] , \key[92] , \key[91] , \key[90] , \key[89] , 
        \key[88] , \key[87] , \key[86] , \key[85] , \key[84] , \key[83] , 
        \key[82] , \key[81] , \key[80] , \key[79] , \key[78] , \key[77] , 
        \key[76] , \key[75] , \key[74] , \key[73] , \key[72] , \key[71] , 
        \key[70] , \key[69] , \key[68] , \key[67] , \key[66] , \key[65] , 
        \key[64] , \key[63] , \key[62] , \key[61] , \key[60] , \key[59] , 
        \key[58] , \key[57] , \key[56] , \key[55] , \key[54] , \key[53] , 
        \key[52] , \key[51] , \key[50] , \key[49] , \key[48] , \key[47] , 
        \key[46] , \key[45] , \key[44] , \key[43] , \key[42] , \key[41] , 
        \key[40] , \key[39] , \key[38] , \key[37] , \key[36] , \key[35] , 
        \key[34] , \key[33] , \key[32] , \key[31] , \key[30] , \key[29] , 
        \key[28] , \key[27] , \key[26] , \key[25] , \key[24] , \key[23] , 
        \key[22] , \key[21] , \key[20] , \key[19] , \key[18] , \key[17] , 
        \key[16] , \key[15] , \key[14] , \key[13] , \key[12] , \key[11] , 
        \key[10] , \key[9] , \key[8] , \key[7] , \key[6] , \key[5] , \key[4] , 
        \key[3] , \key[2] , \key[1] , \key[0] , \text_in[127] , \text_in[126] , 
        \text_in[125] , \text_in[124] , \text_in[123] , \text_in[122] , 
        \text_in[121] , \text_in[120] , \text_in[119] , \text_in[118] , 
        \text_in[117] , \text_in[116] , \text_in[115] , \text_in[114] , 
        \text_in[113] , \text_in[112] , \text_in[111] , \text_in[110] , 
        \text_in[109] , \text_in[108] , \text_in[107] , \text_in[106] , 
        \text_in[105] , \text_in[104] , \text_in[103] , \text_in[102] , 
        \text_in[101] , \text_in[100] , \text_in[99] , \text_in[98] , 
        \text_in[97] , \text_in[96] , \text_in[95] , \text_in[94] , 
        \text_in[93] , \text_in[92] , \text_in[91] , \text_in[90] , 
        \text_in[89] , \text_in[88] , \text_in[87] , \text_in[86] , 
        \text_in[85] , \text_in[84] , \text_in[83] , \text_in[82] , 
        \text_in[81] , \text_in[80] , \text_in[79] , \text_in[78] , 
        \text_in[77] , \text_in[76] , \text_in[75] , \text_in[74] , 
        \text_in[73] , \text_in[72] , \text_in[71] , \text_in[70] , 
        \text_in[69] , \text_in[68] , \text_in[67] , \text_in[66] , 
        \text_in[65] , \text_in[64] , \text_in[63] , \text_in[62] , 
        \text_in[61] , \text_in[60] , \text_in[59] , \text_in[58] , 
        \text_in[57] , \text_in[56] , \text_in[55] , \text_in[54] , 
        \text_in[53] , \text_in[52] , \text_in[51] , \text_in[50] , 
        \text_in[49] , \text_in[48] , \text_in[47] , \text_in[46] , 
        \text_in[45] , \text_in[44] , \text_in[43] , \text_in[42] , 
        \text_in[41] , \text_in[40] , \text_in[39] , \text_in[38] , 
        \text_in[37] , \text_in[36] , \text_in[35] , \text_in[34] , 
        \text_in[33] , \text_in[32] , \text_in[31] , \text_in[30] , 
        \text_in[29] , \text_in[28] , \text_in[27] , \text_in[26] , 
        \text_in[25] , \text_in[24] , \text_in[23] , \text_in[22] , 
        \text_in[21] , \text_in[20] , \text_in[19] , \text_in[18] , 
        \text_in[17] , \text_in[16] , \text_in[15] , \text_in[14] , 
        \text_in[13] , \text_in[12] , \text_in[11] , \text_in[10] , 
        \text_in[9] , \text_in[8] , \text_in[7] , \text_in[6] , \text_in[5] , 
        \text_in[4] , \text_in[3] , \text_in[2] , \text_in[1] , \text_in[0] , 
        \text_out[127] , \text_out[126] , \text_out[125] , \text_out[124] , 
        \text_out[123] , \text_out[122] , \text_out[121] , \text_out[120] , 
        \text_out[119] , \text_out[118] , \text_out[117] , \text_out[116] , 
        \text_out[115] , \text_out[114] , \text_out[113] , \text_out[112] , 
        \text_out[111] , \text_out[110] , \text_out[109] , \text_out[108] , 
        \text_out[107] , \text_out[106] , \text_out[105] , \text_out[104] , 
        \text_out[103] , \text_out[102] , \text_out[101] , \text_out[100] , 
        \text_out[99] , \text_out[98] , \text_out[97] , \text_out[96] , 
        \text_out[95] , \text_out[94] , \text_out[93] , \text_out[92] , 
        \text_out[91] , \text_out[90] , \text_out[89] , \text_out[88] , 
        \text_out[87] , \text_out[86] , \text_out[85] , \text_out[84] , 
        \text_out[83] , \text_out[82] , \text_out[81] , \text_out[80] , 
        \text_out[79] , \text_out[78] , \text_out[77] , \text_out[76] , 
        \text_out[75] , \text_out[74] , \text_out[73] , \text_out[72] , 
        \text_out[71] , \text_out[70] , \text_out[69] , \text_out[68] , 
        \text_out[67] , \text_out[66] , \text_out[65] , \text_out[64] , 
        \text_out[63] , \text_out[62] , \text_out[61] , \text_out[60] , 
        \text_out[59] , \text_out[58] , \text_out[57] , \text_out[56] , 
        \text_out[55] , \text_out[54] , \text_out[53] , \text_out[52] , 
        \text_out[51] , \text_out[50] , \text_out[49] , \text_out[48] , 
        \text_out[47] , \text_out[46] , \text_out[45] , \text_out[44] , 
        \text_out[43] , \text_out[42] , \text_out[41] , \text_out[40] , 
        \text_out[39] , \text_out[38] , \text_out[37] , \text_out[36] , 
        \text_out[35] , \text_out[34] , \text_out[33] , \text_out[32] , 
        \text_out[31] , \text_out[30] , \text_out[29] , \text_out[28] , 
        \text_out[27] , \text_out[26] , \text_out[25] , \text_out[24] , 
        \text_out[23] , \text_out[22] , \text_out[21] , \text_out[20] , 
        \text_out[19] , \text_out[18] , \text_out[17] , \text_out[16] , 
        \text_out[15] , \text_out[14] , \text_out[13] , \text_out[12] , 
        \text_out[11] , \text_out[10] , \text_out[9] , \text_out[8] , 
        \text_out[7] , \text_out[6] , \text_out[5] , \text_out[4] , 
        \text_out[3] , \text_out[2] , \text_out[1] , \text_out[0]  );
  input clk, rst, ld, \key[127] , \key[126] , \key[125] , \key[124] ,
         \key[123] , \key[122] , \key[121] , \key[120] , \key[119] ,
         \key[118] , \key[117] , \key[116] , \key[115] , \key[114] ,
         \key[113] , \key[112] , \key[111] , \key[110] , \key[109] ,
         \key[108] , \key[107] , \key[106] , \key[105] , \key[104] ,
         \key[103] , \key[102] , \key[101] , \key[100] , \key[99] , \key[98] ,
         \key[97] , \key[96] , \key[95] , \key[94] , \key[93] , \key[92] ,
         \key[91] , \key[90] , \key[89] , \key[88] , \key[87] , \key[86] ,
         \key[85] , \key[84] , \key[83] , \key[82] , \key[81] , \key[80] ,
         \key[79] , \key[78] , \key[77] , \key[76] , \key[75] , \key[74] ,
         \key[73] , \key[72] , \key[71] , \key[70] , \key[69] , \key[68] ,
         \key[67] , \key[66] , \key[65] , \key[64] , \key[63] , \key[62] ,
         \key[61] , \key[60] , \key[59] , \key[58] , \key[57] , \key[56] ,
         \key[55] , \key[54] , \key[53] , \key[52] , \key[51] , \key[50] ,
         \key[49] , \key[48] , \key[47] , \key[46] , \key[45] , \key[44] ,
         \key[43] , \key[42] , \key[41] , \key[40] , \key[39] , \key[38] ,
         \key[37] , \key[36] , \key[35] , \key[34] , \key[33] , \key[32] ,
         \key[31] , \key[30] , \key[29] , \key[28] , \key[27] , \key[26] ,
         \key[25] , \key[24] , \key[23] , \key[22] , \key[21] , \key[20] ,
         \key[19] , \key[18] , \key[17] , \key[16] , \key[15] , \key[14] ,
         \key[13] , \key[12] , \key[11] , \key[10] , \key[9] , \key[8] ,
         \key[7] , \key[6] , \key[5] , \key[4] , \key[3] , \key[2] , \key[1] ,
         \key[0] , \text_in[127] , \text_in[126] , \text_in[125] ,
         \text_in[124] , \text_in[123] , \text_in[122] , \text_in[121] ,
         \text_in[120] , \text_in[119] , \text_in[118] , \text_in[117] ,
         \text_in[116] , \text_in[115] , \text_in[114] , \text_in[113] ,
         \text_in[112] , \text_in[111] , \text_in[110] , \text_in[109] ,
         \text_in[108] , \text_in[107] , \text_in[106] , \text_in[105] ,
         \text_in[104] , \text_in[103] , \text_in[102] , \text_in[101] ,
         \text_in[100] , \text_in[99] , \text_in[98] , \text_in[97] ,
         \text_in[96] , \text_in[95] , \text_in[94] , \text_in[93] ,
         \text_in[92] , \text_in[91] , \text_in[90] , \text_in[89] ,
         \text_in[88] , \text_in[87] , \text_in[86] , \text_in[85] ,
         \text_in[84] , \text_in[83] , \text_in[82] , \text_in[81] ,
         \text_in[80] , \text_in[79] , \text_in[78] , \text_in[77] ,
         \text_in[76] , \text_in[75] , \text_in[74] , \text_in[73] ,
         \text_in[72] , \text_in[71] , \text_in[70] , \text_in[69] ,
         \text_in[68] , \text_in[67] , \text_in[66] , \text_in[65] ,
         \text_in[64] , \text_in[63] , \text_in[62] , \text_in[61] ,
         \text_in[60] , \text_in[59] , \text_in[58] , \text_in[57] ,
         \text_in[56] , \text_in[55] , \text_in[54] , \text_in[53] ,
         \text_in[52] , \text_in[51] , \text_in[50] , \text_in[49] ,
         \text_in[48] , \text_in[47] , \text_in[46] , \text_in[45] ,
         \text_in[44] , \text_in[43] , \text_in[42] , \text_in[41] ,
         \text_in[40] , \text_in[39] , \text_in[38] , \text_in[37] ,
         \text_in[36] , \text_in[35] , \text_in[34] , \text_in[33] ,
         \text_in[32] , \text_in[31] , \text_in[30] , \text_in[29] ,
         \text_in[28] , \text_in[27] , \text_in[26] , \text_in[25] ,
         \text_in[24] , \text_in[23] , \text_in[22] , \text_in[21] ,
         \text_in[20] , \text_in[19] , \text_in[18] , \text_in[17] ,
         \text_in[16] , \text_in[15] , \text_in[14] , \text_in[13] ,
         \text_in[12] , \text_in[11] , \text_in[10] , \text_in[9] ,
         \text_in[8] , \text_in[7] , \text_in[6] , \text_in[5] , \text_in[4] ,
         \text_in[3] , \text_in[2] , \text_in[1] , \text_in[0] ;
  output done, \text_out[127] , \text_out[126] , \text_out[125] ,
         \text_out[124] , \text_out[123] , \text_out[122] , \text_out[121] ,
         \text_out[120] , \text_out[119] , \text_out[118] , \text_out[117] ,
         \text_out[116] , \text_out[115] , \text_out[114] , \text_out[113] ,
         \text_out[112] , \text_out[111] , \text_out[110] , \text_out[109] ,
         \text_out[108] , \text_out[107] , \text_out[106] , \text_out[105] ,
         \text_out[104] , \text_out[103] , \text_out[102] , \text_out[101] ,
         \text_out[100] , \text_out[99] , \text_out[98] , \text_out[97] ,
         \text_out[96] , \text_out[95] , \text_out[94] , \text_out[93] ,
         \text_out[92] , \text_out[91] , \text_out[90] , \text_out[89] ,
         \text_out[88] , \text_out[87] , \text_out[86] , \text_out[85] ,
         \text_out[84] , \text_out[83] , \text_out[82] , \text_out[81] ,
         \text_out[80] , \text_out[79] , \text_out[78] , \text_out[77] ,
         \text_out[76] , \text_out[75] , \text_out[74] , \text_out[73] ,
         \text_out[72] , \text_out[71] , \text_out[70] , \text_out[69] ,
         \text_out[68] , \text_out[67] , \text_out[66] , \text_out[65] ,
         \text_out[64] , \text_out[63] , \text_out[62] , \text_out[61] ,
         \text_out[60] , \text_out[59] , \text_out[58] , \text_out[57] ,
         \text_out[56] , \text_out[55] , \text_out[54] , \text_out[53] ,
         \text_out[52] , \text_out[51] , \text_out[50] , \text_out[49] ,
         \text_out[48] , \text_out[47] , \text_out[46] , \text_out[45] ,
         \text_out[44] , \text_out[43] , \text_out[42] , \text_out[41] ,
         \text_out[40] , \text_out[39] , \text_out[38] , \text_out[37] ,
         \text_out[36] , \text_out[35] , \text_out[34] , \text_out[33] ,
         \text_out[32] , \text_out[31] , \text_out[30] , \text_out[29] ,
         \text_out[28] , \text_out[27] , \text_out[26] , \text_out[25] ,
         \text_out[24] , \text_out[23] , \text_out[22] , \text_out[21] ,
         \text_out[20] , \text_out[19] , \text_out[18] , \text_out[17] ,
         \text_out[16] , \text_out[15] , \text_out[14] , \text_out[13] ,
         \text_out[12] , \text_out[11] , \text_out[10] , \text_out[9] ,
         \text_out[8] , \text_out[7] , \text_out[6] , \text_out[5] ,
         \text_out[4] , \text_out[3] , \text_out[2] , \text_out[1] ,
         \text_out[0] ;
  wire   N23, N34, N35, N36, N37, N38, N39, N40, N41, N50, N51, N52, N53, N54,
         N55, N56, N57, N66, N67, N68, N69, N70, N71, N72, N73, N82, N83, N84,
         N85, N86, N87, N88, N89, N98, N99, N100, N101, N102, N103, N104, N105,
         N114, N115, N116, N117, N118, N119, N120, N121, N130, N131, N132,
         N133, N134, N135, N136, N137, N146, N147, N148, N149, N150, N151,
         N152, N153, N162, N163, N164, N165, N166, N167, N168, N169, N178,
         N179, N180, N181, N182, N183, N184, N185, N194, N195, N196, N197,
         N198, N199, N200, N201, N210, N211, N212, N213, N214, N215, N216,
         N217, N226, N227, N228, N229, N230, N231, N232, N233, N242, N243,
         N244, N245, N246, N247, N248, N249, N258, N259, N260, N261, N262,
         N263, N264, N265, N274, N275, N276, N277, N278, N279, N280, N281,
         N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410,
         N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421,
         N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443,
         N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465,
         N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476,
         N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487,
         N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498,
         N499, N500, N501, N502, N503, N504, N505, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1351, n1352, n1353, n1354, \u0/N271 ,
         \u0/N270 , \u0/N269 , \u0/N268 , \u0/N267 , \u0/N266 , \u0/N265 ,
         \u0/N264 , \u0/N263 , \u0/N262 , \u0/N261 , \u0/N260 , \u0/N259 ,
         \u0/N258 , \u0/N257 , \u0/N256 , \u0/N255 , \u0/N254 , \u0/N253 ,
         \u0/N252 , \u0/N251 , \u0/N250 , \u0/N249 , \u0/N248 , \u0/N247 ,
         \u0/N246 , \u0/N245 , \u0/N244 , \u0/N243 , \u0/N242 , \u0/N241 ,
         \u0/N240 , \u0/N205 , \u0/N204 , \u0/N203 , \u0/N202 , \u0/N201 ,
         \u0/N200 , \u0/N199 , \u0/N198 , \u0/N197 , \u0/N196 , \u0/N195 ,
         \u0/N194 , \u0/N193 , \u0/N192 , \u0/N191 , \u0/N190 , \u0/N189 ,
         \u0/N188 , \u0/N187 , \u0/N186 , \u0/N185 , \u0/N184 , \u0/N183 ,
         \u0/N182 , \u0/N181 , \u0/N180 , \u0/N179 , \u0/N178 , \u0/N177 ,
         \u0/N176 , \u0/N175 , \u0/N174 , \u0/N139 , \u0/N138 , \u0/N137 ,
         \u0/N136 , \u0/N135 , \u0/N134 , \u0/N133 , \u0/N132 , \u0/N131 ,
         \u0/N130 , \u0/N129 , \u0/N128 , \u0/N127 , \u0/N126 , \u0/N125 ,
         \u0/N124 , \u0/N123 , \u0/N122 , \u0/N121 , \u0/N120 , \u0/N119 ,
         \u0/N118 , \u0/N117 , \u0/N116 , \u0/N115 , \u0/N114 , \u0/N113 ,
         \u0/N112 , \u0/N111 , \u0/N110 , \u0/N109 , \u0/N108 , \u0/N73 ,
         \u0/N72 , \u0/N71 , \u0/N70 , \u0/N69 , \u0/N68 , \u0/N67 , \u0/N66 ,
         \u0/N65 , \u0/N64 , \u0/N63 , \u0/N62 , \u0/N61 , \u0/N60 , \u0/N59 ,
         \u0/N58 , \u0/N57 , \u0/N56 , \u0/N55 , \u0/N54 , \u0/N53 , \u0/N52 ,
         \u0/N51 , \u0/N50 , \u0/N49 , \u0/N48 , \u0/N47 , \u0/N46 , \u0/N45 ,
         \u0/N44 , \u0/N43 , \u0/N42 , \u0/r0/n3 , \u0/r0/N81 , \u0/r0/N80 ,
         \u0/r0/N79 , \u0/r0/N78 , \u0/r0/N77 , \u0/r0/N76 , \u0/r0/N75 ,
         \u0/r0/N74 , \u0/r0/N73 , \u0/r0/N72 , \u0/r0/N71 , \u0/r0/N70 ,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588;


  dffs1 \dcnt_reg[0]  ( .DIN(n1354), .CLK(clk), .Q(n15579), .QN(n1449) );
  dffs1 \dcnt_reg[1]  ( .DIN(n1352), .CLK(clk), .Q(n15577), .QN(n1409) );
  dffs1 \dcnt_reg[3]  ( .DIN(n1353), .CLK(clk), .Q(n15578), .QN(n1526) );
  dffs1 \dcnt_reg[2]  ( .DIN(n1351), .CLK(clk), .QN(n1360) );
  dffs1 done_reg ( .DIN(N23), .CLK(clk), .Q(done) );
  dffs1 \text_in_r_reg[127]  ( .DIN(n1346), .CLK(clk), .Q(text_in_r[127]) );
  dffs1 \text_in_r_reg[126]  ( .DIN(n1345), .CLK(clk), .Q(text_in_r[126]) );
  dffs1 \text_in_r_reg[125]  ( .DIN(n1344), .CLK(clk), .Q(text_in_r[125]) );
  dffs1 \text_in_r_reg[124]  ( .DIN(n1343), .CLK(clk), .Q(text_in_r[124]) );
  dffs1 \text_in_r_reg[123]  ( .DIN(n1342), .CLK(clk), .Q(text_in_r[123]) );
  dffs1 \text_in_r_reg[122]  ( .DIN(n1341), .CLK(clk), .Q(text_in_r[122]) );
  dffs1 \text_in_r_reg[121]  ( .DIN(n1340), .CLK(clk), .Q(text_in_r[121]) );
  dffs1 \text_in_r_reg[120]  ( .DIN(n1339), .CLK(clk), .Q(text_in_r[120]) );
  dffs1 \text_in_r_reg[119]  ( .DIN(n1338), .CLK(clk), .Q(text_in_r[119]) );
  dffs1 \text_in_r_reg[118]  ( .DIN(n1337), .CLK(clk), .Q(text_in_r[118]) );
  dffs1 \text_in_r_reg[117]  ( .DIN(n1336), .CLK(clk), .Q(text_in_r[117]) );
  dffs1 \text_in_r_reg[116]  ( .DIN(n1335), .CLK(clk), .Q(text_in_r[116]) );
  dffs1 \text_in_r_reg[115]  ( .DIN(n1334), .CLK(clk), .Q(text_in_r[115]) );
  dffs1 \text_in_r_reg[114]  ( .DIN(n1333), .CLK(clk), .Q(text_in_r[114]) );
  dffs1 \text_in_r_reg[113]  ( .DIN(n1332), .CLK(clk), .Q(text_in_r[113]) );
  dffs1 \text_in_r_reg[112]  ( .DIN(n1331), .CLK(clk), .Q(text_in_r[112]) );
  dffs1 \text_in_r_reg[111]  ( .DIN(n1330), .CLK(clk), .Q(text_in_r[111]) );
  dffs1 \text_in_r_reg[110]  ( .DIN(n1329), .CLK(clk), .Q(text_in_r[110]) );
  dffs1 \text_in_r_reg[109]  ( .DIN(n1328), .CLK(clk), .Q(text_in_r[109]) );
  dffs1 \text_in_r_reg[108]  ( .DIN(n1327), .CLK(clk), .Q(text_in_r[108]) );
  dffs1 \text_in_r_reg[107]  ( .DIN(n1326), .CLK(clk), .Q(text_in_r[107]) );
  dffs1 \text_in_r_reg[106]  ( .DIN(n1325), .CLK(clk), .Q(text_in_r[106]) );
  dffs1 \text_in_r_reg[105]  ( .DIN(n1324), .CLK(clk), .Q(text_in_r[105]) );
  dffs1 \text_in_r_reg[104]  ( .DIN(n1323), .CLK(clk), .Q(text_in_r[104]) );
  dffs1 \text_in_r_reg[103]  ( .DIN(n1322), .CLK(clk), .Q(text_in_r[103]) );
  dffs1 \text_in_r_reg[102]  ( .DIN(n1321), .CLK(clk), .Q(text_in_r[102]) );
  dffs1 \text_in_r_reg[101]  ( .DIN(n1320), .CLK(clk), .Q(text_in_r[101]) );
  dffs1 \text_in_r_reg[100]  ( .DIN(n1319), .CLK(clk), .Q(text_in_r[100]) );
  dffs1 \text_in_r_reg[99]  ( .DIN(n1318), .CLK(clk), .Q(text_in_r[99]) );
  dffs1 \text_in_r_reg[98]  ( .DIN(n1317), .CLK(clk), .Q(text_in_r[98]) );
  dffs1 \text_in_r_reg[97]  ( .DIN(n1316), .CLK(clk), .Q(text_in_r[97]) );
  dffs1 \text_in_r_reg[96]  ( .DIN(n1315), .CLK(clk), .Q(text_in_r[96]) );
  dffs1 \text_in_r_reg[95]  ( .DIN(n1314), .CLK(clk), .Q(text_in_r[95]) );
  dffs1 \text_in_r_reg[94]  ( .DIN(n1313), .CLK(clk), .Q(text_in_r[94]) );
  dffs1 \text_in_r_reg[93]  ( .DIN(n1312), .CLK(clk), .Q(text_in_r[93]) );
  dffs1 \text_in_r_reg[92]  ( .DIN(n1311), .CLK(clk), .Q(text_in_r[92]) );
  dffs1 \text_in_r_reg[91]  ( .DIN(n1310), .CLK(clk), .Q(text_in_r[91]) );
  dffs1 \text_in_r_reg[90]  ( .DIN(n1309), .CLK(clk), .Q(text_in_r[90]) );
  dffs1 \text_in_r_reg[89]  ( .DIN(n1308), .CLK(clk), .Q(text_in_r[89]) );
  dffs1 \text_in_r_reg[88]  ( .DIN(n1307), .CLK(clk), .Q(text_in_r[88]) );
  dffs1 \text_in_r_reg[87]  ( .DIN(n1306), .CLK(clk), .Q(text_in_r[87]) );
  dffs1 \text_in_r_reg[86]  ( .DIN(n1305), .CLK(clk), .Q(text_in_r[86]) );
  dffs1 \text_in_r_reg[85]  ( .DIN(n1304), .CLK(clk), .Q(text_in_r[85]) );
  dffs1 \text_in_r_reg[84]  ( .DIN(n1303), .CLK(clk), .Q(text_in_r[84]) );
  dffs1 \text_in_r_reg[83]  ( .DIN(n1302), .CLK(clk), .Q(text_in_r[83]) );
  dffs1 \text_in_r_reg[82]  ( .DIN(n1301), .CLK(clk), .Q(text_in_r[82]) );
  dffs1 \text_in_r_reg[81]  ( .DIN(n1300), .CLK(clk), .Q(text_in_r[81]) );
  dffs1 \text_in_r_reg[80]  ( .DIN(n1299), .CLK(clk), .Q(text_in_r[80]) );
  dffs1 \text_in_r_reg[79]  ( .DIN(n1298), .CLK(clk), .Q(text_in_r[79]) );
  dffs1 \text_in_r_reg[78]  ( .DIN(n1297), .CLK(clk), .Q(text_in_r[78]) );
  dffs1 \text_in_r_reg[77]  ( .DIN(n1296), .CLK(clk), .Q(text_in_r[77]) );
  dffs1 \text_in_r_reg[76]  ( .DIN(n1295), .CLK(clk), .Q(text_in_r[76]) );
  dffs1 \text_in_r_reg[75]  ( .DIN(n1294), .CLK(clk), .Q(text_in_r[75]) );
  dffs1 \text_in_r_reg[74]  ( .DIN(n1293), .CLK(clk), .Q(text_in_r[74]) );
  dffs1 \text_in_r_reg[73]  ( .DIN(n1292), .CLK(clk), .Q(text_in_r[73]) );
  dffs1 \text_in_r_reg[72]  ( .DIN(n1291), .CLK(clk), .Q(text_in_r[72]) );
  dffs1 \text_in_r_reg[71]  ( .DIN(n1290), .CLK(clk), .Q(text_in_r[71]) );
  dffs1 \text_in_r_reg[70]  ( .DIN(n1289), .CLK(clk), .Q(text_in_r[70]) );
  dffs1 \text_in_r_reg[69]  ( .DIN(n1288), .CLK(clk), .Q(text_in_r[69]) );
  dffs1 \text_in_r_reg[68]  ( .DIN(n1287), .CLK(clk), .Q(text_in_r[68]) );
  dffs1 \text_in_r_reg[67]  ( .DIN(n1286), .CLK(clk), .Q(text_in_r[67]) );
  dffs1 \text_in_r_reg[66]  ( .DIN(n1285), .CLK(clk), .Q(text_in_r[66]) );
  dffs1 \text_in_r_reg[65]  ( .DIN(n1284), .CLK(clk), .Q(text_in_r[65]) );
  dffs1 \text_in_r_reg[64]  ( .DIN(n1283), .CLK(clk), .Q(text_in_r[64]) );
  dffs1 \text_in_r_reg[63]  ( .DIN(n1282), .CLK(clk), .Q(text_in_r[63]) );
  dffs1 \text_in_r_reg[62]  ( .DIN(n1281), .CLK(clk), .Q(text_in_r[62]) );
  dffs1 \text_in_r_reg[61]  ( .DIN(n1280), .CLK(clk), .Q(text_in_r[61]) );
  dffs1 \text_in_r_reg[60]  ( .DIN(n1279), .CLK(clk), .Q(text_in_r[60]) );
  dffs1 \text_in_r_reg[59]  ( .DIN(n1278), .CLK(clk), .Q(text_in_r[59]) );
  dffs1 \text_in_r_reg[58]  ( .DIN(n1277), .CLK(clk), .Q(text_in_r[58]) );
  dffs1 \text_in_r_reg[57]  ( .DIN(n1276), .CLK(clk), .Q(text_in_r[57]) );
  dffs1 \text_in_r_reg[56]  ( .DIN(n1275), .CLK(clk), .Q(text_in_r[56]) );
  dffs1 \text_in_r_reg[55]  ( .DIN(n1274), .CLK(clk), .Q(text_in_r[55]) );
  dffs1 \text_in_r_reg[54]  ( .DIN(n1273), .CLK(clk), .Q(text_in_r[54]) );
  dffs1 \text_in_r_reg[53]  ( .DIN(n1272), .CLK(clk), .Q(text_in_r[53]) );
  dffs1 \text_in_r_reg[52]  ( .DIN(n1271), .CLK(clk), .Q(text_in_r[52]) );
  dffs1 \text_in_r_reg[51]  ( .DIN(n1270), .CLK(clk), .Q(text_in_r[51]) );
  dffs1 \text_in_r_reg[50]  ( .DIN(n1269), .CLK(clk), .Q(text_in_r[50]) );
  dffs1 \text_in_r_reg[49]  ( .DIN(n1268), .CLK(clk), .Q(text_in_r[49]) );
  dffs1 \text_in_r_reg[48]  ( .DIN(n1267), .CLK(clk), .Q(text_in_r[48]) );
  dffs1 \text_in_r_reg[47]  ( .DIN(n1266), .CLK(clk), .Q(text_in_r[47]) );
  dffs1 \text_in_r_reg[46]  ( .DIN(n1265), .CLK(clk), .Q(text_in_r[46]) );
  dffs1 \text_in_r_reg[45]  ( .DIN(n1264), .CLK(clk), .Q(text_in_r[45]) );
  dffs1 \text_in_r_reg[44]  ( .DIN(n1263), .CLK(clk), .Q(text_in_r[44]) );
  dffs1 \text_in_r_reg[43]  ( .DIN(n1262), .CLK(clk), .Q(text_in_r[43]) );
  dffs1 \text_in_r_reg[42]  ( .DIN(n1261), .CLK(clk), .Q(text_in_r[42]) );
  dffs1 \text_in_r_reg[41]  ( .DIN(n1260), .CLK(clk), .Q(text_in_r[41]) );
  dffs1 \text_in_r_reg[40]  ( .DIN(n1259), .CLK(clk), .Q(text_in_r[40]) );
  dffs1 \text_in_r_reg[39]  ( .DIN(n1258), .CLK(clk), .Q(text_in_r[39]) );
  dffs1 \text_in_r_reg[38]  ( .DIN(n1257), .CLK(clk), .Q(text_in_r[38]) );
  dffs1 \text_in_r_reg[37]  ( .DIN(n1256), .CLK(clk), .Q(text_in_r[37]) );
  dffs1 \text_in_r_reg[36]  ( .DIN(n1255), .CLK(clk), .Q(text_in_r[36]) );
  dffs1 \text_in_r_reg[35]  ( .DIN(n1254), .CLK(clk), .Q(text_in_r[35]) );
  dffs1 \text_in_r_reg[34]  ( .DIN(n1253), .CLK(clk), .Q(text_in_r[34]) );
  dffs1 \text_in_r_reg[33]  ( .DIN(n1252), .CLK(clk), .Q(text_in_r[33]) );
  dffs1 \text_in_r_reg[32]  ( .DIN(n1251), .CLK(clk), .Q(text_in_r[32]) );
  dffs1 \text_in_r_reg[31]  ( .DIN(n1250), .CLK(clk), .Q(text_in_r[31]) );
  dffs1 \text_in_r_reg[30]  ( .DIN(n1249), .CLK(clk), .Q(text_in_r[30]) );
  dffs1 \text_in_r_reg[29]  ( .DIN(n1248), .CLK(clk), .Q(text_in_r[29]) );
  dffs1 \text_in_r_reg[28]  ( .DIN(n1247), .CLK(clk), .Q(text_in_r[28]) );
  dffs1 \text_in_r_reg[27]  ( .DIN(n1246), .CLK(clk), .Q(text_in_r[27]) );
  dffs1 \text_in_r_reg[26]  ( .DIN(n1245), .CLK(clk), .Q(text_in_r[26]) );
  dffs1 \text_in_r_reg[25]  ( .DIN(n1244), .CLK(clk), .Q(text_in_r[25]) );
  dffs1 \text_in_r_reg[24]  ( .DIN(n1243), .CLK(clk), .Q(text_in_r[24]) );
  dffs1 \text_in_r_reg[23]  ( .DIN(n1242), .CLK(clk), .Q(text_in_r[23]) );
  dffs1 \text_in_r_reg[22]  ( .DIN(n1241), .CLK(clk), .Q(text_in_r[22]) );
  dffs1 \text_in_r_reg[21]  ( .DIN(n1240), .CLK(clk), .Q(text_in_r[21]) );
  dffs1 \text_in_r_reg[20]  ( .DIN(n1239), .CLK(clk), .Q(text_in_r[20]) );
  dffs1 \text_in_r_reg[19]  ( .DIN(n1238), .CLK(clk), .Q(text_in_r[19]) );
  dffs1 \text_in_r_reg[18]  ( .DIN(n1237), .CLK(clk), .Q(text_in_r[18]) );
  dffs1 \text_in_r_reg[17]  ( .DIN(n1236), .CLK(clk), .Q(text_in_r[17]) );
  dffs1 \text_in_r_reg[16]  ( .DIN(n1235), .CLK(clk), .Q(text_in_r[16]) );
  dffs1 \text_in_r_reg[15]  ( .DIN(n1234), .CLK(clk), .Q(text_in_r[15]) );
  dffs1 \text_in_r_reg[14]  ( .DIN(n1233), .CLK(clk), .Q(text_in_r[14]) );
  dffs1 \text_in_r_reg[13]  ( .DIN(n1232), .CLK(clk), .Q(text_in_r[13]) );
  dffs1 \text_in_r_reg[12]  ( .DIN(n1231), .CLK(clk), .Q(text_in_r[12]) );
  dffs1 \text_in_r_reg[11]  ( .DIN(n1230), .CLK(clk), .Q(text_in_r[11]) );
  dffs1 \text_in_r_reg[10]  ( .DIN(n1229), .CLK(clk), .Q(text_in_r[10]) );
  dffs1 \text_in_r_reg[9]  ( .DIN(n1228), .CLK(clk), .Q(text_in_r[9]) );
  dffs1 \text_in_r_reg[8]  ( .DIN(n1227), .CLK(clk), .Q(text_in_r[8]) );
  dffs1 \text_in_r_reg[7]  ( .DIN(n1226), .CLK(clk), .Q(text_in_r[7]) );
  dffs1 \text_in_r_reg[6]  ( .DIN(n1225), .CLK(clk), .Q(text_in_r[6]) );
  dffs1 \text_in_r_reg[5]  ( .DIN(n1224), .CLK(clk), .Q(text_in_r[5]) );
  dffs1 \text_in_r_reg[4]  ( .DIN(n1223), .CLK(clk), .Q(text_in_r[4]) );
  dffs1 \text_in_r_reg[3]  ( .DIN(n1222), .CLK(clk), .Q(text_in_r[3]) );
  dffs1 \text_in_r_reg[2]  ( .DIN(n1221), .CLK(clk), .Q(text_in_r[2]) );
  dffs1 \text_in_r_reg[1]  ( .DIN(n1220), .CLK(clk), .Q(text_in_r[1]) );
  dffs1 \text_in_r_reg[0]  ( .DIN(n1219), .CLK(clk), .Q(text_in_r[0]) );
  dffs1 ld_r_reg ( .DIN(ld), .CLK(clk), .Q(n15580), .QN(n1543) );
  dffs1 \sa00_reg[0]  ( .DIN(N274), .CLK(clk), .Q(sa00[0]), .QN(n1363) );
  dffs1 \sa10_reg[7]  ( .DIN(N265), .CLK(clk), .Q(sa10[7]), .QN(n1516) );
  dffs1 \sa03_reg[7]  ( .DIN(N89), .CLK(clk), .Q(sa03[7]), .QN(n1515) );
  dffs1 \sa13_reg[7]  ( .DIN(N73), .CLK(clk), .Q(sa13[7]), .QN(n1422) );
  dffs1 \sa02_reg[7]  ( .DIN(N153), .CLK(clk), .Q(sa02[7]), .QN(n1524) );
  dffs1 \sa12_reg[7]  ( .DIN(N137), .CLK(clk), .Q(sa12[7]), .QN(n1521) );
  dffs1 \sa01_reg[7]  ( .DIN(N217), .CLK(clk), .Q(sa01[7]), .QN(n1522) );
  dffs1 \sa11_reg[7]  ( .DIN(N201), .CLK(clk), .Q(sa11[7]), .QN(n1518) );
  dffs1 \sa30_reg[7]  ( .DIN(N233), .CLK(clk), .Q(sa30[7]) );
  dffs1 \sa21_reg[7]  ( .DIN(N185), .CLK(clk), .Q(sa21[7]), .QN(n1517) );
  dffs1 \sa23_reg[0]  ( .DIN(N50), .CLK(clk), .Q(sa23[0]), .QN(n1367) );
  dffs1 \sa31_reg[0]  ( .DIN(N162), .CLK(clk), .Q(sa31[0]), .QN(n1379) );
  dffs1 \sa01_reg[0]  ( .DIN(N210), .CLK(clk), .Q(sa01[0]), .QN(n1366) );
  dffs1 \sa31_reg[1]  ( .DIN(N163), .CLK(clk), .Q(sa31[1]), .QN(n1421) );
  dffs1 \sa01_reg[1]  ( .DIN(N211), .CLK(clk), .Q(sa01[1]), .QN(n1434) );
  dffs1 \sa21_reg[2]  ( .DIN(N180), .CLK(clk), .Q(sa21[2]), .QN(n1390) );
  dffs1 \sa31_reg[2]  ( .DIN(N164), .CLK(clk), .Q(sa31[2]), .QN(n1418) );
  dffs1 \sa01_reg[2]  ( .DIN(N212), .CLK(clk), .Q(sa01[2]), .QN(n1447) );
  dffs1 \sa11_reg[2]  ( .DIN(N196), .CLK(clk), .Q(sa11[2]), .QN(n1443) );
  dffs1 \sa31_reg[3]  ( .DIN(N165), .CLK(clk), .Q(sa31[3]), .QN(n1378) );
  dffs1 \sa01_reg[3]  ( .DIN(N213), .CLK(clk), .Q(sa01[3]) );
  dffs1 \sa31_reg[4]  ( .DIN(N166), .CLK(clk), .Q(sa31[4]), .QN(n1511) );
  dffs1 \sa01_reg[4]  ( .DIN(N214), .CLK(clk), .Q(sa01[4]), .QN(n1535) );
  dffs1 \sa21_reg[5]  ( .DIN(N183), .CLK(clk), .Q(sa21[5]), .QN(n1399) );
  dffs1 \sa31_reg[5]  ( .DIN(N167), .CLK(clk), .Q(sa31[5]), .QN(n1408) );
  dffs1 \sa01_reg[5]  ( .DIN(N215), .CLK(clk), .Q(sa01[5]), .QN(n1404) );
  dffs1 \sa11_reg[5]  ( .DIN(N199), .CLK(clk), .Q(sa11[5]), .QN(n1400) );
  dffs1 \sa21_reg[6]  ( .DIN(N184), .CLK(clk), .Q(sa21[6]) );
  dffs1 \sa31_reg[6]  ( .DIN(N168), .CLK(clk), .Q(sa31[6]) );
  dffs1 \sa01_reg[6]  ( .DIN(N216), .CLK(clk), .Q(sa01[6]) );
  dffs1 \sa11_reg[6]  ( .DIN(N200), .CLK(clk), .Q(sa11[6]) );
  dffs1 \sa31_reg[7]  ( .DIN(N169), .CLK(clk), .Q(sa31[7]), .QN(n1539) );
  dffs1 \sa22_reg[7]  ( .DIN(N121), .CLK(clk), .Q(sa22[7]), .QN(n1520) );
  dffs1 \sa20_reg[0]  ( .DIN(N242), .CLK(clk), .Q(sa20[0]), .QN(n1359) );
  dffs1 \sa02_reg[0]  ( .DIN(N146), .CLK(clk), .Q(sa02[0]), .QN(n1380) );
  dffs1 \sa32_reg[0]  ( .DIN(N98), .CLK(clk), .Q(sa32[0]), .QN(n1395) );
  dffs1 \sa02_reg[1]  ( .DIN(N147), .CLK(clk), .Q(sa02[1]), .QN(n1420) );
  dffs1 \sa22_reg[2]  ( .DIN(N116), .CLK(clk), .Q(sa22[2]), .QN(n1445) );
  dffs1 \sa32_reg[1]  ( .DIN(N99), .CLK(clk), .Q(sa32[1]), .QN(n1394) );
  dffs1 \sa32_reg[2]  ( .DIN(N100), .CLK(clk), .Q(sa32[2]), .QN(n1513) );
  dffs1 \sa02_reg[2]  ( .DIN(N148), .CLK(clk), .Q(sa02[2]), .QN(n1417) );
  dffs1 \sa12_reg[2]  ( .DIN(N132), .CLK(clk), .Q(sa12[2]), .QN(n1446) );
  dffs1 \sa32_reg[3]  ( .DIN(N101), .CLK(clk), .Q(sa32[3]), .QN(n1512) );
  dffs1 \sa02_reg[3]  ( .DIN(N149), .CLK(clk), .Q(sa02[3]), .QN(n1377) );
  dffs1 \sa32_reg[4]  ( .DIN(N102), .CLK(clk), .Q(sa32[4]) );
  dffs1 \sa02_reg[4]  ( .DIN(N150), .CLK(clk), .Q(sa02[4]), .QN(n1406) );
  dffs1 \sa22_reg[5]  ( .DIN(N119), .CLK(clk), .Q(sa22[5]), .QN(n1402) );
  dffs1 \sa32_reg[5]  ( .DIN(N103), .CLK(clk), .Q(sa32[5]), .QN(n1381) );
  dffs1 \sa02_reg[5]  ( .DIN(N151), .CLK(clk), .Q(sa02[5]), .QN(n1525) );
  dffs1 \sa12_reg[5]  ( .DIN(N135), .CLK(clk), .Q(sa12[5]), .QN(n1403) );
  dffs1 \sa22_reg[6]  ( .DIN(N120), .CLK(clk), .Q(sa22[6]) );
  dffs1 \sa32_reg[6]  ( .DIN(N104), .CLK(clk), .Q(sa32[6]), .QN(n1425) );
  dffs1 \sa02_reg[6]  ( .DIN(N152), .CLK(clk), .Q(sa02[6]), .QN(n1407) );
  dffs1 \sa12_reg[6]  ( .DIN(N136), .CLK(clk), .Q(sa12[6]) );
  dffs1 \sa32_reg[7]  ( .DIN(N105), .CLK(clk), .Q(sa32[7]) );
  dffs1 \sa03_reg[0]  ( .DIN(N82), .CLK(clk), .Q(sa03[0]), .QN(n1355) );
  dffs1 \sa33_reg[2]  ( .DIN(N36), .CLK(clk), .Q(sa33[2]), .QN(n1537) );
  dffs1 \sa23_reg[1]  ( .DIN(N51), .CLK(clk), .Q(sa23[1]), .QN(n1435) );
  dffs1 \sa03_reg[1]  ( .DIN(N83), .CLK(clk), .Q(sa03[1]), .QN(n1424) );
  dffs1 \sa23_reg[2]  ( .DIN(N52), .CLK(clk), .Q(sa23[2]), .QN(n1448) );
  dffs1 \sa03_reg[2]  ( .DIN(N84), .CLK(clk), .Q(sa03[2]), .QN(n1388) );
  dffs1 \sa13_reg[2]  ( .DIN(N68), .CLK(clk), .Q(sa13[2]), .QN(n1386) );
  dffs1 \sa23_reg[3]  ( .DIN(N53), .CLK(clk), .Q(sa23[3]) );
  dffs1 \sa03_reg[3]  ( .DIN(N85), .CLK(clk), .Q(sa03[3]), .QN(n1508) );
  dffs1 \sa33_reg[5]  ( .DIN(N39), .CLK(clk), .Q(sa33[5]), .QN(n1382) );
  dffs1 \sa23_reg[4]  ( .DIN(N54), .CLK(clk), .Q(sa23[4]), .QN(n1536) );
  dffs1 \sa03_reg[4]  ( .DIN(N86), .CLK(clk), .Q(sa03[4]), .QN(n1396) );
  dffs1 \sa33_reg[6]  ( .DIN(N40), .CLK(clk), .Q(sa33[6]), .QN(n1428) );
  dffs1 \sa23_reg[5]  ( .DIN(N55), .CLK(clk), .Q(sa23[5]), .QN(n1405) );
  dffs1 \sa03_reg[5]  ( .DIN(N87), .CLK(clk), .Q(sa03[5]), .QN(n1397) );
  dffs1 \sa13_reg[5]  ( .DIN(N71), .CLK(clk), .Q(sa13[5]), .QN(n1384) );
  dffs1 \sa33_reg[7]  ( .DIN(N41), .CLK(clk), .Q(sa33[7]) );
  dffs1 \sa23_reg[6]  ( .DIN(N56), .CLK(clk), .Q(sa23[6]) );
  dffs1 \sa03_reg[6]  ( .DIN(N88), .CLK(clk), .Q(sa03[6]), .QN(n1514) );
  dffs1 \sa13_reg[6]  ( .DIN(N72), .CLK(clk), .QN(n1370) );
  dffs1 \sa33_reg[4]  ( .DIN(N38), .CLK(clk), .Q(sa33[4]) );
  dffs1 \sa33_reg[3]  ( .DIN(N37), .CLK(clk), .Q(sa33[3]) );
  dffs1 \sa33_reg[1]  ( .DIN(N35), .CLK(clk), .Q(sa33[1]), .QN(n1529) );
  dffs1 \sa33_reg[0]  ( .DIN(N34), .CLK(clk), .Q(sa33[0]) );
  dffs1 \sa30_reg[2]  ( .DIN(N228), .CLK(clk), .Q(sa30[2]), .QN(n1538) );
  dffs1 \sa20_reg[1]  ( .DIN(N243), .CLK(clk), .Q(sa20[1]), .QN(n1507) );
  dffs1 \sa00_reg[1]  ( .DIN(N275), .CLK(clk), .Q(sa00[1]), .QN(n1430) );
  dffs1 \sa20_reg[2]  ( .DIN(N244), .CLK(clk), .Q(sa20[2]), .QN(n1387) );
  dffs1 \sa00_reg[2]  ( .DIN(N276), .CLK(clk), .Q(sa00[2]), .QN(n1444) );
  dffs1 \sa10_reg[2]  ( .DIN(N260), .CLK(clk), .Q(sa10[2]), .QN(n1389) );
  dffs1 \sa20_reg[3]  ( .DIN(N245), .CLK(clk), .Q(sa20[3]), .QN(n1437) );
  dffs1 \sa00_reg[3]  ( .DIN(N277), .CLK(clk), .Q(sa00[3]) );
  dffs1 \sa30_reg[5]  ( .DIN(N231), .CLK(clk), .Q(sa30[5]), .QN(n1383) );
  dffs1 \sa20_reg[4]  ( .DIN(N246), .CLK(clk), .Q(sa20[4]) );
  dffs1 \sa00_reg[4]  ( .DIN(N278), .CLK(clk), .Q(sa00[4]), .QN(n1531) );
  dffs1 \sa30_reg[6]  ( .DIN(N232), .CLK(clk), .Q(sa30[6]), .QN(n1432) );
  dffs1 \sa20_reg[5]  ( .DIN(N247), .CLK(clk), .Q(sa20[5]), .QN(n1385) );
  dffs1 \sa00_reg[5]  ( .DIN(N279), .CLK(clk), .Q(sa00[5]), .QN(n1401) );
  dffs1 \sa10_reg[5]  ( .DIN(N263), .CLK(clk), .Q(sa10[5]), .QN(n1398) );
  dffs1 \sa20_reg[6]  ( .DIN(N248), .CLK(clk), .QN(n1371) );
  dffs1 \sa00_reg[6]  ( .DIN(N280), .CLK(clk), .Q(sa00[6]) );
  dffs1 \sa10_reg[6]  ( .DIN(N264), .CLK(clk), .Q(sa10[6]) );
  dffs1 \sa30_reg[4]  ( .DIN(N230), .CLK(clk), .Q(sa30[4]) );
  dffs1 \sa30_reg[3]  ( .DIN(N229), .CLK(clk), .Q(sa30[3]) );
  dffs1 \sa30_reg[1]  ( .DIN(N227), .CLK(clk), .Q(sa30[1]), .QN(n1533) );
  dffs1 \sa30_reg[0]  ( .DIN(N226), .CLK(clk), .Q(sa30[0]) );
  dffs1 \sa20_reg[7]  ( .DIN(N249), .CLK(clk), .Q(sa20[7]), .QN(n1423) );
  dffs1 \sa23_reg[7]  ( .DIN(N57), .CLK(clk), .Q(sa23[7]), .QN(n1523) );
  dffs1 \sa22_reg[4]  ( .DIN(N118), .CLK(clk), .Q(sa22[4]), .QN(n1532) );
  dffs1 \sa22_reg[3]  ( .DIN(N117), .CLK(clk), .Q(sa22[3]) );
  dffs1 \sa22_reg[1]  ( .DIN(N115), .CLK(clk), .Q(sa22[1]), .QN(n1431) );
  dffs1 \sa22_reg[0]  ( .DIN(N114), .CLK(clk), .Q(sa22[0]), .QN(n1364) );
  dffs1 \sa12_reg[4]  ( .DIN(N134), .CLK(clk), .Q(sa12[4]), .QN(n1534) );
  dffs1 \sa12_reg[3]  ( .DIN(N133), .CLK(clk), .Q(sa12[3]) );
  dffs1 \sa12_reg[1]  ( .DIN(N131), .CLK(clk), .Q(sa12[1]), .QN(n1433) );
  dffs1 \sa12_reg[0]  ( .DIN(N130), .CLK(clk), .Q(sa12[0]), .QN(n1365) );
  dffs1 \sa21_reg[4]  ( .DIN(N182), .CLK(clk), .Q(sa21[4]), .QN(n1528) );
  dffs1 \sa21_reg[3]  ( .DIN(N181), .CLK(clk), .Q(sa21[3]), .QN(n1510) );
  dffs1 \sa21_reg[1]  ( .DIN(N179), .CLK(clk), .Q(sa21[1]), .QN(n1427) );
  dffs1 \sa21_reg[0]  ( .DIN(N178), .CLK(clk), .Q(sa21[0]), .QN(n1357) );
  dffs1 \sa11_reg[4]  ( .DIN(N198), .CLK(clk), .Q(sa11[4]), .QN(n1530) );
  dffs1 \sa11_reg[3]  ( .DIN(N197), .CLK(clk), .Q(sa11[3]) );
  dffs1 \sa11_reg[1]  ( .DIN(N195), .CLK(clk), .Q(sa11[1]), .QN(n1429) );
  dffs1 \sa11_reg[0]  ( .DIN(N194), .CLK(clk), .Q(sa11[0]), .QN(n1362) );
  dffs1 \sa13_reg[4]  ( .DIN(N70), .CLK(clk), .Q(sa13[4]) );
  dffs1 \sa13_reg[3]  ( .DIN(N69), .CLK(clk), .Q(sa13[3]), .QN(n1436) );
  dffs1 \sa13_reg[1]  ( .DIN(N67), .CLK(clk), .Q(sa13[1]), .QN(n1506) );
  dffs1 \sa13_reg[0]  ( .DIN(N66), .CLK(clk), .Q(sa13[0]), .QN(n1358) );
  dffs1 \sa10_reg[4]  ( .DIN(N262), .CLK(clk), .Q(sa10[4]), .QN(n1527) );
  dffs1 \sa10_reg[3]  ( .DIN(N261), .CLK(clk), .Q(sa10[3]), .QN(n1509) );
  dffs1 \sa10_reg[1]  ( .DIN(N259), .CLK(clk), .Q(sa10[1]), .QN(n1426) );
  dffs1 \sa10_reg[0]  ( .DIN(N258), .CLK(clk), .Q(sa10[0]), .QN(n1356) );
  dffs1 \sa00_reg[7]  ( .DIN(N281), .CLK(clk), .Q(sa00[7]), .QN(n1519) );
  dffs1 \text_out_reg[127]  ( .DIN(N378), .CLK(clk), .Q(\text_out[127] ) );
  dffs1 \text_out_reg[126]  ( .DIN(N379), .CLK(clk), .Q(\text_out[126] ) );
  dffs1 \text_out_reg[125]  ( .DIN(N380), .CLK(clk), .Q(\text_out[125] ) );
  dffs1 \text_out_reg[124]  ( .DIN(N381), .CLK(clk), .Q(\text_out[124] ) );
  dffs1 \text_out_reg[123]  ( .DIN(N382), .CLK(clk), .Q(\text_out[123] ) );
  dffs1 \text_out_reg[122]  ( .DIN(N383), .CLK(clk), .Q(\text_out[122] ) );
  dffs1 \text_out_reg[121]  ( .DIN(N384), .CLK(clk), .Q(\text_out[121] ) );
  dffs1 \text_out_reg[120]  ( .DIN(N385), .CLK(clk), .Q(\text_out[120] ) );
  dffs1 \text_out_reg[95]  ( .DIN(N386), .CLK(clk), .Q(\text_out[95] ) );
  dffs1 \text_out_reg[94]  ( .DIN(N387), .CLK(clk), .Q(\text_out[94] ) );
  dffs1 \text_out_reg[93]  ( .DIN(N388), .CLK(clk), .Q(\text_out[93] ) );
  dffs1 \text_out_reg[92]  ( .DIN(N389), .CLK(clk), .Q(\text_out[92] ) );
  dffs1 \text_out_reg[91]  ( .DIN(N390), .CLK(clk), .Q(\text_out[91] ) );
  dffs1 \text_out_reg[90]  ( .DIN(N391), .CLK(clk), .Q(\text_out[90] ) );
  dffs1 \text_out_reg[89]  ( .DIN(N392), .CLK(clk), .Q(\text_out[89] ) );
  dffs1 \text_out_reg[88]  ( .DIN(N393), .CLK(clk), .Q(\text_out[88] ) );
  dffs1 \text_out_reg[63]  ( .DIN(N394), .CLK(clk), .Q(\text_out[63] ) );
  dffs1 \text_out_reg[62]  ( .DIN(N395), .CLK(clk), .Q(\text_out[62] ) );
  dffs1 \text_out_reg[61]  ( .DIN(N396), .CLK(clk), .Q(\text_out[61] ) );
  dffs1 \text_out_reg[60]  ( .DIN(N397), .CLK(clk), .Q(\text_out[60] ) );
  dffs1 \text_out_reg[59]  ( .DIN(N398), .CLK(clk), .Q(\text_out[59] ) );
  dffs1 \text_out_reg[58]  ( .DIN(N399), .CLK(clk), .Q(\text_out[58] ) );
  dffs1 \text_out_reg[57]  ( .DIN(N400), .CLK(clk), .Q(\text_out[57] ) );
  dffs1 \text_out_reg[56]  ( .DIN(N401), .CLK(clk), .Q(\text_out[56] ) );
  dffs1 \text_out_reg[31]  ( .DIN(N402), .CLK(clk), .Q(\text_out[31] ) );
  dffs1 \text_out_reg[30]  ( .DIN(N403), .CLK(clk), .Q(\text_out[30] ) );
  dffs1 \text_out_reg[29]  ( .DIN(N404), .CLK(clk), .Q(\text_out[29] ) );
  dffs1 \text_out_reg[28]  ( .DIN(N405), .CLK(clk), .Q(\text_out[28] ) );
  dffs1 \text_out_reg[27]  ( .DIN(N406), .CLK(clk), .Q(\text_out[27] ) );
  dffs1 \text_out_reg[26]  ( .DIN(N407), .CLK(clk), .Q(\text_out[26] ) );
  dffs1 \text_out_reg[25]  ( .DIN(n1545), .CLK(clk), .Q(\text_out[25] ) );
  dffs1 \text_out_reg[24]  ( .DIN(N409), .CLK(clk), .Q(\text_out[24] ) );
  dffs1 \text_out_reg[119]  ( .DIN(N410), .CLK(clk), .Q(\text_out[119] ) );
  dffs1 \text_out_reg[118]  ( .DIN(N411), .CLK(clk), .Q(\text_out[118] ) );
  dffs1 \text_out_reg[117]  ( .DIN(N412), .CLK(clk), .Q(\text_out[117] ) );
  dffs1 \text_out_reg[116]  ( .DIN(N413), .CLK(clk), .Q(\text_out[116] ) );
  dffs1 \text_out_reg[115]  ( .DIN(N414), .CLK(clk), .Q(\text_out[115] ) );
  dffs1 \text_out_reg[114]  ( .DIN(N415), .CLK(clk), .Q(\text_out[114] ) );
  dffs1 \text_out_reg[113]  ( .DIN(N416), .CLK(clk), .Q(\text_out[113] ) );
  dffs1 \text_out_reg[112]  ( .DIN(N417), .CLK(clk), .Q(\text_out[112] ) );
  dffs1 \text_out_reg[87]  ( .DIN(N418), .CLK(clk), .Q(\text_out[87] ) );
  dffs1 \text_out_reg[86]  ( .DIN(N419), .CLK(clk), .Q(\text_out[86] ) );
  dffs1 \text_out_reg[85]  ( .DIN(N420), .CLK(clk), .Q(\text_out[85] ) );
  dffs1 \text_out_reg[84]  ( .DIN(N421), .CLK(clk), .Q(\text_out[84] ) );
  dffs1 \text_out_reg[83]  ( .DIN(N422), .CLK(clk), .Q(\text_out[83] ) );
  dffs1 \text_out_reg[82]  ( .DIN(N423), .CLK(clk), .Q(\text_out[82] ) );
  dffs1 \text_out_reg[81]  ( .DIN(N424), .CLK(clk), .Q(\text_out[81] ) );
  dffs1 \text_out_reg[80]  ( .DIN(N425), .CLK(clk), .Q(\text_out[80] ) );
  dffs1 \text_out_reg[55]  ( .DIN(N426), .CLK(clk), .Q(\text_out[55] ) );
  dffs1 \text_out_reg[54]  ( .DIN(N427), .CLK(clk), .Q(\text_out[54] ) );
  dffs1 \text_out_reg[53]  ( .DIN(N428), .CLK(clk), .Q(\text_out[53] ) );
  dffs1 \text_out_reg[52]  ( .DIN(N429), .CLK(clk), .Q(\text_out[52] ) );
  dffs1 \text_out_reg[51]  ( .DIN(N430), .CLK(clk), .Q(\text_out[51] ) );
  dffs1 \text_out_reg[50]  ( .DIN(N431), .CLK(clk), .Q(\text_out[50] ) );
  dffs1 \text_out_reg[49]  ( .DIN(N432), .CLK(clk), .Q(\text_out[49] ) );
  dffs1 \text_out_reg[48]  ( .DIN(N433), .CLK(clk), .Q(\text_out[48] ) );
  dffs1 \text_out_reg[23]  ( .DIN(N434), .CLK(clk), .Q(\text_out[23] ) );
  dffs1 \text_out_reg[22]  ( .DIN(N435), .CLK(clk), .Q(\text_out[22] ) );
  dffs1 \text_out_reg[21]  ( .DIN(N436), .CLK(clk), .Q(\text_out[21] ) );
  dffs1 \text_out_reg[20]  ( .DIN(N437), .CLK(clk), .Q(\text_out[20] ) );
  dffs1 \text_out_reg[19]  ( .DIN(N438), .CLK(clk), .Q(\text_out[19] ) );
  dffs1 \text_out_reg[18]  ( .DIN(N439), .CLK(clk), .Q(\text_out[18] ) );
  dffs1 \text_out_reg[17]  ( .DIN(n1544), .CLK(clk), .Q(\text_out[17] ) );
  dffs1 \text_out_reg[16]  ( .DIN(N441), .CLK(clk), .Q(\text_out[16] ) );
  dffs1 \text_out_reg[111]  ( .DIN(N442), .CLK(clk), .Q(\text_out[111] ) );
  dffs1 \text_out_reg[110]  ( .DIN(N443), .CLK(clk), .Q(\text_out[110] ) );
  dffs1 \text_out_reg[109]  ( .DIN(N444), .CLK(clk), .Q(\text_out[109] ) );
  dffs1 \text_out_reg[108]  ( .DIN(N445), .CLK(clk), .Q(\text_out[108] ) );
  dffs1 \text_out_reg[107]  ( .DIN(N446), .CLK(clk), .Q(\text_out[107] ) );
  dffs1 \text_out_reg[106]  ( .DIN(N447), .CLK(clk), .Q(\text_out[106] ) );
  dffs1 \text_out_reg[105]  ( .DIN(N448), .CLK(clk), .Q(\text_out[105] ) );
  dffs1 \text_out_reg[104]  ( .DIN(N449), .CLK(clk), .Q(\text_out[104] ) );
  dffs1 \text_out_reg[79]  ( .DIN(N450), .CLK(clk), .Q(\text_out[79] ) );
  dffs1 \text_out_reg[78]  ( .DIN(N451), .CLK(clk), .Q(\text_out[78] ) );
  dffs1 \text_out_reg[77]  ( .DIN(N452), .CLK(clk), .Q(\text_out[77] ) );
  dffs1 \text_out_reg[76]  ( .DIN(N453), .CLK(clk), .Q(\text_out[76] ) );
  dffs1 \text_out_reg[75]  ( .DIN(N454), .CLK(clk), .Q(\text_out[75] ) );
  dffs1 \text_out_reg[74]  ( .DIN(N455), .CLK(clk), .Q(\text_out[74] ) );
  dffs1 \text_out_reg[73]  ( .DIN(N456), .CLK(clk), .Q(\text_out[73] ) );
  dffs1 \text_out_reg[72]  ( .DIN(N457), .CLK(clk), .Q(\text_out[72] ) );
  dffs1 \text_out_reg[47]  ( .DIN(N458), .CLK(clk), .Q(\text_out[47] ) );
  dffs1 \text_out_reg[46]  ( .DIN(N459), .CLK(clk), .Q(\text_out[46] ) );
  dffs1 \text_out_reg[45]  ( .DIN(N460), .CLK(clk), .Q(\text_out[45] ) );
  dffs1 \text_out_reg[44]  ( .DIN(N461), .CLK(clk), .Q(\text_out[44] ) );
  dffs1 \text_out_reg[43]  ( .DIN(N462), .CLK(clk), .Q(\text_out[43] ) );
  dffs1 \text_out_reg[42]  ( .DIN(N463), .CLK(clk), .Q(\text_out[42] ) );
  dffs1 \text_out_reg[41]  ( .DIN(N464), .CLK(clk), .Q(\text_out[41] ) );
  dffs1 \text_out_reg[40]  ( .DIN(N465), .CLK(clk), .Q(\text_out[40] ) );
  dffs1 \text_out_reg[15]  ( .DIN(N466), .CLK(clk), .Q(\text_out[15] ) );
  dffs1 \text_out_reg[14]  ( .DIN(N467), .CLK(clk), .Q(\text_out[14] ) );
  dffs1 \text_out_reg[13]  ( .DIN(N468), .CLK(clk), .Q(\text_out[13] ) );
  dffs1 \text_out_reg[12]  ( .DIN(N469), .CLK(clk), .Q(\text_out[12] ) );
  dffs1 \text_out_reg[11]  ( .DIN(N470), .CLK(clk), .Q(\text_out[11] ) );
  dffs1 \text_out_reg[10]  ( .DIN(N471), .CLK(clk), .Q(\text_out[10] ) );
  dffs1 \text_out_reg[9]  ( .DIN(N472), .CLK(clk), .Q(\text_out[9] ) );
  dffs1 \text_out_reg[8]  ( .DIN(n1549), .CLK(clk), .Q(\text_out[8] ) );
  dffs1 \text_out_reg[103]  ( .DIN(N474), .CLK(clk), .Q(\text_out[103] ) );
  dffs1 \text_out_reg[102]  ( .DIN(N475), .CLK(clk), .Q(\text_out[102] ) );
  dffs1 \text_out_reg[101]  ( .DIN(N476), .CLK(clk), .Q(\text_out[101] ) );
  dffs1 \text_out_reg[100]  ( .DIN(N477), .CLK(clk), .Q(\text_out[100] ) );
  dffs1 \text_out_reg[99]  ( .DIN(N478), .CLK(clk), .Q(\text_out[99] ) );
  dffs1 \text_out_reg[98]  ( .DIN(N479), .CLK(clk), .Q(\text_out[98] ) );
  dffs1 \text_out_reg[97]  ( .DIN(N480), .CLK(clk), .Q(\text_out[97] ) );
  dffs1 \text_out_reg[96]  ( .DIN(N481), .CLK(clk), .Q(\text_out[96] ) );
  dffs1 \text_out_reg[71]  ( .DIN(N482), .CLK(clk), .Q(\text_out[71] ) );
  dffs1 \text_out_reg[70]  ( .DIN(N483), .CLK(clk), .Q(\text_out[70] ) );
  dffs1 \text_out_reg[69]  ( .DIN(N484), .CLK(clk), .Q(\text_out[69] ) );
  dffs1 \text_out_reg[68]  ( .DIN(N485), .CLK(clk), .Q(\text_out[68] ) );
  dffs1 \text_out_reg[67]  ( .DIN(N486), .CLK(clk), .Q(\text_out[67] ) );
  dffs1 \text_out_reg[66]  ( .DIN(N487), .CLK(clk), .Q(\text_out[66] ) );
  dffs1 \text_out_reg[65]  ( .DIN(N488), .CLK(clk), .Q(\text_out[65] ) );
  dffs1 \text_out_reg[64]  ( .DIN(N489), .CLK(clk), .Q(\text_out[64] ) );
  dffs1 \text_out_reg[39]  ( .DIN(N490), .CLK(clk), .Q(\text_out[39] ) );
  dffs1 \text_out_reg[38]  ( .DIN(N491), .CLK(clk), .Q(\text_out[38] ) );
  dffs1 \text_out_reg[37]  ( .DIN(N492), .CLK(clk), .Q(\text_out[37] ) );
  dffs1 \text_out_reg[36]  ( .DIN(N493), .CLK(clk), .Q(\text_out[36] ) );
  dffs1 \text_out_reg[35]  ( .DIN(N494), .CLK(clk), .Q(\text_out[35] ) );
  dffs1 \text_out_reg[34]  ( .DIN(N495), .CLK(clk), .Q(\text_out[34] ) );
  dffs1 \text_out_reg[33]  ( .DIN(N496), .CLK(clk), .Q(\text_out[33] ) );
  dffs1 \text_out_reg[32]  ( .DIN(N497), .CLK(clk), .Q(\text_out[32] ) );
  dffs1 \text_out_reg[7]  ( .DIN(N498), .CLK(clk), .Q(\text_out[7] ) );
  dffs1 \text_out_reg[6]  ( .DIN(N499), .CLK(clk), .Q(\text_out[6] ) );
  dffs1 \text_out_reg[5]  ( .DIN(N500), .CLK(clk), .Q(\text_out[5] ) );
  dffs1 \text_out_reg[4]  ( .DIN(N501), .CLK(clk), .Q(\text_out[4] ) );
  dffs1 \text_out_reg[3]  ( .DIN(N502), .CLK(clk), .Q(\text_out[3] ) );
  dffs1 \text_out_reg[2]  ( .DIN(N503), .CLK(clk), .Q(\text_out[2] ) );
  dffs1 \text_out_reg[1]  ( .DIN(n1550), .CLK(clk), .Q(\text_out[1] ) );
  dffs1 \text_out_reg[0]  ( .DIN(N505), .CLK(clk), .Q(\text_out[0] ) );
  dffs1 \u0/w_reg[1][15]  ( .DIN(\u0/N123 ), .CLK(clk), .Q(w1[15]), .QN(n1491)
         );
  dffs1 \u0/w_reg[2][15]  ( .DIN(\u0/N189 ), .CLK(clk), .Q(w2[15]), .QN(n1458)
         );
  dffs1 \u0/w_reg[1][23]  ( .DIN(\u0/N131 ), .CLK(clk), .Q(w1[23]), .QN(n1487)
         );
  dffs1 \u0/w_reg[2][23]  ( .DIN(\u0/N197 ), .CLK(clk), .Q(w2[23]) );
  dffs1 \u0/w_reg[1][31]  ( .DIN(\u0/N139 ), .CLK(clk), .Q(w1[31]) );
  dffs1 \u0/w_reg[2][31]  ( .DIN(\u0/N205 ), .CLK(clk), .Q(w2[31]), .QN(n1451)
         );
  dffs1 \u0/w_reg[1][7]  ( .DIN(\u0/N115 ), .CLK(clk), .Q(w1[7]) );
  dffs1 \u0/w_reg[2][7]  ( .DIN(\u0/N181 ), .CLK(clk), .Q(w2[7]) );
  dffs1 \u0/w_reg[3][7]  ( .DIN(\u0/N247 ), .CLK(clk), .Q(w3[7]), .QN(n1442)
         );
  dffs1 \u0/w_reg[0][7]  ( .DIN(\u0/N49 ), .CLK(clk), .Q(w0[7]) );
  dffs1 \u0/w_reg[1][6]  ( .DIN(\u0/N114 ), .CLK(clk), .Q(w1[6]), .QN(n1542)
         );
  dffs1 \u0/w_reg[2][6]  ( .DIN(\u0/N180 ), .CLK(clk), .Q(w2[6]) );
  dffs1 \u0/w_reg[3][6]  ( .DIN(\u0/N246 ), .CLK(clk), .Q(w3[6]), .QN(n1391)
         );
  dffs1 \u0/w_reg[0][6]  ( .DIN(\u0/N48 ), .CLK(clk), .Q(w0[6]), .QN(n1504) );
  dffs1 \u0/w_reg[1][5]  ( .DIN(\u0/N113 ), .CLK(clk), .Q(w1[5]), .QN(n1495)
         );
  dffs1 \u0/w_reg[2][5]  ( .DIN(\u0/N179 ), .CLK(clk), .Q(w2[5]), .QN(n1462)
         );
  dffs1 \u0/w_reg[3][5]  ( .DIN(\u0/N245 ), .CLK(clk), .Q(w3[5]), .QN(n1375)
         );
  dffs1 \u0/w_reg[0][5]  ( .DIN(\u0/N47 ), .CLK(clk), .Q(w0[5]), .QN(n1471) );
  dffs1 \u0/w_reg[1][4]  ( .DIN(\u0/N112 ), .CLK(clk), .Q(w1[4]), .QN(n1496)
         );
  dffs1 \u0/w_reg[2][4]  ( .DIN(\u0/N178 ), .CLK(clk), .Q(w2[4]), .QN(n1478)
         );
  dffs1 \u0/w_reg[3][4]  ( .DIN(\u0/N244 ), .CLK(clk), .Q(w3[4]), .QN(n1441)
         );
  dffs1 \u0/w_reg[0][4]  ( .DIN(\u0/N46 ), .CLK(clk), .Q(w0[4]), .QN(n1472) );
  dffs1 \u0/w_reg[1][3]  ( .DIN(\u0/N111 ), .CLK(clk), .Q(w1[3]) );
  dffs1 \u0/w_reg[2][3]  ( .DIN(\u0/N177 ), .CLK(clk), .Q(w2[3]), .QN(n1484)
         );
  dffs1 \u0/w_reg[3][3]  ( .DIN(\u0/N243 ), .CLK(clk), .Q(w3[3]), .QN(n1440)
         );
  dffs1 \u0/w_reg[0][3]  ( .DIN(\u0/N45 ), .CLK(clk), .Q(w0[3]), .QN(n1505) );
  dffs1 \u0/w_reg[1][2]  ( .DIN(\u0/N110 ), .CLK(clk), .Q(w1[2]) );
  dffs1 \u0/w_reg[2][2]  ( .DIN(\u0/N176 ), .CLK(clk), .Q(w2[2]) );
  dffs1 \u0/w_reg[3][2]  ( .DIN(\u0/N242 ), .CLK(clk), .Q(w3[2]), .QN(n1369)
         );
  dffs1 \u0/w_reg[0][2]  ( .DIN(\u0/N44 ), .CLK(clk), .Q(w0[2]) );
  dffs1 \u0/w_reg[1][1]  ( .DIN(\u0/N109 ), .CLK(clk), .Q(w1[1]) );
  dffs1 \u0/w_reg[2][1]  ( .DIN(\u0/N175 ), .CLK(clk), .Q(w2[1]), .QN(n1479)
         );
  dffs1 \u0/w_reg[3][1]  ( .DIN(\u0/N241 ), .CLK(clk), .Q(w3[1]), .QN(n1411)
         );
  dffs1 \u0/w_reg[0][1]  ( .DIN(\u0/N43 ), .CLK(clk), .Q(w0[1]) );
  dffs1 \u0/w_reg[1][0]  ( .DIN(\u0/N108 ), .CLK(clk), .Q(w1[0]), .QN(n1497)
         );
  dffs1 \u0/w_reg[2][0]  ( .DIN(\u0/N174 ), .CLK(clk), .Q(w2[0]), .QN(n1450)
         );
  dffs1 \u0/w_reg[0][0]  ( .DIN(\u0/N42 ), .CLK(clk), .Q(w0[0]), .QN(n1473) );
  dffs1 \u0/w_reg[3][31]  ( .DIN(\u0/N271 ), .CLK(clk), .Q(w3[31]), .QN(n1416)
         );
  dffs1 \u0/w_reg[0][31]  ( .DIN(\u0/N73 ), .CLK(clk), .Q(w0[31]) );
  dffs1 \u0/w_reg[1][30]  ( .DIN(\u0/N138 ), .CLK(clk), .Q(w1[30]) );
  dffs1 \u0/w_reg[2][30]  ( .DIN(\u0/N204 ), .CLK(clk), .Q(w2[30]) );
  dffs1 \u0/w_reg[3][30]  ( .DIN(\u0/N270 ), .CLK(clk), .Q(w3[30]), .QN(n1475)
         );
  dffs1 \u0/w_reg[0][30]  ( .DIN(\u0/N72 ), .CLK(clk), .Q(w0[30]) );
  dffs1 \u0/w_reg[1][29]  ( .DIN(\u0/N137 ), .CLK(clk), .Q(w1[29]), .QN(n1485)
         );
  dffs1 \u0/w_reg[2][29]  ( .DIN(\u0/N203 ), .CLK(clk), .Q(w2[29]), .QN(n1452)
         );
  dffs1 \u0/w_reg[3][29]  ( .DIN(\u0/N269 ), .CLK(clk), .Q(w3[29]), .QN(n1374)
         );
  dffs1 \u0/w_reg[0][29]  ( .DIN(\u0/N71 ), .CLK(clk), .Q(w0[29]), .QN(n1480)
         );
  dffs1 \u0/w_reg[1][28]  ( .DIN(\u0/N136 ), .CLK(clk), .Q(w1[28]), .QN(n1541)
         );
  dffs1 \u0/w_reg[2][28]  ( .DIN(\u0/N202 ), .CLK(clk), .Q(w2[28]), .QN(n1477)
         );
  dffs1 \u0/w_reg[3][28]  ( .DIN(\u0/N268 ), .CLK(clk), .Q(w3[28]), .QN(n1392)
         );
  dffs1 \u0/w_reg[0][28]  ( .DIN(\u0/N70 ), .CLK(clk), .Q(w0[28]), .QN(n1540)
         );
  dffs1 \u0/w_reg[1][27]  ( .DIN(\u0/N135 ), .CLK(clk), .Q(w1[27]) );
  dffs1 \u0/w_reg[2][27]  ( .DIN(\u0/N201 ), .CLK(clk), .Q(w2[27]) );
  dffs1 \u0/w_reg[3][27]  ( .DIN(\u0/N267 ), .CLK(clk), .Q(w3[27]), .QN(n1476)
         );
  dffs1 \u0/w_reg[0][27]  ( .DIN(\u0/N69 ), .CLK(clk), .Q(w0[27]) );
  dffs1 \u0/w_reg[1][26]  ( .DIN(\u0/N134 ), .CLK(clk), .Q(w1[26]) );
  dffs1 \u0/w_reg[2][26]  ( .DIN(\u0/N200 ), .CLK(clk), .Q(w2[26]), .QN(n1453)
         );
  dffs1 \u0/w_reg[3][26]  ( .DIN(\u0/N266 ), .CLK(clk), .Q(w3[26]), .QN(n1548)
         );
  dffs1 \u0/w_reg[0][26]  ( .DIN(\u0/N68 ), .CLK(clk), .Q(w0[26]) );
  dffs1 \u0/w_reg[1][25]  ( .DIN(\u0/N133 ), .CLK(clk), .Q(w1[25]) );
  dffs1 \u0/w_reg[2][25]  ( .DIN(\u0/N199 ), .CLK(clk), .Q(w2[25]) );
  dffs1 \u0/w_reg[3][25]  ( .DIN(\u0/N265 ), .CLK(clk), .Q(w3[25]), .QN(n1410)
         );
  dffs1 \u0/w_reg[0][25]  ( .DIN(\u0/N67 ), .CLK(clk), .Q(w0[25]) );
  dffs1 \u0/w_reg[1][24]  ( .DIN(\u0/N132 ), .CLK(clk), .Q(w1[24]), .QN(n1486)
         );
  dffs1 \u0/w_reg[2][24]  ( .DIN(\u0/N198 ), .CLK(clk), .Q(w2[24]), .QN(n1454)
         );
  dffs1 \u0/w_reg[3][24]  ( .DIN(\u0/N264 ), .CLK(clk), .Q(w3[24]), .QN(n1554)
         );
  dffs1 \u0/w_reg[0][24]  ( .DIN(\u0/N66 ), .CLK(clk), .Q(w0[24]), .QN(n1481)
         );
  dffs1 \u0/w_reg[3][23]  ( .DIN(\u0/N263 ), .CLK(clk), .Q(w3[23]), .QN(n1415)
         );
  dffs1 \u0/w_reg[0][23]  ( .DIN(\u0/N65 ), .CLK(clk), .Q(w0[23]), .QN(n1463)
         );
  dffs1 \u0/w_reg[1][22]  ( .DIN(\u0/N130 ), .CLK(clk), .Q(w1[22]) );
  dffs1 \u0/w_reg[2][22]  ( .DIN(\u0/N196 ), .CLK(clk), .Q(w2[22]), .QN(n1482)
         );
  dffs1 \u0/w_reg[3][22]  ( .DIN(\u0/N262 ), .CLK(clk), .Q(w3[22]), .QN(n1438)
         );
  dffs1 \u0/w_reg[0][22]  ( .DIN(\u0/N64 ), .CLK(clk), .Q(w0[22]) );
  dffs1 \u0/w_reg[1][21]  ( .DIN(\u0/N129 ), .CLK(clk), .Q(w1[21]) );
  dffs1 \u0/w_reg[2][21]  ( .DIN(\u0/N195 ), .CLK(clk), .Q(w2[21]) );
  dffs1 \u0/w_reg[3][21]  ( .DIN(\u0/N261 ), .CLK(clk), .Q(w3[21]), .QN(n1373)
         );
  dffs1 \u0/w_reg[0][21]  ( .DIN(\u0/N63 ), .CLK(clk), .Q(w0[21]) );
  dffs1 \u0/w_reg[1][20]  ( .DIN(\u0/N128 ), .CLK(clk), .Q(w1[20]), .QN(n1488)
         );
  dffs1 \u0/w_reg[2][20]  ( .DIN(\u0/N194 ), .CLK(clk), .Q(w2[20]), .QN(n1455)
         );
  dffs1 \u0/w_reg[3][20]  ( .DIN(\u0/N260 ), .CLK(clk), .Q(w3[20]), .QN(n1376)
         );
  dffs1 \u0/w_reg[0][20]  ( .DIN(\u0/N62 ), .CLK(clk), .Q(w0[20]), .QN(n1464)
         );
  dffs1 \u0/w_reg[1][19]  ( .DIN(\u0/N127 ), .CLK(clk), .Q(w1[19]) );
  dffs1 \u0/w_reg[2][19]  ( .DIN(\u0/N193 ), .CLK(clk), .Q(w2[19]), .QN(n1483)
         );
  dffs1 \u0/w_reg[3][19]  ( .DIN(\u0/N259 ), .CLK(clk), .Q(w3[19]), .QN(n1439)
         );
  dffs1 \u0/w_reg[0][19]  ( .DIN(\u0/N61 ), .CLK(clk), .Q(w0[19]), .QN(n1500)
         );
  dffs1 \u0/w_reg[1][18]  ( .DIN(\u0/N126 ), .CLK(clk), .Q(w1[18]), .QN(n1489)
         );
  dffs1 \u0/w_reg[2][18]  ( .DIN(\u0/N192 ), .CLK(clk), .Q(w2[18]) );
  dffs1 \u0/w_reg[3][18]  ( .DIN(\u0/N258 ), .CLK(clk), .Q(w3[18]), .QN(n1368)
         );
  dffs1 \u0/w_reg[0][18]  ( .DIN(\u0/N60 ), .CLK(clk), .Q(w0[18]), .QN(n1465)
         );
  dffs1 \u0/w_reg[1][17]  ( .DIN(\u0/N125 ), .CLK(clk), .Q(w1[17]) );
  dffs1 \u0/w_reg[2][17]  ( .DIN(\u0/N191 ), .CLK(clk), .Q(w2[17]), .QN(n1456)
         );
  dffs1 \u0/w_reg[3][17]  ( .DIN(\u0/N257 ), .CLK(clk), .Q(w3[17]), .QN(n1412)
         );
  dffs1 \u0/w_reg[0][17]  ( .DIN(\u0/N59 ), .CLK(clk), .Q(w0[17]), .QN(n1501)
         );
  dffs1 \u0/w_reg[1][16]  ( .DIN(\u0/N124 ), .CLK(clk), .Q(w1[16]), .QN(n1490)
         );
  dffs1 \u0/w_reg[2][16]  ( .DIN(\u0/N190 ), .CLK(clk), .Q(w2[16]), .QN(n1457)
         );
  dffs1 \u0/w_reg[3][16]  ( .DIN(\u0/N256 ), .CLK(clk), .Q(w3[16]), .QN(n1558)
         );
  dffs1 \u0/w_reg[0][16]  ( .DIN(\u0/N58 ), .CLK(clk), .Q(w0[16]), .QN(n1466)
         );
  dffs1 \u0/w_reg[3][15]  ( .DIN(\u0/N255 ), .CLK(clk), .Q(w3[15]), .QN(n1414)
         );
  dffs1 \u0/w_reg[0][15]  ( .DIN(\u0/N57 ), .CLK(clk), .Q(w0[15]), .QN(n1467)
         );
  dffs1 \u0/w_reg[1][14]  ( .DIN(\u0/N122 ), .CLK(clk), .Q(w1[14]) );
  dffs1 \u0/w_reg[2][14]  ( .DIN(\u0/N188 ), .CLK(clk), .Q(w2[14]) );
  dffs1 \u0/w_reg[3][14]  ( .DIN(\u0/N254 ), .CLK(clk), .Q(w3[14]), .QN(n1474)
         );
  dffs1 \u0/w_reg[0][14]  ( .DIN(\u0/N56 ), .CLK(clk), .Q(w0[14]), .QN(n1502)
         );
  dffs1 \u0/w_reg[1][13]  ( .DIN(\u0/N121 ), .CLK(clk), .Q(w1[13]), .QN(n1492)
         );
  dffs1 \u0/w_reg[2][13]  ( .DIN(\u0/N187 ), .CLK(clk), .Q(w2[13]), .QN(n1459)
         );
  dffs1 \u0/w_reg[3][13]  ( .DIN(\u0/N253 ), .CLK(clk), .Q(w3[13]), .QN(n1372)
         );
  dffs1 \u0/w_reg[0][13]  ( .DIN(\u0/N55 ), .CLK(clk), .Q(w0[13]), .QN(n1468)
         );
  dffs1 \u0/w_reg[1][12]  ( .DIN(\u0/N120 ), .CLK(clk), .Q(w1[12]), .QN(n1493)
         );
  dffs1 \u0/w_reg[2][12]  ( .DIN(\u0/N186 ), .CLK(clk), .Q(w2[12]), .QN(n1460)
         );
  dffs1 \u0/w_reg[3][12]  ( .DIN(\u0/N252 ), .CLK(clk), .Q(w3[12]), .QN(n1393)
         );
  dffs1 \u0/w_reg[0][12]  ( .DIN(\u0/N54 ), .CLK(clk), .Q(w0[12]), .QN(n1469)
         );
  dffs1 \u0/w_reg[1][11]  ( .DIN(\u0/N119 ), .CLK(clk), .Q(w1[11]) );
  dffs1 \u0/w_reg[2][11]  ( .DIN(\u0/N185 ), .CLK(clk), .Q(w2[11]) );
  dffs1 \u0/w_reg[3][11]  ( .DIN(\u0/N251 ), .CLK(clk), .Q(w3[11]), .QN(n1413)
         );
  dffs1 \u0/w_reg[0][11]  ( .DIN(\u0/N53 ), .CLK(clk), .Q(w0[11]) );
  dffs1 \u0/w_reg[1][10]  ( .DIN(\u0/N118 ), .CLK(clk), .Q(w1[10]) );
  dffs1 \u0/w_reg[2][10]  ( .DIN(\u0/N184 ), .CLK(clk), .Q(w2[10]) );
  dffs1 \u0/w_reg[3][10]  ( .DIN(\u0/N250 ), .CLK(clk), .Q(w3[10]), .QN(n1553)
         );
  dffs1 \u0/w_reg[0][10]  ( .DIN(\u0/N52 ), .CLK(clk), .Q(w0[10]), .QN(n1499)
         );
  dffs1 \u0/w_reg[1][9]  ( .DIN(\u0/N117 ), .CLK(clk), .Q(w1[9]) );
  dffs1 \u0/w_reg[2][9]  ( .DIN(\u0/N183 ), .CLK(clk), .Q(w2[9]) );
  dffs1 \u0/w_reg[3][9]  ( .DIN(\u0/N249 ), .CLK(clk), .Q(w3[9]), .QN(n1547)
         );
  dffs1 \u0/w_reg[0][9]  ( .DIN(\u0/N51 ), .CLK(clk), .Q(w0[9]), .QN(n1503) );
  dffs1 \u0/w_reg[1][8]  ( .DIN(\u0/N116 ), .CLK(clk), .Q(w1[8]), .QN(n1494)
         );
  dffs1 \u0/w_reg[2][8]  ( .DIN(\u0/N182 ), .CLK(clk), .Q(w2[8]), .QN(n1461)
         );
  dffs1 \u0/w_reg[3][8]  ( .DIN(\u0/N248 ), .CLK(clk), .Q(w3[8]), .QN(n1361)
         );
  dffs1 \u0/w_reg[0][8]  ( .DIN(\u0/N50 ), .CLK(clk), .Q(w0[8]), .QN(n1470) );
  dffs1 \u0/w_reg[3][0]  ( .DIN(\u0/N240 ), .CLK(clk), .Q(w3[0]), .QN(n1556)
         );
  dffs1 \u0/r0/out_reg[31]  ( .DIN(\u0/r0/N77 ), .CLK(clk), .QN(n15588) );
  dffs1 \u0/r0/out_reg[29]  ( .DIN(\u0/r0/N75 ), .CLK(clk), .QN(n15586) );
  dffs1 \u0/r0/out_reg[27]  ( .DIN(\u0/r0/N73 ), .CLK(clk), .QN(n15584) );
  dffs1 \u0/r0/out_reg[30]  ( .DIN(\u0/r0/N76 ), .CLK(clk), .QN(n15587) );
  dffs1 \u0/r0/out_reg[28]  ( .DIN(\u0/r0/N74 ), .CLK(clk), .QN(n15585) );
  dffs1 \u0/r0/out_reg[26]  ( .DIN(\u0/r0/N72 ), .CLK(clk), .QN(n15583) );
  dffs1 \u0/r0/out_reg[25]  ( .DIN(\u0/r0/N71 ), .CLK(clk), .QN(n15582) );
  dffs1 \u0/r0/rcnt_reg[3]  ( .DIN(\u0/r0/N81 ), .CLK(clk), .QN(\u0/r0/n3 ) );
  dffs1 \u0/r0/out_reg[24]  ( .DIN(\u0/r0/N70 ), .CLK(clk), .QN(n15581) );
  dffs1 \u0/r0/rcnt_reg[2]  ( .DIN(\u0/r0/N80 ), .CLK(clk), 
        .Q(\u0/r0/rcnt[2]), .QN(n1419) );
  dffs1 \u0/r0/rcnt_reg[1]  ( .DIN(\u0/r0/N79 ), .CLK(clk), 
        .Q(\u0/r0/rcnt[1]) );
  dffs1 \u0/r0/rcnt_reg[0]  ( .DIN(\u0/r0/N78 ), .CLK(clk), 
        .Q(\u0/r0/rcnt[0]), .QN(n1498) );
  xnr2s1 U1609 ( .DIN1(n1412), .DIN2(n4837), .Q(N440) );
  hi1s1 U1610 ( .DIN(N440), .Q(n1544) );
  xnr2s1 U1611 ( .DIN1(n1410), .DIN2(n5223), .Q(N408) );
  hi1s1 U1612 ( .DIN(N408), .Q(n1545) );
  xnr2s1 U1613 ( .DIN1(n4845), .DIN2(n4941), .Q(n4834) );
  hi1s1 U1614 ( .DIN(n4834), .Q(n1546) );
  xnr2s1 U1615 ( .DIN1(n1361), .DIN2(n4931), .Q(N473) );
  hi1s1 U1616 ( .DIN(N473), .Q(n1549) );
  xnr2s1 U1617 ( .DIN1(n1411), .DIN2(n5007), .Q(N504) );
  hi1s1 U1618 ( .DIN(N504), .Q(n1550) );
  xnr2s1 U1619 ( .DIN1(n1412), .DIN2(n4933), .Q(n4932) );
  hi1s1 U1620 ( .DIN(n4932), .Q(n1551) );
  xnr2s1 U1621 ( .DIN1(n4837), .DIN2(n5223), .Q(n4826) );
  hi1s1 U1622 ( .DIN(n4826), .Q(n1552) );
  hi1s1 U1623 ( .DIN(n1554), .Q(n1555) );
  hi1s1 U1624 ( .DIN(n1556), .Q(n1557) );
  hi1s1 U1625 ( .DIN(n1558), .Q(n1559) );
  nb1s1 U1626 ( .DIN(n1588), .Q(n1560) );
  nb1s1 U1627 ( .DIN(n1593), .Q(n1561) );
  nb1s1 U1628 ( .DIN(n1593), .Q(n1562) );
  nb1s1 U1629 ( .DIN(n1593), .Q(n1563) );
  nb1s1 U1630 ( .DIN(n1593), .Q(n1564) );
  nb1s1 U1631 ( .DIN(n1592), .Q(n1565) );
  nb1s1 U1632 ( .DIN(n1592), .Q(n1566) );
  nb1s1 U1633 ( .DIN(n1592), .Q(n1567) );
  nb1s1 U1634 ( .DIN(n1591), .Q(n1568) );
  nb1s1 U1635 ( .DIN(n1591), .Q(n1569) );
  nb1s1 U1636 ( .DIN(n1591), .Q(n1570) );
  nb1s1 U1637 ( .DIN(n1590), .Q(n1571) );
  nb1s1 U1638 ( .DIN(n1590), .Q(n1572) );
  nb1s1 U1639 ( .DIN(n1590), .Q(n1573) );
  nb1s1 U1640 ( .DIN(n1589), .Q(n1574) );
  nb1s1 U1641 ( .DIN(n1589), .Q(n1575) );
  nb1s1 U1642 ( .DIN(n1589), .Q(n1576) );
  nb1s1 U1643 ( .DIN(n1591), .Q(n1577) );
  nb1s1 U1644 ( .DIN(n1590), .Q(n1578) );
  nb1s1 U1645 ( .DIN(n1589), .Q(n1579) );
  nb1s1 U1646 ( .DIN(n1593), .Q(n1580) );
  nb1s1 U1647 ( .DIN(n1592), .Q(n1581) );
  nb1s1 U1648 ( .DIN(n1588), .Q(n1582) );
  nb1s1 U1649 ( .DIN(n1591), .Q(n1583) );
  nb1s1 U1650 ( .DIN(n1590), .Q(n1584) );
  nb1s1 U1651 ( .DIN(n1589), .Q(n1585) );
  nb1s1 U1652 ( .DIN(n1588), .Q(n1586) );
  nb1s1 U1653 ( .DIN(n1588), .Q(n1587) );
  nb1s1 U1654 ( .DIN(n1669), .Q(n1588) );
  nb1s1 U1655 ( .DIN(n1669), .Q(n1589) );
  nb1s1 U1656 ( .DIN(n1669), .Q(n1590) );
  nb1s1 U1657 ( .DIN(n1669), .Q(n1591) );
  nb1s1 U1658 ( .DIN(n1669), .Q(n1592) );
  nb1s1 U1659 ( .DIN(n1669), .Q(n1593) );
  hi1s1 U1660 ( .DIN(n1640), .Q(n1594) );
  hi1s1 U1661 ( .DIN(n1639), .Q(n1595) );
  hi1s1 U1662 ( .DIN(n1641), .Q(n1596) );
  hi1s1 U1663 ( .DIN(n1639), .Q(n1597) );
  hi1s1 U1664 ( .DIN(n1642), .Q(n1598) );
  hi1s1 U1665 ( .DIN(n1639), .Q(n1599) );
  hi1s1 U1666 ( .DIN(n1642), .Q(n1600) );
  hi1s1 U1667 ( .DIN(n1640), .Q(n1601) );
  hi1s1 U1668 ( .DIN(n1642), .Q(n1602) );
  hi1s1 U1669 ( .DIN(n1640), .Q(n1603) );
  hi1s1 U1670 ( .DIN(n1643), .Q(n1604) );
  hi1s1 U1671 ( .DIN(n1641), .Q(n1605) );
  hi1s1 U1672 ( .DIN(n1643), .Q(n1606) );
  hi1s1 U1673 ( .DIN(n1641), .Q(n1607) );
  hi1s1 U1674 ( .DIN(n1653), .Q(n1608) );
  hi1s1 U1675 ( .DIN(n1652), .Q(n1609) );
  hi1s1 U1676 ( .DIN(n1652), .Q(n1610) );
  hi1s1 U1677 ( .DIN(n1652), .Q(n1611) );
  hi1s1 U1678 ( .DIN(n1651), .Q(n1612) );
  hi1s1 U1679 ( .DIN(n1651), .Q(n1613) );
  hi1s1 U1680 ( .DIN(n1651), .Q(n1614) );
  hi1s1 U1681 ( .DIN(n1650), .Q(n1615) );
  hi1s1 U1682 ( .DIN(n1650), .Q(n1616) );
  hi1s1 U1683 ( .DIN(n1650), .Q(n1617) );
  hi1s1 U1684 ( .DIN(n1649), .Q(n1618) );
  hi1s1 U1685 ( .DIN(n1649), .Q(n1619) );
  hi1s1 U1686 ( .DIN(n1649), .Q(n1620) );
  hi1s1 U1687 ( .DIN(n1648), .Q(n1621) );
  hi1s1 U1688 ( .DIN(n1648), .Q(n1622) );
  hi1s1 U1689 ( .DIN(n1648), .Q(n1623) );
  hi1s1 U1690 ( .DIN(n1647), .Q(n1624) );
  hi1s1 U1691 ( .DIN(n1647), .Q(n1625) );
  hi1s1 U1692 ( .DIN(n1647), .Q(n1626) );
  hi1s1 U1693 ( .DIN(n1646), .Q(n1627) );
  hi1s1 U1694 ( .DIN(n1646), .Q(n1628) );
  hi1s1 U1695 ( .DIN(n1646), .Q(n1629) );
  hi1s1 U1696 ( .DIN(n1645), .Q(n1630) );
  hi1s1 U1697 ( .DIN(n1645), .Q(n1631) );
  hi1s1 U1698 ( .DIN(n1645), .Q(n1632) );
  hi1s1 U1699 ( .DIN(n1644), .Q(n1633) );
  hi1s1 U1700 ( .DIN(n1644), .Q(n1634) );
  hi1s1 U1701 ( .DIN(n1644), .Q(n1635) );
  hi1s1 U1702 ( .DIN(n15580), .Q(n1636) );
  hi1s1 U1703 ( .DIN(n1644), .Q(n1637) );
  hi1s1 U1704 ( .DIN(n1645), .Q(n1638) );
  hi1s1 U1705 ( .DIN(n1646), .Q(n1639) );
  hi1s1 U1706 ( .DIN(n1647), .Q(n1640) );
  hi1s1 U1707 ( .DIN(n1648), .Q(n1641) );
  hi1s1 U1708 ( .DIN(n1653), .Q(n1642) );
  hi1s1 U1709 ( .DIN(n1653), .Q(n1643) );
  hi1s1 U1710 ( .DIN(n1656), .Q(n1644) );
  hi1s1 U1711 ( .DIN(n1656), .Q(n1645) );
  hi1s1 U1712 ( .DIN(n1656), .Q(n1646) );
  hi1s1 U1713 ( .DIN(n1656), .Q(n1647) );
  hi1s1 U1714 ( .DIN(n1655), .Q(n1648) );
  hi1s1 U1715 ( .DIN(n1655), .Q(n1649) );
  hi1s1 U1716 ( .DIN(n1655), .Q(n1650) );
  hi1s1 U1717 ( .DIN(n1654), .Q(n1651) );
  hi1s1 U1718 ( .DIN(n1654), .Q(n1652) );
  hi1s1 U1719 ( .DIN(n1654), .Q(n1653) );
  hi1s1 U1720 ( .DIN(n15580), .Q(n1654) );
  hi1s1 U1721 ( .DIN(n15580), .Q(n1655) );
  hi1s1 U1722 ( .DIN(n15580), .Q(n1656) );
  nnd2s1 U1723 ( .DIN1(n1657), .DIN2(n1658), .Q(\u0/r0/N81 ) );
  or2s1 U1724 ( .DIN1(\u0/r0/N70 ), .DIN2(\u0/r0/n3 ), .Q(n1658) );
  and3s1 U1725 ( .DIN1(n1659), .DIN2(n1498), .DIN3(n1660), .Q(\u0/r0/N77 ) );
  and3s1 U1726 ( .DIN1(\u0/r0/rcnt[0]), .DIN2(n1659), .DIN3(n1660), 
        .Q(\u0/r0/N76 ) );
  nnd2s1 U1727 ( .DIN1(n1661), .DIN2(n1662), .Q(\u0/r0/N75 ) );
  nnd3s1 U1728 ( .DIN1(n1663), .DIN2(n1498), .DIN3(n1660), .Q(n1662) );
  hi1s1 U1729 ( .DIN(n1664), .Q(n1660) );
  nnd2s1 U1730 ( .DIN1(n1661), .DIN2(n1665), .Q(\u0/r0/N74 ) );
  nnd3s1 U1731 ( .DIN1(\u0/r0/rcnt[0]), .DIN2(n1666), .DIN3(n1663), 
        .Q(n1665) );
  nnd2s1 U1732 ( .DIN1(n1664), .DIN2(n1667), .Q(n1666) );
  nnd3s1 U1733 ( .DIN1(n1668), .DIN2(n1560), .DIN3(n1670), .Q(n1667) );
  nnd2s1 U1734 ( .DIN1(\u0/r0/N80 ), .DIN2(n1671), .Q(n1664) );
  nor2s1 U1735 ( .DIN1(n1670), .DIN2(ld), .Q(\u0/r0/N80 ) );
  and3s1 U1736 ( .DIN1(n1672), .DIN2(n1673), .DIN3(n1670), .Q(\u0/r0/N73 ) );
  nnd2s1 U1737 ( .DIN1(\u0/r0/rcnt[0]), .DIN2(n1674), .Q(n1673) );
  nnd3s1 U1738 ( .DIN1(n1663), .DIN2(n1560), .DIN3(n1668), .Q(n1674) );
  nnd2s1 U1739 ( .DIN1(n1675), .DIN2(n1498), .Q(n1672) );
  nnd2s1 U1740 ( .DIN1(\u0/r0/N79 ), .DIN2(n1671), .Q(n1675) );
  nnd2s1 U1741 ( .DIN1(n1661), .DIN2(n1676), .Q(\u0/r0/N72 ) );
  nnd4s1 U1742 ( .DIN1(n1670), .DIN2(\u0/r0/N79 ), .DIN3(\u0/r0/rcnt[0]), 
        .DIN4(n1671), .Q(n1676) );
  hi1s1 U1743 ( .DIN(n1668), .Q(n1671) );
  nor2s1 U1744 ( .DIN1(n1663), .DIN2(ld), .Q(\u0/r0/N79 ) );
  nnd4s1 U1745 ( .DIN1(n1670), .DIN2(\u0/r0/N78 ), .DIN3(n1668), .DIN4(n1663), 
        .Q(n1661) );
  xnr2s1 U1746 ( .DIN1(\u0/r0/n3 ), .DIN2(n1677), .Q(n1668) );
  nor2s1 U1747 ( .DIN1(n1419), .DIN2(n1678), .Q(n1677) );
  nor2s1 U1748 ( .DIN1(ld), .DIN2(\u0/r0/rcnt[0]), .Q(\u0/r0/N78 ) );
  xnr2s1 U1749 ( .DIN1(n1678), .DIN2(n1419), .Q(n1670) );
  nnd2s1 U1750 ( .DIN1(n1657), .DIN2(n1679), .Q(\u0/r0/N71 ) );
  or3s1 U1751 ( .DIN1(n1680), .DIN2(ld), .DIN3(n1681), .Q(n1679) );
  nnd4s1 U1752 ( .DIN1(\u0/r0/n3 ), .DIN2(n1680), .DIN3(n1681), .DIN4(n1560), 
        .Q(n1657) );
  nnd2s1 U1753 ( .DIN1(n1560), .DIN2(n1682), .Q(\u0/r0/N70 ) );
  nnd2s1 U1754 ( .DIN1(n1680), .DIN2(n1681), .Q(n1682) );
  nnd2s1 U1755 ( .DIN1(n1678), .DIN2(n1683), .Q(n1681) );
  nnd2s1 U1756 ( .DIN1(\u0/r0/rcnt[2]), .DIN2(n1659), .Q(n1683) );
  nnd2s1 U1757 ( .DIN1(\u0/r0/rcnt[0]), .DIN2(\u0/r0/rcnt[1]), .Q(n1678)
         );
  xor2s1 U1758 ( .DIN1(n1419), .DIN2(n1663), .Q(n1680) );
  hi1s1 U1759 ( .DIN(n1659), .Q(n1663) );
  xor2s1 U1760 ( .DIN1(\u0/r0/rcnt[1]), .DIN2(\u0/r0/rcnt[0]), .Q(n1659)
         );
  nnd2s1 U1761 ( .DIN1(n1684), .DIN2(n1685), .Q(\u0/N73 ) );
  nnd2s1 U1762 ( .DIN1(\key[127] ), .DIN2(ld), .Q(n1685) );
  or2s1 U1763 ( .DIN1(n1686), .DIN2(ld), .Q(n1684) );
  nnd2s1 U1764 ( .DIN1(n1687), .DIN2(n1688), .Q(\u0/N72 ) );
  nnd2s1 U1765 ( .DIN1(\key[126] ), .DIN2(ld), .Q(n1688) );
  or2s1 U1766 ( .DIN1(n1689), .DIN2(ld), .Q(n1687) );
  nnd2s1 U1767 ( .DIN1(n1690), .DIN2(n1691), .Q(\u0/N71 ) );
  nnd2s1 U1768 ( .DIN1(\key[125] ), .DIN2(ld), .Q(n1691) );
  or2s1 U1769 ( .DIN1(n1692), .DIN2(ld), .Q(n1690) );
  nnd2s1 U1770 ( .DIN1(n1693), .DIN2(n1694), .Q(\u0/N70 ) );
  nnd2s1 U1771 ( .DIN1(\key[124] ), .DIN2(ld), .Q(n1694) );
  or2s1 U1772 ( .DIN1(n1695), .DIN2(ld), .Q(n1693) );
  nnd2s1 U1773 ( .DIN1(n1696), .DIN2(n1697), .Q(\u0/N69 ) );
  nnd2s1 U1774 ( .DIN1(\key[123] ), .DIN2(ld), .Q(n1697) );
  or2s1 U1775 ( .DIN1(n1698), .DIN2(ld), .Q(n1696) );
  nnd2s1 U1776 ( .DIN1(n1699), .DIN2(n1700), .Q(\u0/N68 ) );
  nnd2s1 U1777 ( .DIN1(\key[122] ), .DIN2(ld), .Q(n1700) );
  or2s1 U1778 ( .DIN1(n1701), .DIN2(ld), .Q(n1699) );
  nnd2s1 U1779 ( .DIN1(n1702), .DIN2(n1703), .Q(\u0/N67 ) );
  nnd2s1 U1780 ( .DIN1(\key[121] ), .DIN2(ld), .Q(n1703) );
  or2s1 U1781 ( .DIN1(n1704), .DIN2(ld), .Q(n1702) );
  nnd2s1 U1782 ( .DIN1(n1705), .DIN2(n1706), .Q(\u0/N66 ) );
  nnd2s1 U1783 ( .DIN1(\key[120] ), .DIN2(ld), .Q(n1706) );
  or2s1 U1784 ( .DIN1(n1707), .DIN2(ld), .Q(n1705) );
  nnd2s1 U1785 ( .DIN1(n1708), .DIN2(n1709), .Q(\u0/N65 ) );
  nnd2s1 U1786 ( .DIN1(\key[119] ), .DIN2(ld), .Q(n1709) );
  or2s1 U1787 ( .DIN1(n1710), .DIN2(ld), .Q(n1708) );
  nnd2s1 U1788 ( .DIN1(n1711), .DIN2(n1712), .Q(\u0/N64 ) );
  nnd2s1 U1789 ( .DIN1(\key[118] ), .DIN2(ld), .Q(n1712) );
  or2s1 U1790 ( .DIN1(n1713), .DIN2(ld), .Q(n1711) );
  nnd2s1 U1791 ( .DIN1(n1714), .DIN2(n1715), .Q(\u0/N63 ) );
  nnd2s1 U1792 ( .DIN1(\key[117] ), .DIN2(ld), .Q(n1715) );
  or2s1 U1793 ( .DIN1(n1716), .DIN2(ld), .Q(n1714) );
  nnd2s1 U1794 ( .DIN1(n1717), .DIN2(n1718), .Q(\u0/N62 ) );
  nnd2s1 U1795 ( .DIN1(\key[116] ), .DIN2(ld), .Q(n1718) );
  or2s1 U1796 ( .DIN1(n1719), .DIN2(ld), .Q(n1717) );
  nnd2s1 U1797 ( .DIN1(n1720), .DIN2(n1721), .Q(\u0/N61 ) );
  nnd2s1 U1798 ( .DIN1(\key[115] ), .DIN2(ld), .Q(n1721) );
  or2s1 U1799 ( .DIN1(n1722), .DIN2(ld), .Q(n1720) );
  nnd2s1 U1800 ( .DIN1(n1723), .DIN2(n1724), .Q(\u0/N60 ) );
  nnd2s1 U1801 ( .DIN1(\key[114] ), .DIN2(ld), .Q(n1724) );
  or2s1 U1802 ( .DIN1(n1725), .DIN2(ld), .Q(n1723) );
  nnd2s1 U1803 ( .DIN1(n1726), .DIN2(n1727), .Q(\u0/N59 ) );
  nnd2s1 U1804 ( .DIN1(\key[113] ), .DIN2(ld), .Q(n1727) );
  or2s1 U1805 ( .DIN1(n1728), .DIN2(ld), .Q(n1726) );
  nnd2s1 U1806 ( .DIN1(n1729), .DIN2(n1730), .Q(\u0/N58 ) );
  nnd2s1 U1807 ( .DIN1(\key[112] ), .DIN2(ld), .Q(n1730) );
  or2s1 U1808 ( .DIN1(n1731), .DIN2(ld), .Q(n1729) );
  nnd2s1 U1809 ( .DIN1(n1732), .DIN2(n1733), .Q(\u0/N57 ) );
  nnd2s1 U1810 ( .DIN1(\key[111] ), .DIN2(ld), .Q(n1733) );
  or2s1 U1811 ( .DIN1(n1734), .DIN2(ld), .Q(n1732) );
  nnd2s1 U1812 ( .DIN1(n1735), .DIN2(n1736), .Q(\u0/N56 ) );
  nnd2s1 U1813 ( .DIN1(\key[110] ), .DIN2(ld), .Q(n1736) );
  or2s1 U1814 ( .DIN1(n1737), .DIN2(ld), .Q(n1735) );
  nnd2s1 U1815 ( .DIN1(n1738), .DIN2(n1739), .Q(\u0/N55 ) );
  nnd2s1 U1816 ( .DIN1(\key[109] ), .DIN2(ld), .Q(n1739) );
  or2s1 U1817 ( .DIN1(n1740), .DIN2(ld), .Q(n1738) );
  nnd2s1 U1818 ( .DIN1(n1741), .DIN2(n1742), .Q(\u0/N54 ) );
  nnd2s1 U1819 ( .DIN1(\key[108] ), .DIN2(ld), .Q(n1742) );
  or2s1 U1820 ( .DIN1(n1743), .DIN2(ld), .Q(n1741) );
  nnd2s1 U1821 ( .DIN1(n1744), .DIN2(n1745), .Q(\u0/N53 ) );
  nnd2s1 U1822 ( .DIN1(\key[107] ), .DIN2(ld), .Q(n1745) );
  or2s1 U1823 ( .DIN1(n1746), .DIN2(ld), .Q(n1744) );
  nnd2s1 U1824 ( .DIN1(n1747), .DIN2(n1748), .Q(\u0/N52 ) );
  nnd2s1 U1825 ( .DIN1(\key[106] ), .DIN2(ld), .Q(n1748) );
  or2s1 U1826 ( .DIN1(n1749), .DIN2(ld), .Q(n1747) );
  nnd2s1 U1827 ( .DIN1(n1750), .DIN2(n1751), .Q(\u0/N51 ) );
  nnd2s1 U1828 ( .DIN1(\key[105] ), .DIN2(ld), .Q(n1751) );
  or2s1 U1829 ( .DIN1(n1752), .DIN2(ld), .Q(n1750) );
  nnd2s1 U1830 ( .DIN1(n1753), .DIN2(n1754), .Q(\u0/N50 ) );
  nnd2s1 U1831 ( .DIN1(\key[104] ), .DIN2(ld), .Q(n1754) );
  or2s1 U1832 ( .DIN1(n1755), .DIN2(ld), .Q(n1753) );
  nnd2s1 U1833 ( .DIN1(n1756), .DIN2(n1757), .Q(\u0/N49 ) );
  nnd2s1 U1834 ( .DIN1(\key[103] ), .DIN2(ld), .Q(n1757) );
  or2s1 U1835 ( .DIN1(n1758), .DIN2(ld), .Q(n1756) );
  nnd2s1 U1836 ( .DIN1(n1759), .DIN2(n1760), .Q(\u0/N48 ) );
  nnd2s1 U1837 ( .DIN1(\key[102] ), .DIN2(ld), .Q(n1760) );
  or2s1 U1838 ( .DIN1(n1761), .DIN2(ld), .Q(n1759) );
  nnd2s1 U1839 ( .DIN1(n1762), .DIN2(n1763), .Q(\u0/N47 ) );
  nnd2s1 U1840 ( .DIN1(\key[101] ), .DIN2(ld), .Q(n1763) );
  or2s1 U1841 ( .DIN1(n1764), .DIN2(ld), .Q(n1762) );
  nnd2s1 U1842 ( .DIN1(n1765), .DIN2(n1766), .Q(\u0/N46 ) );
  nnd2s1 U1843 ( .DIN1(\key[100] ), .DIN2(ld), .Q(n1766) );
  or2s1 U1844 ( .DIN1(n1767), .DIN2(ld), .Q(n1765) );
  nnd2s1 U1845 ( .DIN1(n1768), .DIN2(n1769), .Q(\u0/N45 ) );
  nnd2s1 U1846 ( .DIN1(\key[99] ), .DIN2(ld), .Q(n1769) );
  or2s1 U1847 ( .DIN1(n1770), .DIN2(ld), .Q(n1768) );
  nnd2s1 U1848 ( .DIN1(n1771), .DIN2(n1772), .Q(\u0/N44 ) );
  nnd2s1 U1849 ( .DIN1(\key[98] ), .DIN2(ld), .Q(n1772) );
  or2s1 U1850 ( .DIN1(n1773), .DIN2(ld), .Q(n1771) );
  nnd2s1 U1851 ( .DIN1(n1774), .DIN2(n1775), .Q(\u0/N43 ) );
  nnd2s1 U1852 ( .DIN1(\key[97] ), .DIN2(ld), .Q(n1775) );
  or2s1 U1853 ( .DIN1(n1776), .DIN2(ld), .Q(n1774) );
  nnd2s1 U1854 ( .DIN1(n1777), .DIN2(n1778), .Q(\u0/N42 ) );
  nnd2s1 U1855 ( .DIN1(\key[96] ), .DIN2(ld), .Q(n1778) );
  or2s1 U1856 ( .DIN1(n1779), .DIN2(ld), .Q(n1777) );
  nnd2s1 U1857 ( .DIN1(n1780), .DIN2(n1781), .Q(\u0/N271 ) );
  nnd2s1 U1858 ( .DIN1(\key[31] ), .DIN2(ld), .Q(n1781) );
  nnd2s1 U1859 ( .DIN1(n1782), .DIN2(n1561), .Q(n1780) );
  xor2s1 U1860 ( .DIN1(n1416), .DIN2(n1783), .Q(n1782) );
  nnd2s1 U1861 ( .DIN1(n1784), .DIN2(n1785), .Q(\u0/N270 ) );
  nnd2s1 U1862 ( .DIN1(\key[30] ), .DIN2(ld), .Q(n1785) );
  nnd2s1 U1863 ( .DIN1(n1786), .DIN2(n1561), .Q(n1784) );
  xor2s1 U1864 ( .DIN1(n1475), .DIN2(n1787), .Q(n1786) );
  nnd2s1 U1865 ( .DIN1(n1788), .DIN2(n1789), .Q(\u0/N269 ) );
  nnd2s1 U1866 ( .DIN1(\key[29] ), .DIN2(ld), .Q(n1789) );
  nnd2s1 U1867 ( .DIN1(n1790), .DIN2(n1561), .Q(n1788) );
  xor2s1 U1868 ( .DIN1(n1374), .DIN2(n1791), .Q(n1790) );
  nnd2s1 U1869 ( .DIN1(n1792), .DIN2(n1793), .Q(\u0/N268 ) );
  nnd2s1 U1870 ( .DIN1(\key[28] ), .DIN2(ld), .Q(n1793) );
  nnd2s1 U1871 ( .DIN1(n1794), .DIN2(n1561), .Q(n1792) );
  xor2s1 U1872 ( .DIN1(n1392), .DIN2(n1795), .Q(n1794) );
  nnd2s1 U1873 ( .DIN1(n1796), .DIN2(n1797), .Q(\u0/N267 ) );
  nnd2s1 U1874 ( .DIN1(\key[27] ), .DIN2(ld), .Q(n1797) );
  nnd2s1 U1875 ( .DIN1(n1798), .DIN2(n1561), .Q(n1796) );
  xor2s1 U1876 ( .DIN1(n1476), .DIN2(n1799), .Q(n1798) );
  nnd2s1 U1877 ( .DIN1(n1800), .DIN2(n1801), .Q(\u0/N266 ) );
  nnd2s1 U1878 ( .DIN1(\key[26] ), .DIN2(ld), .Q(n1801) );
  nnd2s1 U1879 ( .DIN1(n1802), .DIN2(n1561), .Q(n1800) );
  xor2s1 U1880 ( .DIN1(n1548), .DIN2(n1803), .Q(n1802) );
  nnd2s1 U1881 ( .DIN1(n1804), .DIN2(n1805), .Q(\u0/N265 ) );
  nnd2s1 U1882 ( .DIN1(\key[25] ), .DIN2(ld), .Q(n1805) );
  nnd2s1 U1883 ( .DIN1(n1806), .DIN2(n1561), .Q(n1804) );
  xor2s1 U1884 ( .DIN1(n1410), .DIN2(n1807), .Q(n1806) );
  nnd2s1 U1885 ( .DIN1(n1808), .DIN2(n1809), .Q(\u0/N264 ) );
  nnd2s1 U1886 ( .DIN1(\key[24] ), .DIN2(ld), .Q(n1809) );
  nnd2s1 U1887 ( .DIN1(n1810), .DIN2(n1562), .Q(n1808) );
  xor2s1 U1888 ( .DIN1(n1554), .DIN2(n1811), .Q(n1810) );
  nnd2s1 U1889 ( .DIN1(n1812), .DIN2(n1813), .Q(\u0/N263 ) );
  nnd2s1 U1890 ( .DIN1(\key[23] ), .DIN2(ld), .Q(n1813) );
  nnd2s1 U1891 ( .DIN1(n1814), .DIN2(n1562), .Q(n1812) );
  xor2s1 U1892 ( .DIN1(n1415), .DIN2(n1815), .Q(n1814) );
  nnd2s1 U1893 ( .DIN1(n1816), .DIN2(n1817), .Q(\u0/N262 ) );
  nnd2s1 U1894 ( .DIN1(\key[22] ), .DIN2(ld), .Q(n1817) );
  nnd2s1 U1895 ( .DIN1(n1818), .DIN2(n1562), .Q(n1816) );
  xor2s1 U1896 ( .DIN1(n1438), .DIN2(n1819), .Q(n1818) );
  nnd2s1 U1897 ( .DIN1(n1820), .DIN2(n1821), .Q(\u0/N261 ) );
  nnd2s1 U1898 ( .DIN1(\key[21] ), .DIN2(ld), .Q(n1821) );
  nnd2s1 U1899 ( .DIN1(n1822), .DIN2(n1562), .Q(n1820) );
  xor2s1 U1900 ( .DIN1(n1373), .DIN2(n1823), .Q(n1822) );
  nnd2s1 U1901 ( .DIN1(n1824), .DIN2(n1825), .Q(\u0/N260 ) );
  nnd2s1 U1902 ( .DIN1(\key[20] ), .DIN2(ld), .Q(n1825) );
  nnd2s1 U1903 ( .DIN1(n1826), .DIN2(n1562), .Q(n1824) );
  xor2s1 U1904 ( .DIN1(n1376), .DIN2(n1827), .Q(n1826) );
  nnd2s1 U1905 ( .DIN1(n1828), .DIN2(n1829), .Q(\u0/N259 ) );
  nnd2s1 U1906 ( .DIN1(\key[19] ), .DIN2(ld), .Q(n1829) );
  nnd2s1 U1907 ( .DIN1(n1830), .DIN2(n1562), .Q(n1828) );
  xor2s1 U1908 ( .DIN1(n1439), .DIN2(n1831), .Q(n1830) );
  nnd2s1 U1909 ( .DIN1(n1832), .DIN2(n1833), .Q(\u0/N258 ) );
  nnd2s1 U1910 ( .DIN1(\key[18] ), .DIN2(ld), .Q(n1833) );
  nnd2s1 U1911 ( .DIN1(n1834), .DIN2(n1562), .Q(n1832) );
  xor2s1 U1912 ( .DIN1(n1368), .DIN2(n1835), .Q(n1834) );
  nnd2s1 U1913 ( .DIN1(n1836), .DIN2(n1837), .Q(\u0/N257 ) );
  nnd2s1 U1914 ( .DIN1(\key[17] ), .DIN2(ld), .Q(n1837) );
  nnd2s1 U1915 ( .DIN1(n1838), .DIN2(n1563), .Q(n1836) );
  xor2s1 U1916 ( .DIN1(n1412), .DIN2(n1839), .Q(n1838) );
  nnd2s1 U1917 ( .DIN1(n1840), .DIN2(n1841), .Q(\u0/N256 ) );
  nnd2s1 U1918 ( .DIN1(\key[16] ), .DIN2(ld), .Q(n1841) );
  nnd2s1 U1919 ( .DIN1(n1842), .DIN2(n1563), .Q(n1840) );
  xor2s1 U1920 ( .DIN1(n1558), .DIN2(n1843), .Q(n1842) );
  nnd2s1 U1921 ( .DIN1(n1844), .DIN2(n1845), .Q(\u0/N255 ) );
  nnd2s1 U1922 ( .DIN1(\key[15] ), .DIN2(ld), .Q(n1845) );
  nnd2s1 U1923 ( .DIN1(n1846), .DIN2(n1563), .Q(n1844) );
  xor2s1 U1924 ( .DIN1(n1414), .DIN2(n1847), .Q(n1846) );
  nnd2s1 U1925 ( .DIN1(n1848), .DIN2(n1849), .Q(\u0/N254 ) );
  nnd2s1 U1926 ( .DIN1(\key[14] ), .DIN2(ld), .Q(n1849) );
  nnd2s1 U1927 ( .DIN1(n1850), .DIN2(n1563), .Q(n1848) );
  xor2s1 U1928 ( .DIN1(n1474), .DIN2(n1851), .Q(n1850) );
  nnd2s1 U1929 ( .DIN1(n1852), .DIN2(n1853), .Q(\u0/N253 ) );
  nnd2s1 U1930 ( .DIN1(\key[13] ), .DIN2(ld), .Q(n1853) );
  nnd2s1 U1931 ( .DIN1(n1854), .DIN2(n1563), .Q(n1852) );
  xor2s1 U1932 ( .DIN1(n1372), .DIN2(n1855), .Q(n1854) );
  nnd2s1 U1933 ( .DIN1(n1856), .DIN2(n1857), .Q(\u0/N252 ) );
  nnd2s1 U1934 ( .DIN1(\key[12] ), .DIN2(ld), .Q(n1857) );
  nnd2s1 U1935 ( .DIN1(n1858), .DIN2(n1563), .Q(n1856) );
  xor2s1 U1936 ( .DIN1(n1393), .DIN2(n1859), .Q(n1858) );
  nnd2s1 U1937 ( .DIN1(n1860), .DIN2(n1861), .Q(\u0/N251 ) );
  nnd2s1 U1938 ( .DIN1(\key[11] ), .DIN2(ld), .Q(n1861) );
  nnd2s1 U1939 ( .DIN1(n1862), .DIN2(n1563), .Q(n1860) );
  xor2s1 U1940 ( .DIN1(n1413), .DIN2(n1863), .Q(n1862) );
  nnd2s1 U1941 ( .DIN1(n1864), .DIN2(n1865), .Q(\u0/N250 ) );
  nnd2s1 U1942 ( .DIN1(\key[10] ), .DIN2(ld), .Q(n1865) );
  nnd2s1 U1943 ( .DIN1(n1866), .DIN2(n1564), .Q(n1864) );
  xor2s1 U1944 ( .DIN1(n1553), .DIN2(n1867), .Q(n1866) );
  nnd2s1 U1945 ( .DIN1(n1868), .DIN2(n1869), .Q(\u0/N249 ) );
  nnd2s1 U1946 ( .DIN1(\key[9] ), .DIN2(ld), .Q(n1869) );
  nnd2s1 U1947 ( .DIN1(n1870), .DIN2(n1564), .Q(n1868) );
  xor2s1 U1948 ( .DIN1(n1547), .DIN2(n1871), .Q(n1870) );
  nnd2s1 U1949 ( .DIN1(n1872), .DIN2(n1873), .Q(\u0/N248 ) );
  nnd2s1 U1950 ( .DIN1(\key[8] ), .DIN2(ld), .Q(n1873) );
  nnd2s1 U1951 ( .DIN1(n1874), .DIN2(n1564), .Q(n1872) );
  xor2s1 U1952 ( .DIN1(n1361), .DIN2(n1875), .Q(n1874) );
  nnd2s1 U1953 ( .DIN1(n1876), .DIN2(n1877), .Q(\u0/N247 ) );
  nnd2s1 U1954 ( .DIN1(\key[7] ), .DIN2(ld), .Q(n1877) );
  nnd2s1 U1955 ( .DIN1(n1878), .DIN2(n1564), .Q(n1876) );
  xor2s1 U1956 ( .DIN1(n1442), .DIN2(n1879), .Q(n1878) );
  nnd2s1 U1957 ( .DIN1(n1880), .DIN2(n1881), .Q(\u0/N246 ) );
  nnd2s1 U1958 ( .DIN1(\key[6] ), .DIN2(ld), .Q(n1881) );
  nnd2s1 U1959 ( .DIN1(n1882), .DIN2(n1564), .Q(n1880) );
  xor2s1 U1960 ( .DIN1(n1391), .DIN2(n1883), .Q(n1882) );
  nnd2s1 U1961 ( .DIN1(n1884), .DIN2(n1885), .Q(\u0/N245 ) );
  nnd2s1 U1962 ( .DIN1(\key[5] ), .DIN2(ld), .Q(n1885) );
  nnd2s1 U1963 ( .DIN1(n1886), .DIN2(n1564), .Q(n1884) );
  xor2s1 U1964 ( .DIN1(n1375), .DIN2(n1887), .Q(n1886) );
  nnd2s1 U1965 ( .DIN1(n1888), .DIN2(n1889), .Q(\u0/N244 ) );
  nnd2s1 U1966 ( .DIN1(\key[4] ), .DIN2(ld), .Q(n1889) );
  nnd2s1 U1967 ( .DIN1(n1890), .DIN2(n1564), .Q(n1888) );
  xor2s1 U1968 ( .DIN1(n1441), .DIN2(n1891), .Q(n1890) );
  nnd2s1 U1969 ( .DIN1(n1892), .DIN2(n1893), .Q(\u0/N243 ) );
  nnd2s1 U1970 ( .DIN1(\key[3] ), .DIN2(ld), .Q(n1893) );
  nnd2s1 U1971 ( .DIN1(n1894), .DIN2(n1565), .Q(n1892) );
  xor2s1 U1972 ( .DIN1(n1440), .DIN2(n1895), .Q(n1894) );
  nnd2s1 U1973 ( .DIN1(n1896), .DIN2(n1897), .Q(\u0/N242 ) );
  nnd2s1 U1974 ( .DIN1(\key[2] ), .DIN2(ld), .Q(n1897) );
  nnd2s1 U1975 ( .DIN1(n1898), .DIN2(n1565), .Q(n1896) );
  xor2s1 U1976 ( .DIN1(n1369), .DIN2(n1899), .Q(n1898) );
  nnd2s1 U1977 ( .DIN1(n1900), .DIN2(n1901), .Q(\u0/N241 ) );
  nnd2s1 U1978 ( .DIN1(\key[1] ), .DIN2(ld), .Q(n1901) );
  nnd2s1 U1979 ( .DIN1(n1902), .DIN2(n1565), .Q(n1900) );
  xor2s1 U1980 ( .DIN1(n1411), .DIN2(n1903), .Q(n1902) );
  nnd2s1 U1981 ( .DIN1(n1904), .DIN2(n1905), .Q(\u0/N240 ) );
  nnd2s1 U1982 ( .DIN1(\key[0] ), .DIN2(ld), .Q(n1905) );
  nnd2s1 U1983 ( .DIN1(n1906), .DIN2(n1565), .Q(n1904) );
  xor2s1 U1984 ( .DIN1(n1556), .DIN2(n1907), .Q(n1906) );
  nnd2s1 U1985 ( .DIN1(n1908), .DIN2(n1909), .Q(\u0/N205 ) );
  nnd2s1 U1986 ( .DIN1(\key[63] ), .DIN2(ld), .Q(n1909) );
  or2s1 U1987 ( .DIN1(n1783), .DIN2(ld), .Q(n1908) );
  xor2s1 U1988 ( .DIN1(n1451), .DIN2(n1910), .Q(n1783) );
  nnd2s1 U1989 ( .DIN1(n1911), .DIN2(n1912), .Q(\u0/N204 ) );
  nnd2s1 U1990 ( .DIN1(\key[62] ), .DIN2(ld), .Q(n1912) );
  or2s1 U1991 ( .DIN1(n1787), .DIN2(ld), .Q(n1911) );
  xnr2s1 U1992 ( .DIN1(w2[30]), .DIN2(n1913), .Q(n1787) );
  nnd2s1 U1993 ( .DIN1(n1914), .DIN2(n1915), .Q(\u0/N203 ) );
  nnd2s1 U1994 ( .DIN1(\key[61] ), .DIN2(ld), .Q(n1915) );
  or2s1 U1995 ( .DIN1(n1791), .DIN2(ld), .Q(n1914) );
  xor2s1 U1996 ( .DIN1(n1452), .DIN2(n1916), .Q(n1791) );
  nnd2s1 U1997 ( .DIN1(n1917), .DIN2(n1918), .Q(\u0/N202 ) );
  nnd2s1 U1998 ( .DIN1(\key[60] ), .DIN2(ld), .Q(n1918) );
  or2s1 U1999 ( .DIN1(n1795), .DIN2(ld), .Q(n1917) );
  xor2s1 U2000 ( .DIN1(n1477), .DIN2(n1919), .Q(n1795) );
  nnd2s1 U2001 ( .DIN1(n1920), .DIN2(n1921), .Q(\u0/N201 ) );
  nnd2s1 U2002 ( .DIN1(\key[59] ), .DIN2(ld), .Q(n1921) );
  or2s1 U2003 ( .DIN1(n1799), .DIN2(ld), .Q(n1920) );
  xnr2s1 U2004 ( .DIN1(w2[27]), .DIN2(n1922), .Q(n1799) );
  nnd2s1 U2005 ( .DIN1(n1923), .DIN2(n1924), .Q(\u0/N200 ) );
  nnd2s1 U2006 ( .DIN1(\key[58] ), .DIN2(ld), .Q(n1924) );
  or2s1 U2007 ( .DIN1(n1803), .DIN2(ld), .Q(n1923) );
  xor2s1 U2008 ( .DIN1(n1453), .DIN2(n1925), .Q(n1803) );
  nnd2s1 U2009 ( .DIN1(n1926), .DIN2(n1927), .Q(\u0/N199 ) );
  nnd2s1 U2010 ( .DIN1(\key[57] ), .DIN2(ld), .Q(n1927) );
  or2s1 U2011 ( .DIN1(n1807), .DIN2(ld), .Q(n1926) );
  xnr2s1 U2012 ( .DIN1(w2[25]), .DIN2(n1928), .Q(n1807) );
  nnd2s1 U2013 ( .DIN1(n1929), .DIN2(n1930), .Q(\u0/N198 ) );
  nnd2s1 U2014 ( .DIN1(\key[56] ), .DIN2(ld), .Q(n1930) );
  or2s1 U2015 ( .DIN1(n1811), .DIN2(ld), .Q(n1929) );
  xor2s1 U2016 ( .DIN1(n1454), .DIN2(n1931), .Q(n1811) );
  nnd2s1 U2017 ( .DIN1(n1932), .DIN2(n1933), .Q(\u0/N197 ) );
  nnd2s1 U2018 ( .DIN1(\key[55] ), .DIN2(ld), .Q(n1933) );
  or2s1 U2019 ( .DIN1(n1815), .DIN2(ld), .Q(n1932) );
  xnr2s1 U2020 ( .DIN1(w2[23]), .DIN2(n1934), .Q(n1815) );
  nnd2s1 U2021 ( .DIN1(n1935), .DIN2(n1936), .Q(\u0/N196 ) );
  nnd2s1 U2022 ( .DIN1(\key[54] ), .DIN2(ld), .Q(n1936) );
  or2s1 U2023 ( .DIN1(n1819), .DIN2(ld), .Q(n1935) );
  xor2s1 U2024 ( .DIN1(n1482), .DIN2(n1937), .Q(n1819) );
  nnd2s1 U2025 ( .DIN1(n1938), .DIN2(n1939), .Q(\u0/N195 ) );
  nnd2s1 U2026 ( .DIN1(\key[53] ), .DIN2(ld), .Q(n1939) );
  or2s1 U2027 ( .DIN1(n1823), .DIN2(ld), .Q(n1938) );
  xnr2s1 U2028 ( .DIN1(w2[21]), .DIN2(n1940), .Q(n1823) );
  nnd2s1 U2029 ( .DIN1(n1941), .DIN2(n1942), .Q(\u0/N194 ) );
  nnd2s1 U2030 ( .DIN1(\key[52] ), .DIN2(ld), .Q(n1942) );
  or2s1 U2031 ( .DIN1(n1827), .DIN2(ld), .Q(n1941) );
  xor2s1 U2032 ( .DIN1(n1455), .DIN2(n1943), .Q(n1827) );
  nnd2s1 U2033 ( .DIN1(n1944), .DIN2(n1945), .Q(\u0/N193 ) );
  nnd2s1 U2034 ( .DIN1(\key[51] ), .DIN2(ld), .Q(n1945) );
  or2s1 U2035 ( .DIN1(n1831), .DIN2(ld), .Q(n1944) );
  xor2s1 U2036 ( .DIN1(n1483), .DIN2(n1946), .Q(n1831) );
  nnd2s1 U2037 ( .DIN1(n1947), .DIN2(n1948), .Q(\u0/N192 ) );
  nnd2s1 U2038 ( .DIN1(\key[50] ), .DIN2(ld), .Q(n1948) );
  or2s1 U2039 ( .DIN1(n1835), .DIN2(ld), .Q(n1947) );
  xnr2s1 U2040 ( .DIN1(w2[18]), .DIN2(n1949), .Q(n1835) );
  nnd2s1 U2041 ( .DIN1(n1950), .DIN2(n1951), .Q(\u0/N191 ) );
  nnd2s1 U2042 ( .DIN1(\key[49] ), .DIN2(ld), .Q(n1951) );
  or2s1 U2043 ( .DIN1(n1839), .DIN2(ld), .Q(n1950) );
  xor2s1 U2044 ( .DIN1(n1456), .DIN2(n1952), .Q(n1839) );
  nnd2s1 U2045 ( .DIN1(n1953), .DIN2(n1954), .Q(\u0/N190 ) );
  nnd2s1 U2046 ( .DIN1(\key[48] ), .DIN2(ld), .Q(n1954) );
  or2s1 U2047 ( .DIN1(n1843), .DIN2(ld), .Q(n1953) );
  xor2s1 U2048 ( .DIN1(n1457), .DIN2(n1955), .Q(n1843) );
  nnd2s1 U2049 ( .DIN1(n1956), .DIN2(n1957), .Q(\u0/N189 ) );
  nnd2s1 U2050 ( .DIN1(\key[47] ), .DIN2(ld), .Q(n1957) );
  or2s1 U2051 ( .DIN1(n1847), .DIN2(ld), .Q(n1956) );
  xor2s1 U2052 ( .DIN1(n1458), .DIN2(n1958), .Q(n1847) );
  nnd2s1 U2053 ( .DIN1(n1959), .DIN2(n1960), .Q(\u0/N188 ) );
  nnd2s1 U2054 ( .DIN1(\key[46] ), .DIN2(ld), .Q(n1960) );
  or2s1 U2055 ( .DIN1(n1851), .DIN2(ld), .Q(n1959) );
  xnr2s1 U2056 ( .DIN1(w2[14]), .DIN2(n1961), .Q(n1851) );
  nnd2s1 U2057 ( .DIN1(n1962), .DIN2(n1963), .Q(\u0/N187 ) );
  nnd2s1 U2058 ( .DIN1(\key[45] ), .DIN2(ld), .Q(n1963) );
  or2s1 U2059 ( .DIN1(n1855), .DIN2(ld), .Q(n1962) );
  xor2s1 U2060 ( .DIN1(n1459), .DIN2(n1964), .Q(n1855) );
  nnd2s1 U2061 ( .DIN1(n1965), .DIN2(n1966), .Q(\u0/N186 ) );
  nnd2s1 U2062 ( .DIN1(\key[44] ), .DIN2(ld), .Q(n1966) );
  or2s1 U2063 ( .DIN1(n1859), .DIN2(ld), .Q(n1965) );
  xor2s1 U2064 ( .DIN1(n1460), .DIN2(n1967), .Q(n1859) );
  nnd2s1 U2065 ( .DIN1(n1968), .DIN2(n1969), .Q(\u0/N185 ) );
  nnd2s1 U2066 ( .DIN1(\key[43] ), .DIN2(ld), .Q(n1969) );
  or2s1 U2067 ( .DIN1(n1863), .DIN2(ld), .Q(n1968) );
  xnr2s1 U2068 ( .DIN1(w2[11]), .DIN2(n1970), .Q(n1863) );
  nnd2s1 U2069 ( .DIN1(n1971), .DIN2(n1972), .Q(\u0/N184 ) );
  nnd2s1 U2070 ( .DIN1(\key[42] ), .DIN2(ld), .Q(n1972) );
  or2s1 U2071 ( .DIN1(n1867), .DIN2(ld), .Q(n1971) );
  xnr2s1 U2072 ( .DIN1(w2[10]), .DIN2(n1973), .Q(n1867) );
  nnd2s1 U2073 ( .DIN1(n1974), .DIN2(n1975), .Q(\u0/N183 ) );
  nnd2s1 U2074 ( .DIN1(\key[41] ), .DIN2(ld), .Q(n1975) );
  or2s1 U2075 ( .DIN1(n1871), .DIN2(ld), .Q(n1974) );
  xnr2s1 U2076 ( .DIN1(w2[9]), .DIN2(n1976), .Q(n1871) );
  nnd2s1 U2077 ( .DIN1(n1977), .DIN2(n1978), .Q(\u0/N182 ) );
  nnd2s1 U2078 ( .DIN1(\key[40] ), .DIN2(ld), .Q(n1978) );
  or2s1 U2079 ( .DIN1(n1875), .DIN2(ld), .Q(n1977) );
  xor2s1 U2080 ( .DIN1(n1461), .DIN2(n1979), .Q(n1875) );
  nnd2s1 U2081 ( .DIN1(n1980), .DIN2(n1981), .Q(\u0/N181 ) );
  nnd2s1 U2082 ( .DIN1(\key[39] ), .DIN2(ld), .Q(n1981) );
  or2s1 U2083 ( .DIN1(n1879), .DIN2(ld), .Q(n1980) );
  xnr2s1 U2084 ( .DIN1(w2[7]), .DIN2(n1982), .Q(n1879) );
  nnd2s1 U2085 ( .DIN1(n1983), .DIN2(n1984), .Q(\u0/N180 ) );
  nnd2s1 U2086 ( .DIN1(\key[38] ), .DIN2(ld), .Q(n1984) );
  or2s1 U2087 ( .DIN1(n1883), .DIN2(ld), .Q(n1983) );
  xnr2s1 U2088 ( .DIN1(w2[6]), .DIN2(n1985), .Q(n1883) );
  nnd2s1 U2089 ( .DIN1(n1986), .DIN2(n1987), .Q(\u0/N179 ) );
  nnd2s1 U2090 ( .DIN1(\key[37] ), .DIN2(ld), .Q(n1987) );
  or2s1 U2091 ( .DIN1(n1887), .DIN2(ld), .Q(n1986) );
  xor2s1 U2092 ( .DIN1(n1462), .DIN2(n1988), .Q(n1887) );
  nnd2s1 U2093 ( .DIN1(n1989), .DIN2(n1990), .Q(\u0/N178 ) );
  nnd2s1 U2094 ( .DIN1(\key[36] ), .DIN2(ld), .Q(n1990) );
  or2s1 U2095 ( .DIN1(n1891), .DIN2(ld), .Q(n1989) );
  xor2s1 U2096 ( .DIN1(n1478), .DIN2(n1991), .Q(n1891) );
  nnd2s1 U2097 ( .DIN1(n1992), .DIN2(n1993), .Q(\u0/N177 ) );
  nnd2s1 U2098 ( .DIN1(\key[35] ), .DIN2(ld), .Q(n1993) );
  or2s1 U2099 ( .DIN1(n1895), .DIN2(ld), .Q(n1992) );
  xor2s1 U2100 ( .DIN1(n1484), .DIN2(n1994), .Q(n1895) );
  nnd2s1 U2101 ( .DIN1(n1995), .DIN2(n1996), .Q(\u0/N176 ) );
  nnd2s1 U2102 ( .DIN1(\key[34] ), .DIN2(ld), .Q(n1996) );
  or2s1 U2103 ( .DIN1(n1899), .DIN2(ld), .Q(n1995) );
  xnr2s1 U2104 ( .DIN1(w2[2]), .DIN2(n1997), .Q(n1899) );
  nnd2s1 U2105 ( .DIN1(n1998), .DIN2(n1999), .Q(\u0/N175 ) );
  nnd2s1 U2106 ( .DIN1(\key[33] ), .DIN2(ld), .Q(n1999) );
  or2s1 U2107 ( .DIN1(n1903), .DIN2(ld), .Q(n1998) );
  xor2s1 U2108 ( .DIN1(n1479), .DIN2(n2000), .Q(n1903) );
  nnd2s1 U2109 ( .DIN1(n2001), .DIN2(n2002), .Q(\u0/N174 ) );
  nnd2s1 U2110 ( .DIN1(\key[32] ), .DIN2(ld), .Q(n2002) );
  or2s1 U2111 ( .DIN1(n1907), .DIN2(ld), .Q(n2001) );
  xor2s1 U2112 ( .DIN1(n1450), .DIN2(n2003), .Q(n1907) );
  nnd2s1 U2113 ( .DIN1(n2004), .DIN2(n2005), .Q(\u0/N139 ) );
  nnd2s1 U2114 ( .DIN1(\key[95] ), .DIN2(ld), .Q(n2005) );
  nnd2s1 U2115 ( .DIN1(n1910), .DIN2(n1565), .Q(n2004) );
  xnr2s1 U2116 ( .DIN1(w1[31]), .DIN2(n1686), .Q(n1910) );
  xnr2s1 U2117 ( .DIN1(n2006), .DIN2(n2007), .Q(n1686) );
  nor4s1 U2118 ( .DIN1(n2008), .DIN2(n2009), .DIN3(n2010), .DIN4(n2011), 
        .Q(n2007) );
  nnd3s1 U2119 ( .DIN1(n2012), .DIN2(n2013), .DIN3(n2014), .Q(n2011) );
  nnd4s1 U2120 ( .DIN1(n2015), .DIN2(n2016), .DIN3(n2017), .DIN4(n2018), 
        .Q(n2010) );
  nnd2s1 U2121 ( .DIN1(n2019), .DIN2(n2020), .Q(n2017) );
  nnd2s1 U2122 ( .DIN1(n2021), .DIN2(n2022), .Q(n2016) );
  nnd4s1 U2123 ( .DIN1(n2023), .DIN2(n2024), .DIN3(n2025), .DIN4(n2026), 
        .Q(n2009) );
  nnd2s1 U2124 ( .DIN1(n2027), .DIN2(n2028), .Q(n2026) );
  nnd2s1 U2125 ( .DIN1(n2029), .DIN2(n2030), .Q(n2025) );
  nnd2s1 U2126 ( .DIN1(n2031), .DIN2(n2032), .Q(n2024) );
  nnd4s1 U2127 ( .DIN1(n2033), .DIN2(n2034), .DIN3(n2035), .DIN4(n2036), 
        .Q(n2008) );
  nnd2s1 U2128 ( .DIN1(n2037), .DIN2(n2038), .Q(n2036) );
  nnd2s1 U2129 ( .DIN1(n2039), .DIN2(n2040), .Q(n2038) );
  nnd2s1 U2130 ( .DIN1(n2041), .DIN2(n2042), .Q(n2035) );
  nnd2s1 U2131 ( .DIN1(n2043), .DIN2(n2044), .Q(n2042) );
  nnd2s1 U2132 ( .DIN1(n2045), .DIN2(n2046), .Q(n2034) );
  nnd2s1 U2133 ( .DIN1(n2047), .DIN2(n2048), .Q(n2046) );
  nnd2s1 U2134 ( .DIN1(n2049), .DIN2(n2050), .Q(n2033) );
  xor2s1 U2135 ( .DIN1(n15588), .DIN2(w0[31]), .Q(n2006) );
  nnd2s1 U2136 ( .DIN1(n2051), .DIN2(n2052), .Q(\u0/N138 ) );
  nnd2s1 U2137 ( .DIN1(\key[94] ), .DIN2(ld), .Q(n2052) );
  nnd2s1 U2138 ( .DIN1(n1913), .DIN2(n1565), .Q(n2051) );
  xnr2s1 U2139 ( .DIN1(w1[30]), .DIN2(n1689), .Q(n1913) );
  xnr2s1 U2140 ( .DIN1(n2053), .DIN2(n2054), .Q(n1689) );
  nor4s1 U2141 ( .DIN1(n2055), .DIN2(n2056), .DIN3(n2057), .DIN4(n2058), 
        .Q(n2054) );
  nnd3s1 U2142 ( .DIN1(n2059), .DIN2(n2060), .DIN3(n2061), .Q(n2058) );
  nnd3s1 U2143 ( .DIN1(n2062), .DIN2(n2063), .DIN3(n2064), .Q(n2057) );
  nnd2s1 U2144 ( .DIN1(n2065), .DIN2(n2029), .Q(n2063) );
  nnd2s1 U2145 ( .DIN1(n2020), .DIN2(n2066), .Q(n2062) );
  nnd3s1 U2146 ( .DIN1(n2067), .DIN2(n2068), .DIN3(n2069), .Q(n2056) );
  or2s1 U2147 ( .DIN1(n2070), .DIN2(n2071), .Q(n2069) );
  or2s1 U2148 ( .DIN1(n2044), .DIN2(n2072), .Q(n2068) );
  nnd2s1 U2149 ( .DIN1(n2045), .DIN2(n2073), .Q(n2067) );
  nnd3s1 U2150 ( .DIN1(n2074), .DIN2(n2075), .DIN3(n2076), .Q(n2055) );
  nnd2s1 U2151 ( .DIN1(n2077), .DIN2(n2078), .Q(n2076) );
  nnd2s1 U2152 ( .DIN1(n2079), .DIN2(n2080), .Q(n2078) );
  nnd2s1 U2153 ( .DIN1(n2081), .DIN2(n2082), .Q(n2075) );
  nnd2s1 U2154 ( .DIN1(n2083), .DIN2(n2084), .Q(n2082) );
  nnd2s1 U2155 ( .DIN1(n2021), .DIN2(n2085), .Q(n2074) );
  nnd2s1 U2156 ( .DIN1(n2086), .DIN2(n2087), .Q(n2085) );
  hi1s1 U2157 ( .DIN(n2088), .Q(n2087) );
  xor2s1 U2158 ( .DIN1(n15587), .DIN2(w0[30]), .Q(n2053) );
  nnd2s1 U2159 ( .DIN1(n2089), .DIN2(n2090), .Q(\u0/N137 ) );
  nnd2s1 U2160 ( .DIN1(\key[93] ), .DIN2(ld), .Q(n2090) );
  nnd2s1 U2161 ( .DIN1(n1916), .DIN2(n1565), .Q(n2089) );
  xnr2s1 U2162 ( .DIN1(w1[29]), .DIN2(n1692), .Q(n1916) );
  xnr2s1 U2163 ( .DIN1(n2091), .DIN2(n2092), .Q(n1692) );
  nor4s1 U2164 ( .DIN1(n2093), .DIN2(n2094), .DIN3(n2095), .DIN4(n2096), 
        .Q(n2092) );
  nnd3s1 U2165 ( .DIN1(n2097), .DIN2(n2060), .DIN3(n2098), .Q(n2096) );
  nor2s1 U2166 ( .DIN1(n2099), .DIN2(n2100), .Q(n2060) );
  nnd4s1 U2167 ( .DIN1(n2101), .DIN2(n2102), .DIN3(n2103), .DIN4(n2104), 
        .Q(n2100) );
  or2s1 U2168 ( .DIN1(n2105), .DIN2(n2106), .Q(n2104) );
  nnd2s1 U2169 ( .DIN1(n2107), .DIN2(n2108), .Q(n2103) );
  nnd2s1 U2170 ( .DIN1(n2109), .DIN2(n2020), .Q(n2102) );
  nnd2s1 U2171 ( .DIN1(n2032), .DIN2(n2110), .Q(n2101) );
  nnd4s1 U2172 ( .DIN1(n2111), .DIN2(n2112), .DIN3(n2113), .DIN4(n2114), 
        .Q(n2099) );
  nnd2s1 U2173 ( .DIN1(n2031), .DIN2(n2115), .Q(n2114) );
  nnd2s1 U2174 ( .DIN1(n2083), .DIN2(n2116), .Q(n2115) );
  nnd2s1 U2175 ( .DIN1(n2117), .DIN2(n2118), .Q(n2113) );
  nnd2s1 U2176 ( .DIN1(n2079), .DIN2(n2119), .Q(n2118) );
  nnd2s1 U2177 ( .DIN1(n2120), .DIN2(n2121), .Q(n2112) );
  nnd2s1 U2178 ( .DIN1(n2122), .DIN2(n2123), .Q(n2121) );
  nnd2s1 U2179 ( .DIN1(n2041), .DIN2(n2124), .Q(n2111) );
  nnd3s1 U2180 ( .DIN1(n2083), .DIN2(n2125), .DIN3(n2126), .Q(n2124) );
  nnd4s1 U2181 ( .DIN1(n2127), .DIN2(n2128), .DIN3(n2129), .DIN4(n2018), 
        .Q(n2095) );
  nnd2s1 U2182 ( .DIN1(n2109), .DIN2(n2081), .Q(n2018) );
  nnd2s1 U2183 ( .DIN1(n2077), .DIN2(n2120), .Q(n2129) );
  nnd2s1 U2184 ( .DIN1(n2107), .DIN2(n2022), .Q(n2128) );
  nnd4s1 U2185 ( .DIN1(n2130), .DIN2(n2131), .DIN3(n2132), .DIN4(n2133), 
        .Q(n2094) );
  nnd2s1 U2186 ( .DIN1(n2134), .DIN2(n2135), .Q(n2133) );
  nnd2s1 U2187 ( .DIN1(n2032), .DIN2(n2136), .Q(n2132) );
  nnd2s1 U2188 ( .DIN1(n2019), .DIN2(n2137), .Q(n2131) );
  nnd2s1 U2189 ( .DIN1(n2065), .DIN2(n2110), .Q(n2130) );
  nnd4s1 U2190 ( .DIN1(n2138), .DIN2(n2139), .DIN3(n2140), .DIN4(n2141), 
        .Q(n2093) );
  nnd2s1 U2191 ( .DIN1(n2049), .DIN2(n2142), .Q(n2141) );
  nnd2s1 U2192 ( .DIN1(n2080), .DIN2(n2143), .Q(n2142) );
  nnd2s1 U2193 ( .DIN1(n2144), .DIN2(n2145), .Q(n2140) );
  nnd2s1 U2194 ( .DIN1(n2045), .DIN2(n2146), .Q(n2139) );
  nnd2s1 U2195 ( .DIN1(n2147), .DIN2(n2040), .Q(n2146) );
  nnd2s1 U2196 ( .DIN1(n2029), .DIN2(n2148), .Q(n2138) );
  xor2s1 U2197 ( .DIN1(n15586), .DIN2(w0[29]), .Q(n2091) );
  nnd2s1 U2198 ( .DIN1(n2149), .DIN2(n2150), .Q(\u0/N136 ) );
  nnd2s1 U2199 ( .DIN1(\key[92] ), .DIN2(ld), .Q(n2150) );
  nnd2s1 U2200 ( .DIN1(n1919), .DIN2(n1566), .Q(n2149) );
  xnr2s1 U2201 ( .DIN1(w1[28]), .DIN2(n1695), .Q(n1919) );
  xnr2s1 U2202 ( .DIN1(n2151), .DIN2(n2152), .Q(n1695) );
  nor4s1 U2203 ( .DIN1(n2153), .DIN2(n2154), .DIN3(n2155), .DIN4(n2156), 
        .Q(n2152) );
  nnd3s1 U2204 ( .DIN1(n2097), .DIN2(n2061), .DIN3(n2157), .Q(n2156) );
  and4s1 U2205 ( .DIN1(n2158), .DIN2(n2159), .DIN3(n2160), .DIN4(n2161), 
        .Q(n2061) );
  and4s1 U2206 ( .DIN1(n2162), .DIN2(n2163), .DIN3(n2164), .DIN4(n2165), 
        .Q(n2161) );
  nnd2s1 U2207 ( .DIN1(n2027), .DIN2(n2065), .Q(n2165) );
  nnd2s1 U2208 ( .DIN1(n2107), .DIN2(n2166), .Q(n2163) );
  nnd2s1 U2209 ( .DIN1(n2117), .DIN2(n2028), .Q(n2162) );
  and3s1 U2210 ( .DIN1(n2167), .DIN2(n2168), .DIN3(n2169), .Q(n2160) );
  nnd2s1 U2211 ( .DIN1(n2134), .DIN2(n2170), .Q(n2169) );
  nnd2s1 U2212 ( .DIN1(n2171), .DIN2(n2043), .Q(n2170) );
  nnd2s1 U2213 ( .DIN1(n2041), .DIN2(n2172), .Q(n2168) );
  nnd2s1 U2214 ( .DIN1(n2173), .DIN2(n2143), .Q(n2172) );
  nnd2s1 U2215 ( .DIN1(n2109), .DIN2(n2174), .Q(n2167) );
  nnd2s1 U2216 ( .DIN1(n2175), .DIN2(n2040), .Q(n2174) );
  nnd2s1 U2217 ( .DIN1(n2020), .DIN2(n2176), .Q(n2159) );
  nnd3s1 U2218 ( .DIN1(n2177), .DIN2(n2080), .DIN3(n2083), .Q(n2176) );
  nnd2s1 U2219 ( .DIN1(n2049), .DIN2(n2178), .Q(n2158) );
  nor3s1 U2220 ( .DIN1(n2179), .DIN2(n2180), .DIN3(n2181), .Q(n2097) );
  nnd4s1 U2221 ( .DIN1(n2059), .DIN2(n2182), .DIN3(n2183), .DIN4(n2184), 
        .Q(n2181) );
  and3s1 U2222 ( .DIN1(n2185), .DIN2(n2186), .DIN3(n2187), .Q(n2184) );
  nnd2s1 U2223 ( .DIN1(n2109), .DIN2(n2110), .Q(n2187) );
  nnd2s1 U2224 ( .DIN1(n2188), .DIN2(n2021), .Q(n2186) );
  nnd2s1 U2225 ( .DIN1(n2189), .DIN2(n2032), .Q(n2185) );
  nor2s1 U2226 ( .DIN1(n2190), .DIN2(n2191), .Q(n2059) );
  nnd4s1 U2227 ( .DIN1(n2192), .DIN2(n2193), .DIN3(n2194), .DIN4(n2195), 
        .Q(n2191) );
  nnd2s1 U2228 ( .DIN1(n2077), .DIN2(n2196), .Q(n2195) );
  nnd2s1 U2229 ( .DIN1(n2045), .DIN2(n2197), .Q(n2194) );
  nnd2s1 U2230 ( .DIN1(n2027), .DIN2(n2198), .Q(n2193) );
  nnd2s1 U2231 ( .DIN1(n2041), .DIN2(n2066), .Q(n2192) );
  nnd4s1 U2232 ( .DIN1(n2199), .DIN2(n2200), .DIN3(n2201), .DIN4(n2202), 
        .Q(n2190) );
  nnd2s1 U2233 ( .DIN1(n2065), .DIN2(n2197), .Q(n2202) );
  nnd2s1 U2234 ( .DIN1(n2031), .DIN2(n2203), .Q(n2201) );
  nnd2s1 U2235 ( .DIN1(n2084), .DIN2(n2119), .Q(n2203) );
  nnd2s1 U2236 ( .DIN1(n2019), .DIN2(n2204), .Q(n2200) );
  nnd2s1 U2237 ( .DIN1(n2205), .DIN2(n2206), .Q(n2204) );
  nnd2s1 U2238 ( .DIN1(n2188), .DIN2(n2207), .Q(n2199) );
  nnd3s1 U2239 ( .DIN1(n2048), .DIN2(n2208), .DIN3(n2209), .Q(n2207) );
  nnd3s1 U2240 ( .DIN1(n2210), .DIN2(n2211), .DIN3(n2023), .Q(n2180) );
  nnd2s1 U2241 ( .DIN1(n2117), .DIN2(n2108), .Q(n2023) );
  nnd2s1 U2242 ( .DIN1(n2019), .DIN2(n2212), .Q(n2211) );
  nnd3s1 U2243 ( .DIN1(n2123), .DIN2(n2213), .DIN3(n2072), .Q(n2212) );
  nor2s1 U2244 ( .DIN1(n2144), .DIN2(n2021), .Q(n2072) );
  nnd2s1 U2245 ( .DIN1(n2120), .DIN2(n2049), .Q(n2210) );
  nnd3s1 U2246 ( .DIN1(n2214), .DIN2(n2215), .DIN3(n2216), .Q(n2179) );
  nnd2s1 U2247 ( .DIN1(n2134), .DIN2(n2217), .Q(n2216) );
  nnd2s1 U2248 ( .DIN1(n2105), .DIN2(n2143), .Q(n2217) );
  nnd2s1 U2249 ( .DIN1(n2029), .DIN2(n2218), .Q(n2215) );
  nnd2s1 U2250 ( .DIN1(n2119), .DIN2(n2105), .Q(n2218) );
  nnd2s1 U2251 ( .DIN1(n2077), .DIN2(n2219), .Q(n2214) );
  nnd2s1 U2252 ( .DIN1(n2173), .DIN2(n2084), .Q(n2219) );
  nnd3s1 U2253 ( .DIN1(n2220), .DIN2(n2221), .DIN3(n2222), .Q(n2155) );
  nnd3s1 U2254 ( .DIN1(n2223), .DIN2(n2224), .DIN3(n2225), .Q(n2154) );
  nnd2s1 U2255 ( .DIN1(n2107), .DIN2(n2198), .Q(n2225) );
  nnd2s1 U2256 ( .DIN1(n2029), .DIN2(n2135), .Q(n2224) );
  nnd2s1 U2257 ( .DIN1(n2120), .DIN2(n2136), .Q(n2223) );
  nnd4s1 U2258 ( .DIN1(n2226), .DIN2(n2227), .DIN3(n2228), .DIN4(n2229), 
        .Q(n2153) );
  nnd2s1 U2259 ( .DIN1(n2027), .DIN2(n2230), .Q(n2229) );
  nnd2s1 U2260 ( .DIN1(n2116), .DIN2(n2080), .Q(n2230) );
  nnd2s1 U2261 ( .DIN1(n2065), .DIN2(n2231), .Q(n2228) );
  nnd2s1 U2262 ( .DIN1(n2209), .DIN2(n2205), .Q(n2231) );
  nnd2s1 U2263 ( .DIN1(n2081), .DIN2(n2232), .Q(n2227) );
  nnd2s1 U2264 ( .DIN1(n2037), .DIN2(n2233), .Q(n2226) );
  nnd2s1 U2265 ( .DIN1(n2234), .DIN2(n2206), .Q(n2233) );
  xor2s1 U2266 ( .DIN1(n15585), .DIN2(w0[28]), .Q(n2151) );
  nnd2s1 U2267 ( .DIN1(n2235), .DIN2(n2236), .Q(\u0/N135 ) );
  nnd2s1 U2268 ( .DIN1(\key[91] ), .DIN2(ld), .Q(n2236) );
  nnd2s1 U2269 ( .DIN1(n1922), .DIN2(n1566), .Q(n2235) );
  xnr2s1 U2270 ( .DIN1(w1[27]), .DIN2(n1698), .Q(n1922) );
  xnr2s1 U2271 ( .DIN1(n2237), .DIN2(n2238), .Q(n1698) );
  nor4s1 U2272 ( .DIN1(n2239), .DIN2(n2240), .DIN3(n2241), .DIN4(n2242), 
        .Q(n2238) );
  nnd3s1 U2273 ( .DIN1(n2098), .DIN2(n2183), .DIN3(n2157), .Q(n2242) );
  nor4s1 U2274 ( .DIN1(n2243), .DIN2(n2244), .DIN3(n2245), .DIN4(n2246), 
        .Q(n2157) );
  nnd4s1 U2275 ( .DIN1(n2247), .DIN2(n2248), .DIN3(n2249), .DIN4(n2250), 
        .Q(n2246) );
  nnd2s1 U2276 ( .DIN1(n2032), .DIN2(n2081), .Q(n2250) );
  nor2s1 U2277 ( .DIN1(n2251), .DIN2(n2252), .Q(n2249) );
  nor2s1 U2278 ( .DIN1(n2080), .DIN2(n2253), .Q(n2252) );
  nor2s1 U2279 ( .DIN1(n2143), .DIN2(n2254), .Q(n2251) );
  nnd2s1 U2280 ( .DIN1(n2022), .DIN2(n2110), .Q(n2248) );
  nnd2s1 U2281 ( .DIN1(n2117), .DIN2(n2045), .Q(n2247) );
  nnd3s1 U2282 ( .DIN1(n2255), .DIN2(n2256), .DIN3(n2257), .Q(n2245) );
  nnd2s1 U2283 ( .DIN1(n2144), .DIN2(n2148), .Q(n2257) );
  nnd2s1 U2284 ( .DIN1(n2030), .DIN2(n2258), .Q(n2256) );
  nnd3s1 U2285 ( .DIN1(n2208), .DIN2(n2175), .DIN3(n2253), .Q(n2258) );
  nnd2s1 U2286 ( .DIN1(n2189), .DIN2(n2259), .Q(n2255) );
  nnd3s1 U2287 ( .DIN1(n2105), .DIN2(n2044), .DIN3(n2079), .Q(n2259) );
  nor2s1 U2288 ( .DIN1(n2105), .DIN2(n2048), .Q(n2244) );
  nor2s1 U2289 ( .DIN1(n2260), .DIN2(n2261), .Q(n2243) );
  nor4s1 U2290 ( .DIN1(n2262), .DIN2(n2263), .DIN3(n2264), .DIN4(n2265), 
        .Q(n2183) );
  nnd4s1 U2291 ( .DIN1(n2266), .DIN2(n2267), .DIN3(n2268), .DIN4(n2269), 
        .Q(n2265) );
  nor2s1 U2292 ( .DIN1(n2270), .DIN2(n2271), .Q(n2269) );
  nor2s1 U2293 ( .DIN1(n2253), .DIN2(n2261), .Q(n2271) );
  nor2s1 U2294 ( .DIN1(n2147), .DIN2(n2044), .Q(n2270) );
  nnd2s1 U2295 ( .DIN1(n2066), .DIN2(n2049), .Q(n2267) );
  nnd2s1 U2296 ( .DIN1(n2120), .DIN2(n2029), .Q(n2266) );
  nnd3s1 U2297 ( .DIN1(n2272), .DIN2(n2273), .DIN3(n2274), .Q(n2264) );
  nnd2s1 U2298 ( .DIN1(n2108), .DIN2(n2275), .Q(n2274) );
  nnd2s1 U2299 ( .DIN1(n2209), .DIN2(n2123), .Q(n2275) );
  nnd2s1 U2300 ( .DIN1(n2065), .DIN2(n2276), .Q(n2273) );
  nnd2s1 U2301 ( .DIN1(n2234), .DIN2(n2175), .Q(n2276) );
  nnd2s1 U2302 ( .DIN1(n2031), .DIN2(n2145), .Q(n2272) );
  nnd2s1 U2303 ( .DIN1(n2125), .DIN2(n2277), .Q(n2145) );
  nor2s1 U2304 ( .DIN1(n2278), .DIN2(n2084), .Q(n2263) );
  nor2s1 U2305 ( .DIN1(n2020), .DIN2(n2041), .Q(n2278) );
  nor2s1 U2306 ( .DIN1(n2279), .DIN2(n2206), .Q(n2262) );
  and2s1 U2307 ( .DIN1(n2105), .DIN2(n2280), .Q(n2279) );
  nor4s1 U2308 ( .DIN1(n2281), .DIN2(n2282), .DIN3(n2283), .DIN4(n2284), 
        .Q(n2098) );
  nnd4s1 U2309 ( .DIN1(n2285), .DIN2(n2286), .DIN3(n2287), .DIN4(n2288), 
        .Q(n2284) );
  nnd2s1 U2310 ( .DIN1(n2188), .DIN2(n2110), .Q(n2288) );
  nor2s1 U2311 ( .DIN1(n2289), .DIN2(n2290), .Q(n2287) );
  nor2s1 U2312 ( .DIN1(n2084), .DIN2(n2291), .Q(n2289) );
  nnd2s1 U2313 ( .DIN1(n2109), .DIN2(n2117), .Q(n2286) );
  nnd2s1 U2314 ( .DIN1(n2107), .DIN2(n2037), .Q(n2285) );
  nnd3s1 U2315 ( .DIN1(n2292), .DIN2(n2293), .DIN3(n2294), .Q(n2283) );
  nnd2s1 U2316 ( .DIN1(n2029), .DIN2(n2295), .Q(n2294) );
  nnd2s1 U2317 ( .DIN1(n2045), .DIN2(n2296), .Q(n2293) );
  nnd2s1 U2318 ( .DIN1(n2206), .DIN2(n2175), .Q(n2296) );
  nnd2s1 U2319 ( .DIN1(n2189), .DIN2(n2297), .Q(n2292) );
  nnd3s1 U2320 ( .DIN1(n2177), .DIN2(n2261), .DIN3(n2298), .Q(n2297) );
  nor2s1 U2321 ( .DIN1(n2044), .DIN2(n2048), .Q(n2282) );
  nor2s1 U2322 ( .DIN1(n2086), .DIN2(n2040), .Q(n2281) );
  nnd3s1 U2323 ( .DIN1(n2299), .DIN2(n2300), .DIN3(n2064), .Q(n2241) );
  nor3s1 U2324 ( .DIN1(n2301), .DIN2(n2302), .DIN3(n2303), .Q(n2064) );
  nnd4s1 U2325 ( .DIN1(n2182), .DIN2(n2127), .DIN3(n2222), .DIN4(n2304), 
        .Q(n2303) );
  and3s1 U2326 ( .DIN1(n2305), .DIN2(n2306), .DIN3(n2307), .Q(n2304) );
  nnd2s1 U2327 ( .DIN1(n2107), .DIN2(n2028), .Q(n2307) );
  nnd2s1 U2328 ( .DIN1(n2019), .DIN2(n2081), .Q(n2305) );
  nor4s1 U2329 ( .DIN1(n2308), .DIN2(n2309), .DIN3(n2310), .DIN4(n2311), 
        .Q(n2222) );
  nnd4s1 U2330 ( .DIN1(n2312), .DIN2(n2313), .DIN3(n2314), .DIN4(n2315), 
        .Q(n2311) );
  nnd2s1 U2331 ( .DIN1(n2107), .DIN2(n2316), .Q(n2315) );
  nnd2s1 U2332 ( .DIN1(n2317), .DIN2(n2177), .Q(n2316) );
  nor2s1 U2333 ( .DIN1(n2318), .DIN2(n2319), .Q(n2314) );
  nor2s1 U2334 ( .DIN1(n2320), .DIN2(n2147), .Q(n2319) );
  nor2s1 U2335 ( .DIN1(n2019), .DIN2(n2088), .Q(n2320) );
  nor2s1 U2336 ( .DIN1(n2321), .DIN2(n2047), .Q(n2318) );
  nor2s1 U2337 ( .DIN1(n2178), .DIN2(n2120), .Q(n2321) );
  nnd2s1 U2338 ( .DIN1(n2037), .DIN2(n2322), .Q(n2313) );
  nnd3s1 U2339 ( .DIN1(n2048), .DIN2(n2205), .DIN3(n2291), .Q(n2322) );
  nnd2s1 U2340 ( .DIN1(n2189), .DIN2(n2178), .Q(n2312) );
  nnd3s1 U2341 ( .DIN1(n2323), .DIN2(n2324), .DIN3(n2325), .Q(n2310) );
  nnd2s1 U2342 ( .DIN1(n2326), .DIN2(n2144), .Q(n2325) );
  nnd2s1 U2343 ( .DIN1(n2027), .DIN2(n2030), .Q(n2324) );
  nnd2s1 U2344 ( .DIN1(n2031), .DIN2(n2065), .Q(n2323) );
  nor2s1 U2345 ( .DIN1(n2253), .DIN2(n2084), .Q(n2309) );
  nor2s1 U2346 ( .DIN1(n2261), .DIN2(n2234), .Q(n2308) );
  nor4s1 U2347 ( .DIN1(n2327), .DIN2(n2328), .DIN3(n2329), .DIN4(n2330), 
        .Q(n2127) );
  nnd4s1 U2348 ( .DIN1(n2331), .DIN2(n2332), .DIN3(n2333), .DIN4(n2334), 
        .Q(n2330) );
  nnd2s1 U2349 ( .DIN1(n2028), .DIN2(n2049), .Q(n2334) );
  nnd2s1 U2350 ( .DIN1(n2081), .DIN2(n2108), .Q(n2333) );
  nnd2s1 U2351 ( .DIN1(n2134), .DIN2(n2037), .Q(n2332) );
  nnd2s1 U2352 ( .DIN1(n2107), .DIN2(n2109), .Q(n2331) );
  nnd3s1 U2353 ( .DIN1(n2335), .DIN2(n2336), .DIN3(n2337), .Q(n2329) );
  nnd2s1 U2354 ( .DIN1(n2021), .DIN2(n2338), .Q(n2337) );
  nnd3s1 U2355 ( .DIN1(n2119), .DIN2(n2084), .DIN3(n2277), .Q(n2338) );
  nnd2s1 U2356 ( .DIN1(n2137), .DIN2(n2339), .Q(n2336) );
  nnd2s1 U2357 ( .DIN1(n2280), .DIN2(n2119), .Q(n2339) );
  nor2s1 U2358 ( .DIN1(n2326), .DIN2(n2178), .Q(n2280) );
  nnd2s1 U2359 ( .DIN1(n2188), .DIN2(n2340), .Q(n2335) );
  nnd2s1 U2360 ( .DIN1(n2254), .DIN2(n2234), .Q(n2340) );
  nor2s1 U2361 ( .DIN1(n2177), .DIN2(n2209), .Q(n2328) );
  nor2s1 U2362 ( .DIN1(n2126), .DIN2(n2206), .Q(n2327) );
  hi1s1 U2363 ( .DIN(n2050), .Q(n2126) );
  nor2s1 U2364 ( .DIN1(n2341), .DIN2(n2342), .Q(n2182) );
  nnd4s1 U2365 ( .DIN1(n2343), .DIN2(n2344), .DIN3(n2345), .DIN4(n2346), 
        .Q(n2342) );
  nnd2s1 U2366 ( .DIN1(n2028), .DIN2(n2347), .Q(n2346) );
  nnd3s1 U2367 ( .DIN1(n2206), .DIN2(n2253), .DIN3(n2291), .Q(n2347) );
  nnd2s1 U2368 ( .DIN1(n2027), .DIN2(n2120), .Q(n2344) );
  nnd4s1 U2369 ( .DIN1(n2348), .DIN2(n2349), .DIN3(n2350), .DIN4(n2351), 
        .Q(n2341) );
  nnd2s1 U2370 ( .DIN1(n2049), .DIN2(n2352), .Q(n2351) );
  nnd2s1 U2371 ( .DIN1(n2353), .DIN2(n2084), .Q(n2352) );
  nnd2s1 U2372 ( .DIN1(n2020), .DIN2(n2354), .Q(n2350) );
  nnd2s1 U2373 ( .DIN1(n2045), .DIN2(n2355), .Q(n2349) );
  nnd2s1 U2374 ( .DIN1(n2209), .DIN2(n2291), .Q(n2355) );
  nnd2s1 U2375 ( .DIN1(n2188), .DIN2(n2356), .Q(n2348) );
  nnd2s1 U2376 ( .DIN1(n2071), .DIN2(n2205), .Q(n2356) );
  nnd3s1 U2377 ( .DIN1(n2357), .DIN2(n2358), .DIN3(n2359), .Q(n2302) );
  nnd2s1 U2378 ( .DIN1(n2029), .DIN2(n2037), .Q(n2359) );
  nnd2s1 U2379 ( .DIN1(n2178), .DIN2(n2360), .Q(n2358) );
  nnd3s1 U2380 ( .DIN1(n2253), .DIN2(n2048), .DIN3(n2361), .Q(n2360) );
  or2s1 U2381 ( .DIN1(n2119), .DIN2(n2362), .Q(n2357) );
  nnd3s1 U2382 ( .DIN1(n2363), .DIN2(n2364), .DIN3(n2365), .Q(n2301) );
  nnd2s1 U2383 ( .DIN1(n2045), .DIN2(n2366), .Q(n2365) );
  nnd2s1 U2384 ( .DIN1(n2213), .DIN2(n2208), .Q(n2366) );
  nnd2s1 U2385 ( .DIN1(n2117), .DIN2(n2367), .Q(n2364) );
  or2s1 U2386 ( .DIN1(n2148), .DIN2(n2030), .Q(n2367) );
  nnd2s1 U2387 ( .DIN1(n2084), .DIN2(n2070), .Q(n2148) );
  nnd2s1 U2388 ( .DIN1(n2144), .DIN2(n2368), .Q(n2363) );
  nnd2s1 U2389 ( .DIN1(n2043), .DIN2(n2105), .Q(n2368) );
  nnd2s1 U2390 ( .DIN1(n2081), .DIN2(n2066), .Q(n2300) );
  nnd2s1 U2391 ( .DIN1(n2041), .DIN2(n2109), .Q(n2299) );
  nnd3s1 U2392 ( .DIN1(n2369), .DIN2(n2370), .DIN3(n2371), .Q(n2240) );
  nnd2s1 U2393 ( .DIN1(n2326), .DIN2(n2049), .Q(n2371) );
  nnd2s1 U2394 ( .DIN1(n2166), .DIN2(n2372), .Q(n2370) );
  nnd4s1 U2395 ( .DIN1(n2373), .DIN2(n2374), .DIN3(n2375), .DIN4(n2376), 
        .Q(n2239) );
  nnd2s1 U2396 ( .DIN1(n2137), .DIN2(n2377), .Q(n2376) );
  nnd2s1 U2397 ( .DIN1(n2086), .DIN2(n2143), .Q(n2377) );
  nor2s1 U2398 ( .DIN1(n2120), .DIN2(n2108), .Q(n2086) );
  nnd2s1 U2399 ( .DIN1(n2108), .DIN2(n2378), .Q(n2375) );
  nnd2s1 U2400 ( .DIN1(n2122), .DIN2(n2208), .Q(n2378) );
  nnd2s1 U2401 ( .DIN1(n2022), .DIN2(n2379), .Q(n2374) );
  nnd2s1 U2402 ( .DIN1(n2123), .DIN2(n2048), .Q(n2379) );
  nnd2s1 U2403 ( .DIN1(n2037), .DIN2(n2197), .Q(n2373) );
  xor2s1 U2404 ( .DIN1(n15584), .DIN2(w0[27]), .Q(n2237) );
  nnd2s1 U2405 ( .DIN1(n2380), .DIN2(n2381), .Q(\u0/N134 ) );
  nnd2s1 U2406 ( .DIN1(\key[90] ), .DIN2(ld), .Q(n2381) );
  nnd2s1 U2407 ( .DIN1(n1925), .DIN2(n1566), .Q(n2380) );
  xnr2s1 U2408 ( .DIN1(w1[26]), .DIN2(n1701), .Q(n1925) );
  xnr2s1 U2409 ( .DIN1(n2382), .DIN2(n2383), .Q(n1701) );
  nor4s1 U2410 ( .DIN1(n2384), .DIN2(n2385), .DIN3(n2386), .DIN4(n2387), 
        .Q(n2383) );
  nnd3s1 U2411 ( .DIN1(n2388), .DIN2(n2389), .DIN3(n2390), .Q(n2387) );
  nnd3s1 U2412 ( .DIN1(n2391), .DIN2(n2392), .DIN3(n2015), .Q(n2386) );
  nor3s1 U2413 ( .DIN1(n2393), .DIN2(n2394), .DIN3(n2395), .Q(n2015) );
  nnd4s1 U2414 ( .DIN1(n2396), .DIN2(n2397), .DIN3(n2398), .DIN4(n2399), 
        .Q(n2395) );
  and3s1 U2415 ( .DIN1(n2400), .DIN2(n2401), .DIN3(n2402), .Q(n2399) );
  nnd2s1 U2416 ( .DIN1(n2077), .DIN2(n2022), .Q(n2402) );
  nnd2s1 U2417 ( .DIN1(n2027), .DIN2(n2109), .Q(n2401) );
  nnd2s1 U2418 ( .DIN1(n2041), .DIN2(n2108), .Q(n2400) );
  nnd3s1 U2419 ( .DIN1(n2403), .DIN2(n2404), .DIN3(n2345), .Q(n2394) );
  nnd2s1 U2420 ( .DIN1(n2107), .DIN2(n2178), .Q(n2345) );
  or2s1 U2421 ( .DIN1(n2047), .DIN2(n2353), .Q(n2404) );
  nor2s1 U2422 ( .DIN1(n2019), .DIN2(n2030), .Q(n2353) );
  nnd2s1 U2423 ( .DIN1(n2137), .DIN2(n2088), .Q(n2403) );
  nnd2s1 U2424 ( .DIN1(n2125), .DIN2(n2079), .Q(n2088) );
  nnd4s1 U2425 ( .DIN1(n2405), .DIN2(n2406), .DIN3(n2407), .DIN4(n2408), 
        .Q(n2393) );
  nnd2s1 U2426 ( .DIN1(n2166), .DIN2(n2409), .Q(n2408) );
  nnd2s1 U2427 ( .DIN1(n2021), .DIN2(n2410), .Q(n2407) );
  nnd2s1 U2428 ( .DIN1(n2079), .DIN2(n2143), .Q(n2410) );
  nnd2s1 U2429 ( .DIN1(n2120), .DIN2(n2411), .Q(n2406) );
  nnd2s1 U2430 ( .DIN1(n2123), .DIN2(n2040), .Q(n2411) );
  nnd2s1 U2431 ( .DIN1(n2045), .DIN2(n2412), .Q(n2405) );
  nnd2s1 U2432 ( .DIN1(n2361), .DIN2(n2253), .Q(n2412) );
  hi1s1 U2433 ( .DIN(n2136), .Q(n2361) );
  nnd2s1 U2434 ( .DIN1(n2205), .DIN2(n2147), .Q(n2136) );
  nnd2s1 U2435 ( .DIN1(n2041), .DIN2(n2032), .Q(n2392) );
  nnd2s1 U2436 ( .DIN1(n2037), .DIN2(n2110), .Q(n2391) );
  nnd3s1 U2437 ( .DIN1(n2413), .DIN2(n2414), .DIN3(n2415), .Q(n2385) );
  nnd2s1 U2438 ( .DIN1(n2109), .DIN2(n2029), .Q(n2415) );
  or2s1 U2439 ( .DIN1(n2043), .DIN2(n2039), .Q(n2414) );
  nor2s1 U2440 ( .DIN1(n2077), .DIN2(n2081), .Q(n2039) );
  nnd2s1 U2441 ( .DIN1(n2188), .DIN2(n2049), .Q(n2413) );
  nnd4s1 U2442 ( .DIN1(n2416), .DIN2(n2417), .DIN3(n2418), .DIN4(n2419), 
        .Q(n2384) );
  nnd2s1 U2443 ( .DIN1(n2326), .DIN2(n2420), .Q(n2419) );
  nnd2s1 U2444 ( .DIN1(n2362), .DIN2(n2205), .Q(n2420) );
  nnd2s1 U2445 ( .DIN1(n2020), .DIN2(n2421), .Q(n2418) );
  nnd2s1 U2446 ( .DIN1(n2173), .DIN2(n2080), .Q(n2421) );
  nor2s1 U2447 ( .DIN1(n2028), .DIN2(n2178), .Q(n2173) );
  nnd2s1 U2448 ( .DIN1(n2021), .DIN2(n2422), .Q(n2417) );
  nnd2s1 U2449 ( .DIN1(n2022), .DIN2(n2409), .Q(n2416) );
  nnd2s1 U2450 ( .DIN1(n2209), .DIN2(n2040), .Q(n2409) );
  xor2s1 U2451 ( .DIN1(n15583), .DIN2(w0[26]), .Q(n2382) );
  nnd2s1 U2452 ( .DIN1(n2423), .DIN2(n2424), .Q(\u0/N133 ) );
  nnd2s1 U2453 ( .DIN1(\key[89] ), .DIN2(ld), .Q(n2424) );
  nnd2s1 U2454 ( .DIN1(n1928), .DIN2(n1566), .Q(n2423) );
  xnr2s1 U2455 ( .DIN1(w1[25]), .DIN2(n1704), .Q(n1928) );
  xnr2s1 U2456 ( .DIN1(n2425), .DIN2(n2426), .Q(n1704) );
  nor4s1 U2457 ( .DIN1(n2427), .DIN2(n2428), .DIN3(n2429), .DIN4(n2430), 
        .Q(n2426) );
  nnd3s1 U2458 ( .DIN1(n2390), .DIN2(n2012), .DIN3(n2431), .Q(n2430) );
  nor2s1 U2459 ( .DIN1(n2432), .DIN2(n2433), .Q(n2012) );
  nnd4s1 U2460 ( .DIN1(n2434), .DIN2(n2435), .DIN3(n2436), .DIN4(n2437), 
        .Q(n2433) );
  nnd2s1 U2461 ( .DIN1(n2032), .DIN2(n2197), .Q(n2437) );
  nnd2s1 U2462 ( .DIN1(n2123), .DIN2(n2047), .Q(n2197) );
  nnd2s1 U2463 ( .DIN1(n2028), .DIN2(n2029), .Q(n2436) );
  nnd2s1 U2464 ( .DIN1(n2021), .DIN2(n2120), .Q(n2435) );
  nnd2s1 U2465 ( .DIN1(n2188), .DIN2(n2144), .Q(n2434) );
  nnd4s1 U2466 ( .DIN1(n2438), .DIN2(n2439), .DIN3(n2440), .DIN4(n2441), 
        .Q(n2432) );
  nnd2s1 U2467 ( .DIN1(n2065), .DIN2(n2442), .Q(n2441) );
  or2s1 U2468 ( .DIN1(n2372), .DIN2(n2031), .Q(n2442) );
  nnd2s1 U2469 ( .DIN1(n2110), .DIN2(n2443), .Q(n2440) );
  nnd2s1 U2470 ( .DIN1(n2070), .DIN2(n2119), .Q(n2443) );
  nnd2s1 U2471 ( .DIN1(n2022), .DIN2(n2444), .Q(n2439) );
  nnd2s1 U2472 ( .DIN1(n2213), .DIN2(n2048), .Q(n2444) );
  nnd2s1 U2473 ( .DIN1(n2045), .DIN2(n2445), .Q(n2438) );
  nnd3s1 U2474 ( .DIN1(n2209), .DIN2(n2213), .DIN3(n2446), .Q(n2445) );
  nor4s1 U2475 ( .DIN1(n2447), .DIN2(n2448), .DIN3(n2449), .DIN4(n2450), 
        .Q(n2390) );
  nnd4s1 U2476 ( .DIN1(n2451), .DIN2(n2343), .DIN3(n2452), .DIN4(n2453), 
        .Q(n2450) );
  nnd2s1 U2477 ( .DIN1(n2134), .DIN2(n2050), .Q(n2453) );
  nnd2s1 U2478 ( .DIN1(n2137), .DIN2(n2022), .Q(n2452) );
  nnd2s1 U2479 ( .DIN1(n2031), .DIN2(n2326), .Q(n2343) );
  nnd2s1 U2480 ( .DIN1(n2077), .DIN2(n2166), .Q(n2451) );
  nnd3s1 U2481 ( .DIN1(n2454), .DIN2(n2455), .DIN3(n2456), .Q(n2449) );
  nnd2s1 U2482 ( .DIN1(n2037), .DIN2(n2457), .Q(n2456) );
  nnd2s1 U2483 ( .DIN1(n2027), .DIN2(n2458), .Q(n2455) );
  nnd2s1 U2484 ( .DIN1(n2083), .DIN2(n2080), .Q(n2458) );
  nnd2s1 U2485 ( .DIN1(n2066), .DIN2(n2459), .Q(n2454) );
  nnd2s1 U2486 ( .DIN1(n2071), .DIN2(n2047), .Q(n2459) );
  nor2s1 U2487 ( .DIN1(n2260), .DIN2(n2116), .Q(n2448) );
  nor2s1 U2488 ( .DIN1(n2144), .DIN2(n2137), .Q(n2260) );
  nor2s1 U2489 ( .DIN1(n2460), .DIN2(n2254), .Q(n2447) );
  nor2s1 U2490 ( .DIN1(n2120), .DIN2(n2109), .Q(n2460) );
  nnd3s1 U2491 ( .DIN1(n2461), .DIN2(n2220), .DIN3(n2397), .Q(n2429) );
  nor2s1 U2492 ( .DIN1(n2462), .DIN2(n2463), .Q(n2397) );
  nnd4s1 U2493 ( .DIN1(n2464), .DIN2(n2465), .DIN3(n2369), .DIN4(n2466), 
        .Q(n2463) );
  nnd2s1 U2494 ( .DIN1(n2066), .DIN2(n2073), .Q(n2466) );
  nnd2s1 U2495 ( .DIN1(n2234), .DIN2(n2048), .Q(n2073) );
  nnd2s1 U2496 ( .DIN1(n2077), .DIN2(n2030), .Q(n2369) );
  nnd2s1 U2497 ( .DIN1(n2189), .DIN2(n2166), .Q(n2465) );
  nnd2s1 U2498 ( .DIN1(n2022), .DIN2(n2081), .Q(n2464) );
  nnd4s1 U2499 ( .DIN1(n2467), .DIN2(n2468), .DIN3(n2469), .DIN4(n2470), 
        .Q(n2462) );
  nnd2s1 U2500 ( .DIN1(n2031), .DIN2(n2471), .Q(n2470) );
  nnd2s1 U2501 ( .DIN1(n2261), .DIN2(n2277), .Q(n2471) );
  nnd2s1 U2502 ( .DIN1(n2134), .DIN2(n2472), .Q(n2469) );
  nnd2s1 U2503 ( .DIN1(n2125), .DIN2(n2143), .Q(n2472) );
  nnd2s1 U2504 ( .DIN1(n2107), .DIN2(n2473), .Q(n2468) );
  nnd3s1 U2505 ( .DIN1(n2070), .DIN2(n2084), .DIN3(n2080), .Q(n2473) );
  nnd2s1 U2506 ( .DIN1(n2117), .DIN2(n2474), .Q(n2467) );
  nnd4s1 U2507 ( .DIN1(n2083), .DIN2(n2105), .DIN3(n2177), .DIN4(n2125), 
        .Q(n2474) );
  nnd2s1 U2508 ( .DIN1(n2032), .DIN2(n2134), .Q(n2220) );
  nnd2s1 U2509 ( .DIN1(n2189), .DIN2(n2045), .Q(n2461) );
  nnd3s1 U2510 ( .DIN1(n2475), .DIN2(n2476), .DIN3(n2477), .Q(n2428) );
  nnd2s1 U2511 ( .DIN1(n2077), .DIN2(n2108), .Q(n2477) );
  nnd2s1 U2512 ( .DIN1(n2031), .DIN2(n2028), .Q(n2476) );
  nnd2s1 U2513 ( .DIN1(n2166), .DIN2(n2020), .Q(n2475) );
  nnd4s1 U2514 ( .DIN1(n2478), .DIN2(n2479), .DIN3(n2480), .DIN4(n2481), 
        .Q(n2427) );
  nnd2s1 U2515 ( .DIN1(n2178), .DIN2(n2482), .Q(n2481) );
  nnd2s1 U2516 ( .DIN1(n2205), .DIN2(n2175), .Q(n2482) );
  nnd2s1 U2517 ( .DIN1(n2037), .DIN2(n2483), .Q(n2480) );
  nnd2s1 U2518 ( .DIN1(n2254), .DIN2(n2209), .Q(n2483) );
  nnd2s1 U2519 ( .DIN1(n2109), .DIN2(n2484), .Q(n2479) );
  nnd2s1 U2520 ( .DIN1(n2106), .DIN2(n2234), .Q(n2484) );
  nor2s1 U2521 ( .DIN1(n2021), .DIN2(n2137), .Q(n2106) );
  nnd2s1 U2522 ( .DIN1(n2120), .DIN2(n2485), .Q(n2478) );
  nnd3s1 U2523 ( .DIN1(n2206), .DIN2(n2208), .DIN3(n2071), .Q(n2485) );
  nor2s1 U2524 ( .DIN1(n2049), .DIN2(n2137), .Q(n2071) );
  xor2s1 U2525 ( .DIN1(n15582), .DIN2(w0[25]), .Q(n2425) );
  nnd2s1 U2526 ( .DIN1(n2486), .DIN2(n2487), .Q(\u0/N132 ) );
  nnd2s1 U2527 ( .DIN1(\key[88] ), .DIN2(ld), .Q(n2487) );
  nnd2s1 U2528 ( .DIN1(n1931), .DIN2(n1566), .Q(n2486) );
  xnr2s1 U2529 ( .DIN1(w1[24]), .DIN2(n1707), .Q(n1931) );
  xnr2s1 U2530 ( .DIN1(n2488), .DIN2(n2489), .Q(n1707) );
  nor4s1 U2531 ( .DIN1(n2490), .DIN2(n2491), .DIN3(n2492), .DIN4(n2493), 
        .Q(n2489) );
  nnd3s1 U2532 ( .DIN1(n2389), .DIN2(n2014), .DIN3(n2431), .Q(n2493) );
  nor3s1 U2533 ( .DIN1(n2494), .DIN2(n2495), .DIN3(n2496), .Q(n2431) );
  nnd4s1 U2534 ( .DIN1(n2013), .DIN2(n2396), .DIN3(n2388), .DIN4(n2497), 
        .Q(n2496) );
  and3s1 U2535 ( .DIN1(n2498), .DIN2(n2499), .DIN3(n2500), .Q(n2497) );
  nnd2s1 U2536 ( .DIN1(n2109), .DIN2(n2134), .Q(n2500) );
  nnd2s1 U2537 ( .DIN1(n2022), .DIN2(n2117), .Q(n2499) );
  nnd2s1 U2538 ( .DIN1(n2189), .DIN2(n2037), .Q(n2498) );
  hi1s1 U2539 ( .DIN(n2125), .Q(n2037) );
  and4s1 U2540 ( .DIN1(n2501), .DIN2(n2502), .DIN3(n2503), .DIN4(n2504), 
        .Q(n2388) );
  and4s1 U2541 ( .DIN1(n2505), .DIN2(n2506), .DIN3(n2268), .DIN4(n2164), 
        .Q(n2504) );
  nnd2s1 U2542 ( .DIN1(n2031), .DIN2(n2066), .Q(n2164) );
  nnd2s1 U2543 ( .DIN1(n2107), .DIN2(n2019), .Q(n2268) );
  nnd2s1 U2544 ( .DIN1(n2077), .DIN2(n2045), .Q(n2506) );
  nnd2s1 U2545 ( .DIN1(n2189), .DIN2(n2109), .Q(n2505) );
  and3s1 U2546 ( .DIN1(n2507), .DIN2(n2508), .DIN3(n2509), .Q(n2503) );
  nnd2s1 U2547 ( .DIN1(n2032), .DIN2(n2457), .Q(n2509) );
  nnd2s1 U2548 ( .DIN1(n2175), .DIN2(n2147), .Q(n2457) );
  nnd2s1 U2549 ( .DIN1(n2029), .DIN2(n2510), .Q(n2508) );
  nnd2s1 U2550 ( .DIN1(n2298), .DIN2(n2125), .Q(n2510) );
  nor2s1 U2551 ( .DIN1(n2188), .DIN2(n2166), .Q(n2298) );
  nnd2s1 U2552 ( .DIN1(n2326), .DIN2(n2511), .Q(n2507) );
  nnd2s1 U2553 ( .DIN1(n2209), .DIN2(n2047), .Q(n2511) );
  nnd2s1 U2554 ( .DIN1(n2188), .DIN2(n2512), .Q(n2502) );
  nnd2s1 U2555 ( .DIN1(n2234), .DIN2(n2040), .Q(n2512) );
  nnd2s1 U2556 ( .DIN1(n2110), .DIN2(n2513), .Q(n2501) );
  nnd3s1 U2557 ( .DIN1(n2044), .DIN2(n2084), .DIN3(n2080), .Q(n2513) );
  nor4s1 U2558 ( .DIN1(n2514), .DIN2(n2515), .DIN3(n2516), .DIN4(n2517), 
        .Q(n2396) );
  nnd4s1 U2559 ( .DIN1(n2518), .DIN2(n2519), .DIN3(n2520), .DIN4(n2521), 
        .Q(n2517) );
  and3s1 U2560 ( .DIN1(n2522), .DIN2(n2523), .DIN3(n2524), .Q(n2521) );
  nnd2s1 U2561 ( .DIN1(n2027), .DIN2(n2178), .Q(n2524) );
  nnd2s1 U2562 ( .DIN1(n2028), .DIN2(n2525), .Q(n2523) );
  nnd2s1 U2563 ( .DIN1(n2123), .DIN2(n2526), .Q(n2525) );
  nnd2s1 U2564 ( .DIN1(n2041), .DIN2(n2422), .Q(n2522) );
  nnd2s1 U2565 ( .DIN1(n2116), .DIN2(n2119), .Q(n2422) );
  nnd2s1 U2566 ( .DIN1(n2020), .DIN2(n2527), .Q(n2520) );
  nnd2s1 U2567 ( .DIN1(n2083), .DIN2(n2143), .Q(n2527) );
  nnd2s1 U2568 ( .DIN1(n2030), .DIN2(n2528), .Q(n2519) );
  nnd2s1 U2569 ( .DIN1(n2040), .DIN2(n2048), .Q(n2528) );
  nnd2s1 U2570 ( .DIN1(n2326), .DIN2(n2529), .Q(n2518) );
  nnd2s1 U2571 ( .DIN1(n2253), .DIN2(n2254), .Q(n2529) );
  nnd3s1 U2572 ( .DIN1(n2530), .DIN2(n2531), .DIN3(n2532), .Q(n2516) );
  nnd2s1 U2573 ( .DIN1(n2144), .DIN2(n2108), .Q(n2532) );
  nnd2s1 U2574 ( .DIN1(n2137), .DIN2(n2065), .Q(n2531) );
  nnd2s1 U2575 ( .DIN1(n2032), .DIN2(n2049), .Q(n2530) );
  nor2s1 U2576 ( .DIN1(n2206), .DIN2(n2317), .Q(n2515) );
  nor2s1 U2577 ( .DIN1(n2116), .DIN2(n2234), .Q(n2514) );
  nor4s1 U2578 ( .DIN1(n2533), .DIN2(n2534), .DIN3(n2535), .DIN4(n2536), 
        .Q(n2013) );
  nnd4s1 U2579 ( .DIN1(n2537), .DIN2(n2538), .DIN3(n2539), .DIN4(n2540), 
        .Q(n2536) );
  nnd2s1 U2580 ( .DIN1(n2137), .DIN2(n2028), .Q(n2540) );
  nnd2s1 U2581 ( .DIN1(n2021), .DIN2(n2030), .Q(n2539) );
  nnd2s1 U2582 ( .DIN1(n2065), .DIN2(n2049), .Q(n2538) );
  hi1s1 U2583 ( .DIN(n2143), .Q(n2065) );
  nnd2s1 U2584 ( .DIN1(n2019), .DIN2(n2029), .Q(n2537) );
  nnd3s1 U2585 ( .DIN1(n2541), .DIN2(n2542), .DIN3(n2543), .Q(n2535) );
  nnd2s1 U2586 ( .DIN1(n2109), .DIN2(n2544), .Q(n2543) );
  nnd3s1 U2587 ( .DIN1(n2526), .DIN2(n2147), .DIN3(n2206), .Q(n2544) );
  nnd2s1 U2588 ( .DIN1(n2032), .DIN2(n2545), .Q(n2542) );
  nnd2s1 U2589 ( .DIN1(n2205), .DIN2(n2291), .Q(n2545) );
  hi1s1 U2590 ( .DIN(n2070), .Q(n2032) );
  nnd2s1 U2591 ( .DIN1(n2134), .DIN2(n2546), .Q(n2541) );
  nnd2s1 U2592 ( .DIN1(n2043), .DIN2(n2277), .Q(n2546) );
  nor2s1 U2593 ( .DIN1(n2125), .DIN2(n2048), .Q(n2534) );
  and2s1 U2594 ( .DIN1(n2189), .DIN2(n2547), .Q(n2533) );
  nnd4s1 U2595 ( .DIN1(n2143), .DIN2(n2083), .DIN3(n2080), .DIN4(n2084), 
        .Q(n2547) );
  nnd3s1 U2596 ( .DIN1(n2548), .DIN2(n2549), .DIN3(n2550), .Q(n2495) );
  nnd2s1 U2597 ( .DIN1(n2077), .DIN2(n2028), .Q(n2550) );
  nnd2s1 U2598 ( .DIN1(n2326), .DIN2(n2027), .Q(n2549) );
  nnd2s1 U2599 ( .DIN1(n2107), .DIN2(n2066), .Q(n2548) );
  nnd4s1 U2600 ( .DIN1(n2551), .DIN2(n2552), .DIN3(n2553), .DIN4(n2554), 
        .Q(n2494) );
  nnd2s1 U2601 ( .DIN1(n2178), .DIN2(n2555), .Q(n2554) );
  nnd2s1 U2602 ( .DIN1(n2213), .DIN2(n2047), .Q(n2555) );
  nnd2s1 U2603 ( .DIN1(n2188), .DIN2(n2556), .Q(n2553) );
  nnd4s1 U2604 ( .DIN1(n2291), .DIN2(n2254), .DIN3(n2206), .DIN4(n2213), 
        .Q(n2556) );
  nnd2s1 U2605 ( .DIN1(n2144), .DIN2(n2295), .Q(n2552) );
  nnd2s1 U2606 ( .DIN1(n2261), .DIN2(n2044), .Q(n2295) );
  nnd2s1 U2607 ( .DIN1(n2029), .DIN2(n2198), .Q(n2551) );
  nnd2s1 U2608 ( .DIN1(n2070), .DIN2(n2079), .Q(n2198) );
  nor4s1 U2609 ( .DIN1(n2557), .DIN2(n2558), .DIN3(n2559), .DIN4(n2560), 
        .Q(n2014) );
  nnd4s1 U2610 ( .DIN1(n2561), .DIN2(n2562), .DIN3(n2563), .DIN4(n2564), 
        .Q(n2560) );
  nnd2s1 U2611 ( .DIN1(n2045), .DIN2(n2029), .Q(n2564) );
  nor2s1 U2612 ( .DIN1(n2565), .DIN2(n2290), .Q(n2563) );
  nor2s1 U2613 ( .DIN1(n2119), .DIN2(n2047), .Q(n2290) );
  nor2s1 U2614 ( .DIN1(n2105), .DIN2(n2147), .Q(n2565) );
  nnd2s1 U2615 ( .DIN1(n2028), .DIN2(n2134), .Q(n2562) );
  hi1s1 U2616 ( .DIN(n2044), .Q(n2028) );
  nnd2s1 U2617 ( .DIN1(n2117), .DIN2(n2120), .Q(n2561) );
  nnd3s1 U2618 ( .DIN1(n2566), .DIN2(n2567), .DIN3(n2568), .Q(n2559) );
  nnd2s1 U2619 ( .DIN1(n2110), .DIN2(n2196), .Q(n2568) );
  nnd2s1 U2620 ( .DIN1(n2116), .DIN2(n2105), .Q(n2196) );
  nnd2s1 U2621 ( .DIN1(n2030), .DIN2(n2569), .Q(n2567) );
  nnd3s1 U2622 ( .DIN1(n2206), .DIN2(n2213), .DIN3(n2254), .Q(n2569) );
  nnd2s1 U2623 ( .DIN1(n2108), .DIN2(n2570), .Q(n2566) );
  nnd3s1 U2624 ( .DIN1(n2526), .DIN2(n2208), .DIN3(n2253), .Q(n2570) );
  nor2s1 U2625 ( .DIN1(n2526), .DIN2(n2125), .Q(n2558) );
  nnd2s1 U2626 ( .DIN1(n2571), .DIN2(n2572), .Q(n2125) );
  nor2s1 U2627 ( .DIN1(n2362), .DIN2(n2277), .Q(n2557) );
  nor2s1 U2628 ( .DIN1(n2077), .DIN2(n2049), .Q(n2362) );
  nor4s1 U2629 ( .DIN1(n2573), .DIN2(n2574), .DIN3(n2575), .DIN4(n2576), 
        .Q(n2389) );
  nnd4s1 U2630 ( .DIN1(n2577), .DIN2(n2578), .DIN3(n2579), .DIN4(n2580), 
        .Q(n2576) );
  nnd2s1 U2631 ( .DIN1(n2117), .DIN2(n2166), .Q(n2580) );
  nor2s1 U2632 ( .DIN1(n2581), .DIN2(n2582), .Q(n2579) );
  nor2s1 U2633 ( .DIN1(n2048), .DIN2(n2116), .Q(n2582) );
  nor2s1 U2634 ( .DIN1(n2171), .DIN2(n2291), .Q(n2581) );
  nor2s1 U2635 ( .DIN1(n2045), .DIN2(n2166), .Q(n2171) );
  hi1s1 U2636 ( .DIN(n2119), .Q(n2166) );
  nnd2s1 U2637 ( .DIN1(n2022), .DIN2(n2029), .Q(n2578) );
  hi1s1 U2638 ( .DIN(n2084), .Q(n2022) );
  nnd2s1 U2639 ( .DIN1(n2326), .DIN2(n2110), .Q(n2577) );
  nnd3s1 U2640 ( .DIN1(n2583), .DIN2(n2584), .DIN3(n2585), .Q(n2575) );
  nnd2s1 U2641 ( .DIN1(n2020), .DIN2(n2232), .Q(n2585) );
  nnd2s1 U2642 ( .DIN1(n2079), .DIN2(n2177), .Q(n2232) );
  nnd2s1 U2643 ( .DIN1(n2066), .DIN2(n2586), .Q(n2584) );
  nnd2s1 U2644 ( .DIN1(n2253), .DIN2(n2123), .Q(n2586) );
  nnd2s1 U2645 ( .DIN1(n2108), .DIN2(n2587), .Q(n2583) );
  nnd2s1 U2646 ( .DIN1(n2040), .DIN2(n2291), .Q(n2587) );
  hi1s1 U2647 ( .DIN(n2080), .Q(n2108) );
  nor2s1 U2648 ( .DIN1(n2588), .DIN2(n2044), .Q(n2574) );
  nor2s1 U2649 ( .DIN1(n2021), .DIN2(n2107), .Q(n2588) );
  nor2s1 U2650 ( .DIN1(n2589), .DIN2(n2070), .Q(n2573) );
  nnd2s1 U2651 ( .DIN1(n2571), .DIN2(n2590), .Q(n2070) );
  nor2s1 U2652 ( .DIN1(n2027), .DIN2(n2077), .Q(n2589) );
  hi1s1 U2653 ( .DIN(n2234), .Q(n2077) );
  nnd3s1 U2654 ( .DIN1(w3[18]), .DIN2(n1558), .DIN3(n2591), .Q(n2234) );
  hi1s1 U2655 ( .DIN(n2048), .Q(n2027) );
  nnd4s1 U2656 ( .DIN1(n2398), .DIN2(n2592), .DIN3(n2593), .DIN4(n2594), 
        .Q(n2492) );
  nnd2s1 U2657 ( .DIN1(n2019), .DIN2(n2117), .Q(n2594) );
  hi1s1 U2658 ( .DIN(n2205), .Q(n2117) );
  hi1s1 U2659 ( .DIN(n2116), .Q(n2019) );
  nnd2s1 U2660 ( .DIN1(n2107), .DIN2(n2045), .Q(n2593) );
  nnd2s1 U2661 ( .DIN1(n2188), .DIN2(n2134), .Q(n2592) );
  hi1s1 U2662 ( .DIN(n2083), .Q(n2188) );
  and4s1 U2663 ( .DIN1(n2595), .DIN2(n2596), .DIN3(n2597), .DIN4(n2598), 
        .Q(n2398) );
  and4s1 U2664 ( .DIN1(n2599), .DIN2(n2306), .DIN3(n2600), .DIN4(n2601), 
        .Q(n2598) );
  nnd2s1 U2665 ( .DIN1(n2137), .DIN2(n2178), .Q(n2601) );
  nnd2s1 U2666 ( .DIN1(n2029), .DIN2(n2066), .Q(n2600) );
  hi1s1 U2667 ( .DIN(n2105), .Q(n2066) );
  hi1s1 U2668 ( .DIN(n2208), .Q(n2029) );
  nnd3s1 U2669 ( .DIN1(n1558), .DIN2(n1368), .DIN3(n2591), .Q(n2208) );
  nnd2s1 U2670 ( .DIN1(n2041), .DIN2(n2326), .Q(n2306) );
  hi1s1 U2671 ( .DIN(n2079), .Q(n2326) );
  nnd2s1 U2672 ( .DIN1(n2021), .DIN2(n2045), .Q(n2599) );
  hi1s1 U2673 ( .DIN(n2317), .Q(n2045) );
  nnd2s1 U2674 ( .DIN1(n2571), .DIN2(n2602), .Q(n2317) );
  and3s1 U2675 ( .DIN1(n2603), .DIN2(n2604), .DIN3(n2605), .Q(n2597) );
  nnd2s1 U2676 ( .DIN1(n2134), .DIN2(n2606), .Q(n2605) );
  nnd2s1 U2677 ( .DIN1(n2084), .DIN2(n2116), .Q(n2606) );
  hi1s1 U2678 ( .DIN(n2253), .Q(n2134) );
  nnd3s1 U2679 ( .DIN1(n2607), .DIN2(n1412), .DIN3(w3[16]), .Q(n2253) );
  nnd2s1 U2680 ( .DIN1(n2020), .DIN2(n2608), .Q(n2604) );
  nnd2s1 U2681 ( .DIN1(n2043), .DIN2(n2084), .Q(n2608) );
  nnd2s1 U2682 ( .DIN1(n2572), .DIN2(n2609), .Q(n2084) );
  hi1s1 U2683 ( .DIN(n2147), .Q(n2020) );
  nnd3s1 U2684 ( .DIN1(w3[16]), .DIN2(n1412), .DIN3(n2610), .Q(n2147) );
  nnd2s1 U2685 ( .DIN1(n2107), .DIN2(n2354), .Q(n2603) );
  nnd2s1 U2686 ( .DIN1(n2119), .DIN2(n2143), .Q(n2354) );
  hi1s1 U2687 ( .DIN(n2254), .Q(n2107) );
  nnd3s1 U2688 ( .DIN1(w3[16]), .DIN2(n2611), .DIN3(w3[18]), .Q(n2254) );
  nnd2s1 U2689 ( .DIN1(n2081), .DIN2(n2612), .Q(n2596) );
  nnd3s1 U2690 ( .DIN1(n2083), .DIN2(n2044), .DIN3(n2143), .Q(n2612) );
  nnd2s1 U2691 ( .DIN1(n2590), .DIN2(n2609), .Q(n2044) );
  nnd2s1 U2692 ( .DIN1(n2602), .DIN2(n2613), .Q(n2083) );
  hi1s1 U2693 ( .DIN(n2047), .Q(n2081) );
  nnd3s1 U2694 ( .DIN1(w3[18]), .DIN2(w3[16]), .DIN3(n2591), .Q(n2047) );
  or2s1 U2695 ( .DIN1(n2116), .DIN2(n2446), .Q(n2595) );
  nor2s1 U2696 ( .DIN1(n2031), .DIN2(n2049), .Q(n2446) );
  hi1s1 U2697 ( .DIN(n2526), .Q(n2049) );
  nnd3s1 U2698 ( .DIN1(n2611), .DIN2(n1368), .DIN3(w3[16]), .Q(n2526) );
  hi1s1 U2699 ( .DIN(n2040), .Q(n2031) );
  nnd3s1 U2700 ( .DIN1(n2607), .DIN2(n1558), .DIN3(w3[17]), .Q(n2040) );
  nnd4s1 U2701 ( .DIN1(n2221), .DIN2(n2614), .DIN3(n2615), .DIN4(n2616), 
        .Q(n2491) );
  nnd2s1 U2702 ( .DIN1(n2120), .DIN2(n2372), .Q(n2616) );
  nnd2s1 U2703 ( .DIN1(n2209), .DIN2(n2048), .Q(n2372) );
  nnd3s1 U2704 ( .DIN1(w3[17]), .DIN2(w3[16]), .DIN3(n2610), .Q(n2048) );
  hi1s1 U2705 ( .DIN(n2043), .Q(n2120) );
  nnd2s1 U2706 ( .DIN1(n2613), .DIN2(n2617), .Q(n2043) );
  nnd2s1 U2707 ( .DIN1(n2144), .DIN2(n2050), .Q(n2615) );
  nnd2s1 U2708 ( .DIN1(n2119), .DIN2(n2177), .Q(n2050) );
  nnd2s1 U2709 ( .DIN1(n2571), .DIN2(n2617), .Q(n2119) );
  nor2s1 U2710 ( .DIN1(n1376), .DIN2(w3[22]), .Q(n2571) );
  hi1s1 U2711 ( .DIN(n2209), .Q(n2144) );
  nnd3s1 U2712 ( .DIN1(n2611), .DIN2(n1558), .DIN3(w3[18]), .Q(n2209) );
  nnd2s1 U2713 ( .DIN1(n2178), .DIN2(n2110), .Q(n2614) );
  hi1s1 U2714 ( .DIN(n2277), .Q(n2178) );
  nnd2s1 U2715 ( .DIN1(n2602), .DIN2(n2618), .Q(n2277) );
  nnd2s1 U2716 ( .DIN1(n2137), .DIN2(n2030), .Q(n2221) );
  hi1s1 U2717 ( .DIN(n2177), .Q(n2030) );
  nnd2s1 U2718 ( .DIN1(n2609), .DIN2(n2617), .Q(n2177) );
  hi1s1 U2719 ( .DIN(n2291), .Q(n2137) );
  nnd3s1 U2720 ( .DIN1(w3[16]), .DIN2(n1368), .DIN3(n2591), .Q(n2291) );
  nor2s1 U2721 ( .DIN1(n1412), .DIN2(w3[19]), .Q(n2591) );
  nnd4s1 U2722 ( .DIN1(n2619), .DIN2(n2620), .DIN3(n2621), .DIN4(n2622), 
        .Q(n2490) );
  nnd2s1 U2723 ( .DIN1(n2021), .DIN2(n2623), .Q(n2622) );
  nnd2s1 U2724 ( .DIN1(n2080), .DIN2(n2105), .Q(n2623) );
  nnd2s1 U2725 ( .DIN1(n2572), .DIN2(n2618), .Q(n2105) );
  nnd2s1 U2726 ( .DIN1(n2618), .DIN2(n2617), .Q(n2080) );
  nor2s1 U2727 ( .DIN1(n1415), .DIN2(n1373), .Q(n2617) );
  hi1s1 U2728 ( .DIN(n2175), .Q(n2021) );
  nnd3s1 U2729 ( .DIN1(n1558), .DIN2(n1412), .DIN3(n2607), .Q(n2175) );
  nnd2s1 U2730 ( .DIN1(n2109), .DIN2(n2624), .Q(n2621) );
  nnd2s1 U2731 ( .DIN1(n2213), .DIN2(n2205), .Q(n2624) );
  nnd3s1 U2732 ( .DIN1(n1558), .DIN2(n1412), .DIN3(n2610), .Q(n2205) );
  hi1s1 U2733 ( .DIN(n2261), .Q(n2109) );
  nnd2s1 U2734 ( .DIN1(n2602), .DIN2(n2609), .Q(n2261) );
  nor2s1 U2735 ( .DIN1(n1438), .DIN2(w3[20]), .Q(n2609) );
  nor2s1 U2736 ( .DIN1(w3[23]), .DIN2(w3[21]), .Q(n2602) );
  or2s1 U2737 ( .DIN1(n2143), .DIN2(n2122), .Q(n2620) );
  nor2s1 U2738 ( .DIN1(n2041), .DIN2(n2110), .Q(n2122) );
  hi1s1 U2739 ( .DIN(n2206), .Q(n2110) );
  nnd3s1 U2740 ( .DIN1(w3[16]), .DIN2(n2607), .DIN3(w3[17]), .Q(n2206) );
  nor2s1 U2741 ( .DIN1(n1439), .DIN2(w3[18]), .Q(n2607) );
  hi1s1 U2742 ( .DIN(n2213), .Q(n2041) );
  nnd3s1 U2743 ( .DIN1(n1558), .DIN2(n1368), .DIN3(n2611), .Q(n2213) );
  nor2s1 U2744 ( .DIN1(w3[19]), .DIN2(w3[17]), .Q(n2611) );
  nnd2s1 U2745 ( .DIN1(n2590), .DIN2(n2618), .Q(n2143) );
  nor2s1 U2746 ( .DIN1(n1376), .DIN2(n1438), .Q(n2618) );
  nnd2s1 U2747 ( .DIN1(n2189), .DIN2(n2135), .Q(n2619) );
  nnd2s1 U2748 ( .DIN1(n2116), .DIN2(n2079), .Q(n2135) );
  nnd2s1 U2749 ( .DIN1(n2613), .DIN2(n2572), .Q(n2079) );
  nor2s1 U2750 ( .DIN1(n1415), .DIN2(w3[21]), .Q(n2572) );
  nnd2s1 U2751 ( .DIN1(n2590), .DIN2(n2613), .Q(n2116) );
  nor2s1 U2752 ( .DIN1(w3[22]), .DIN2(w3[20]), .Q(n2613) );
  nor2s1 U2753 ( .DIN1(n1373), .DIN2(w3[23]), .Q(n2590) );
  hi1s1 U2754 ( .DIN(n2123), .Q(n2189) );
  nnd3s1 U2755 ( .DIN1(w3[17]), .DIN2(n1558), .DIN3(n2610), .Q(n2123) );
  nor2s1 U2756 ( .DIN1(n1368), .DIN2(n1439), .Q(n2610) );
  xor2s1 U2757 ( .DIN1(n15581), .DIN2(w0[24]), .Q(n2488) );
  nnd2s1 U2758 ( .DIN1(n2625), .DIN2(n2626), .Q(\u0/N131 ) );
  nnd2s1 U2759 ( .DIN1(\key[87] ), .DIN2(ld), .Q(n2626) );
  nnd2s1 U2760 ( .DIN1(n1934), .DIN2(n1566), .Q(n2625) );
  xnr2s1 U2761 ( .DIN1(w1[23]), .DIN2(n1710), .Q(n1934) );
  xnr2s1 U2762 ( .DIN1(n1463), .DIN2(n2627), .Q(n1710) );
  nor4s1 U2763 ( .DIN1(n2628), .DIN2(n2629), .DIN3(n2630), .DIN4(n2631), 
        .Q(n2627) );
  nnd3s1 U2764 ( .DIN1(n2632), .DIN2(n2633), .DIN3(n2634), .Q(n2631) );
  nnd4s1 U2765 ( .DIN1(n2635), .DIN2(n2636), .DIN3(n2637), .DIN4(n2638), 
        .Q(n2630) );
  nnd2s1 U2766 ( .DIN1(n2639), .DIN2(n2640), .Q(n2637) );
  nnd2s1 U2767 ( .DIN1(n2641), .DIN2(n2642), .Q(n2636) );
  nnd4s1 U2768 ( .DIN1(n2643), .DIN2(n2644), .DIN3(n2645), .DIN4(n2646), 
        .Q(n2629) );
  nnd2s1 U2769 ( .DIN1(n2647), .DIN2(n2648), .Q(n2646) );
  nnd2s1 U2770 ( .DIN1(n2649), .DIN2(n2650), .Q(n2645) );
  nnd2s1 U2771 ( .DIN1(n2651), .DIN2(n2652), .Q(n2644) );
  nnd4s1 U2772 ( .DIN1(n2653), .DIN2(n2654), .DIN3(n2655), .DIN4(n2656), 
        .Q(n2628) );
  nnd2s1 U2773 ( .DIN1(n2657), .DIN2(n2658), .Q(n2656) );
  nnd2s1 U2774 ( .DIN1(n2659), .DIN2(n2660), .Q(n2658) );
  nnd2s1 U2775 ( .DIN1(n2661), .DIN2(n2662), .Q(n2655) );
  nnd2s1 U2776 ( .DIN1(n2663), .DIN2(n2664), .Q(n2662) );
  nnd2s1 U2777 ( .DIN1(n2665), .DIN2(n2666), .Q(n2654) );
  nnd2s1 U2778 ( .DIN1(n2667), .DIN2(n2668), .Q(n2666) );
  nnd2s1 U2779 ( .DIN1(n2669), .DIN2(n2670), .Q(n2653) );
  nnd2s1 U2780 ( .DIN1(n2671), .DIN2(n2672), .Q(\u0/N130 ) );
  nnd2s1 U2781 ( .DIN1(\key[86] ), .DIN2(ld), .Q(n2672) );
  nnd2s1 U2782 ( .DIN1(n1937), .DIN2(n1566), .Q(n2671) );
  xnr2s1 U2783 ( .DIN1(w1[22]), .DIN2(n1713), .Q(n1937) );
  xor2s1 U2784 ( .DIN1(w0[22]), .DIN2(n2673), .Q(n1713) );
  nor4s1 U2785 ( .DIN1(n2674), .DIN2(n2675), .DIN3(n2676), .DIN4(n2677), 
        .Q(n2673) );
  nnd3s1 U2786 ( .DIN1(n2678), .DIN2(n2679), .DIN3(n2680), .Q(n2677) );
  nnd3s1 U2787 ( .DIN1(n2681), .DIN2(n2682), .DIN3(n2683), .Q(n2676) );
  nnd2s1 U2788 ( .DIN1(n2684), .DIN2(n2649), .Q(n2682) );
  nnd3s1 U2789 ( .DIN1(n2685), .DIN2(n2686), .DIN3(n2687), .Q(n2675) );
  or2s1 U2790 ( .DIN1(n2688), .DIN2(n2689), .Q(n2687) );
  or2s1 U2791 ( .DIN1(n2664), .DIN2(n2690), .Q(n2686) );
  nnd2s1 U2792 ( .DIN1(n2665), .DIN2(n2691), .Q(n2685) );
  nnd3s1 U2793 ( .DIN1(n2692), .DIN2(n2693), .DIN3(n2694), .Q(n2674) );
  nnd2s1 U2794 ( .DIN1(n2695), .DIN2(n2696), .Q(n2694) );
  nnd2s1 U2795 ( .DIN1(n2697), .DIN2(n2698), .Q(n2696) );
  nnd2s1 U2796 ( .DIN1(n2699), .DIN2(n2700), .Q(n2693) );
  nnd2s1 U2797 ( .DIN1(n2701), .DIN2(n2702), .Q(n2700) );
  nnd2s1 U2798 ( .DIN1(n2641), .DIN2(n2703), .Q(n2692) );
  nnd2s1 U2799 ( .DIN1(n2704), .DIN2(n2705), .Q(n2703) );
  hi1s1 U2800 ( .DIN(n2706), .Q(n2705) );
  nnd2s1 U2801 ( .DIN1(n2707), .DIN2(n2708), .Q(\u0/N129 ) );
  nnd2s1 U2802 ( .DIN1(\key[85] ), .DIN2(ld), .Q(n2708) );
  nnd2s1 U2803 ( .DIN1(n1940), .DIN2(n1567), .Q(n2707) );
  xnr2s1 U2804 ( .DIN1(w1[21]), .DIN2(n1716), .Q(n1940) );
  xor2s1 U2805 ( .DIN1(w0[21]), .DIN2(n2709), .Q(n1716) );
  nor4s1 U2806 ( .DIN1(n2710), .DIN2(n2711), .DIN3(n2712), .DIN4(n2713), 
        .Q(n2709) );
  nnd3s1 U2807 ( .DIN1(n2714), .DIN2(n2679), .DIN3(n2715), .Q(n2713) );
  nor2s1 U2808 ( .DIN1(n2716), .DIN2(n2717), .Q(n2679) );
  nnd4s1 U2809 ( .DIN1(n2718), .DIN2(n2719), .DIN3(n2720), .DIN4(n2721), 
        .Q(n2717) );
  or2s1 U2810 ( .DIN1(n2722), .DIN2(n2723), .Q(n2721) );
  nnd2s1 U2811 ( .DIN1(n2724), .DIN2(n2725), .Q(n2720) );
  nnd2s1 U2812 ( .DIN1(n2726), .DIN2(n2640), .Q(n2719) );
  nnd2s1 U2813 ( .DIN1(n2652), .DIN2(n2727), .Q(n2718) );
  nnd4s1 U2814 ( .DIN1(n2728), .DIN2(n2729), .DIN3(n2730), .DIN4(n2731), 
        .Q(n2716) );
  nnd2s1 U2815 ( .DIN1(n2651), .DIN2(n2732), .Q(n2731) );
  nnd2s1 U2816 ( .DIN1(n2701), .DIN2(n2733), .Q(n2732) );
  nnd2s1 U2817 ( .DIN1(n2734), .DIN2(n2735), .Q(n2730) );
  nnd2s1 U2818 ( .DIN1(n2697), .DIN2(n2736), .Q(n2735) );
  nnd2s1 U2819 ( .DIN1(n2737), .DIN2(n2738), .Q(n2729) );
  nnd2s1 U2820 ( .DIN1(n2739), .DIN2(n2740), .Q(n2738) );
  nnd2s1 U2821 ( .DIN1(n2661), .DIN2(n2741), .Q(n2728) );
  nnd3s1 U2822 ( .DIN1(n2701), .DIN2(n2742), .DIN3(n2743), .Q(n2741) );
  nnd4s1 U2823 ( .DIN1(n2744), .DIN2(n2745), .DIN3(n2746), .DIN4(n2638), 
        .Q(n2712) );
  nnd2s1 U2824 ( .DIN1(n2726), .DIN2(n2699), .Q(n2638) );
  nnd2s1 U2825 ( .DIN1(n2695), .DIN2(n2737), .Q(n2746) );
  nnd2s1 U2826 ( .DIN1(n2724), .DIN2(n2642), .Q(n2745) );
  nnd4s1 U2827 ( .DIN1(n2747), .DIN2(n2748), .DIN3(n2749), .DIN4(n2750), 
        .Q(n2711) );
  nnd2s1 U2828 ( .DIN1(n2751), .DIN2(n2752), .Q(n2750) );
  nnd2s1 U2829 ( .DIN1(n2652), .DIN2(n2753), .Q(n2749) );
  nnd2s1 U2830 ( .DIN1(n2639), .DIN2(n2754), .Q(n2748) );
  nnd2s1 U2831 ( .DIN1(n2684), .DIN2(n2727), .Q(n2747) );
  nnd4s1 U2832 ( .DIN1(n2755), .DIN2(n2756), .DIN3(n2757), .DIN4(n2758), 
        .Q(n2710) );
  nnd2s1 U2833 ( .DIN1(n2669), .DIN2(n2759), .Q(n2758) );
  nnd2s1 U2834 ( .DIN1(n2698), .DIN2(n2760), .Q(n2759) );
  nnd2s1 U2835 ( .DIN1(n2761), .DIN2(n2762), .Q(n2757) );
  nnd2s1 U2836 ( .DIN1(n2665), .DIN2(n2763), .Q(n2756) );
  nnd2s1 U2837 ( .DIN1(n2764), .DIN2(n2660), .Q(n2763) );
  nnd2s1 U2838 ( .DIN1(n2649), .DIN2(n2765), .Q(n2755) );
  nnd2s1 U2839 ( .DIN1(n2766), .DIN2(n2767), .Q(\u0/N128 ) );
  nnd2s1 U2840 ( .DIN1(\key[84] ), .DIN2(ld), .Q(n2767) );
  nnd2s1 U2841 ( .DIN1(n1943), .DIN2(n1567), .Q(n2766) );
  xnr2s1 U2842 ( .DIN1(w1[20]), .DIN2(n1719), .Q(n1943) );
  xnr2s1 U2843 ( .DIN1(n1464), .DIN2(n2768), .Q(n1719) );
  nor4s1 U2844 ( .DIN1(n2769), .DIN2(n2770), .DIN3(n2771), .DIN4(n2772), 
        .Q(n2768) );
  nnd3s1 U2845 ( .DIN1(n2714), .DIN2(n2680), .DIN3(n2773), .Q(n2772) );
  nor4s1 U2846 ( .DIN1(n2774), .DIN2(n2775), .DIN3(n2776), .DIN4(n2777), 
        .Q(n2680) );
  nnd4s1 U2847 ( .DIN1(n2778), .DIN2(n2779), .DIN3(n2780), .DIN4(n2781), 
        .Q(n2777) );
  nnd2s1 U2848 ( .DIN1(n2647), .DIN2(n2684), .Q(n2781) );
  nnd2s1 U2849 ( .DIN1(n2724), .DIN2(n2782), .Q(n2779) );
  nnd2s1 U2850 ( .DIN1(n2734), .DIN2(n2648), .Q(n2778) );
  nnd3s1 U2851 ( .DIN1(n2783), .DIN2(n2784), .DIN3(n2785), .Q(n2776) );
  nnd2s1 U2852 ( .DIN1(n2751), .DIN2(n2786), .Q(n2785) );
  nnd2s1 U2853 ( .DIN1(n2787), .DIN2(n2663), .Q(n2786) );
  nnd2s1 U2854 ( .DIN1(n2661), .DIN2(n2788), .Q(n2784) );
  nnd2s1 U2855 ( .DIN1(n2789), .DIN2(n2760), .Q(n2788) );
  nnd2s1 U2856 ( .DIN1(n2726), .DIN2(n2790), .Q(n2783) );
  nnd2s1 U2857 ( .DIN1(n2791), .DIN2(n2660), .Q(n2790) );
  nor2s1 U2858 ( .DIN1(n2792), .DIN2(n2793), .Q(n2775) );
  and2s1 U2859 ( .DIN1(n2640), .DIN2(n2794), .Q(n2774) );
  nnd3s1 U2860 ( .DIN1(n2795), .DIN2(n2698), .DIN3(n2701), .Q(n2794) );
  nor3s1 U2861 ( .DIN1(n2796), .DIN2(n2797), .DIN3(n2798), .Q(n2714) );
  nnd4s1 U2862 ( .DIN1(n2678), .DIN2(n2799), .DIN3(n2800), .DIN4(n2801), 
        .Q(n2798) );
  and3s1 U2863 ( .DIN1(n2802), .DIN2(n2803), .DIN3(n2804), .Q(n2801) );
  nnd2s1 U2864 ( .DIN1(n2726), .DIN2(n2727), .Q(n2804) );
  nnd2s1 U2865 ( .DIN1(n2805), .DIN2(n2641), .Q(n2803) );
  nnd2s1 U2866 ( .DIN1(n2806), .DIN2(n2652), .Q(n2802) );
  nor2s1 U2867 ( .DIN1(n2807), .DIN2(n2808), .Q(n2678) );
  nnd4s1 U2868 ( .DIN1(n2809), .DIN2(n2810), .DIN3(n2811), .DIN4(n2812), 
        .Q(n2808) );
  nnd2s1 U2869 ( .DIN1(n2695), .DIN2(n2813), .Q(n2812) );
  nnd2s1 U2870 ( .DIN1(n2665), .DIN2(n2814), .Q(n2811) );
  nnd2s1 U2871 ( .DIN1(n2647), .DIN2(n2815), .Q(n2810) );
  nnd2s1 U2872 ( .DIN1(n2661), .DIN2(n2816), .Q(n2809) );
  nnd4s1 U2873 ( .DIN1(n2817), .DIN2(n2818), .DIN3(n2819), .DIN4(n2820), 
        .Q(n2807) );
  nnd2s1 U2874 ( .DIN1(n2684), .DIN2(n2814), .Q(n2820) );
  nnd2s1 U2875 ( .DIN1(n2651), .DIN2(n2821), .Q(n2819) );
  nnd2s1 U2876 ( .DIN1(n2702), .DIN2(n2736), .Q(n2821) );
  nnd2s1 U2877 ( .DIN1(n2639), .DIN2(n2822), .Q(n2818) );
  nnd2s1 U2878 ( .DIN1(n2823), .DIN2(n2824), .Q(n2822) );
  nnd2s1 U2879 ( .DIN1(n2805), .DIN2(n2825), .Q(n2817) );
  nnd3s1 U2880 ( .DIN1(n2668), .DIN2(n2826), .DIN3(n2827), .Q(n2825) );
  nnd3s1 U2881 ( .DIN1(n2828), .DIN2(n2829), .DIN3(n2643), .Q(n2797) );
  nnd2s1 U2882 ( .DIN1(n2734), .DIN2(n2725), .Q(n2643) );
  nnd2s1 U2883 ( .DIN1(n2639), .DIN2(n2830), .Q(n2829) );
  nnd3s1 U2884 ( .DIN1(n2740), .DIN2(n2831), .DIN3(n2690), .Q(n2830) );
  nor2s1 U2885 ( .DIN1(n2761), .DIN2(n2641), .Q(n2690) );
  nnd2s1 U2886 ( .DIN1(n2737), .DIN2(n2669), .Q(n2828) );
  nnd3s1 U2887 ( .DIN1(n2832), .DIN2(n2833), .DIN3(n2834), .Q(n2796) );
  nnd2s1 U2888 ( .DIN1(n2751), .DIN2(n2835), .Q(n2834) );
  nnd2s1 U2889 ( .DIN1(n2722), .DIN2(n2760), .Q(n2835) );
  nnd2s1 U2890 ( .DIN1(n2649), .DIN2(n2836), .Q(n2833) );
  nnd2s1 U2891 ( .DIN1(n2736), .DIN2(n2722), .Q(n2836) );
  nnd2s1 U2892 ( .DIN1(n2695), .DIN2(n2837), .Q(n2832) );
  nnd2s1 U2893 ( .DIN1(n2789), .DIN2(n2702), .Q(n2837) );
  nnd3s1 U2894 ( .DIN1(n2838), .DIN2(n2839), .DIN3(n2840), .Q(n2771) );
  nnd3s1 U2895 ( .DIN1(n2841), .DIN2(n2842), .DIN3(n2843), .Q(n2770) );
  nnd2s1 U2896 ( .DIN1(n2724), .DIN2(n2815), .Q(n2843) );
  nnd2s1 U2897 ( .DIN1(n2649), .DIN2(n2752), .Q(n2842) );
  nnd2s1 U2898 ( .DIN1(n2737), .DIN2(n2753), .Q(n2841) );
  nnd4s1 U2899 ( .DIN1(n2844), .DIN2(n2845), .DIN3(n2846), .DIN4(n2847), 
        .Q(n2769) );
  nnd2s1 U2900 ( .DIN1(n2647), .DIN2(n2848), .Q(n2847) );
  nnd2s1 U2901 ( .DIN1(n2733), .DIN2(n2698), .Q(n2848) );
  nnd2s1 U2902 ( .DIN1(n2684), .DIN2(n2849), .Q(n2846) );
  nnd2s1 U2903 ( .DIN1(n2827), .DIN2(n2823), .Q(n2849) );
  nnd2s1 U2904 ( .DIN1(n2699), .DIN2(n2850), .Q(n2845) );
  nnd2s1 U2905 ( .DIN1(n2657), .DIN2(n2851), .Q(n2844) );
  nnd2s1 U2906 ( .DIN1(n2852), .DIN2(n2824), .Q(n2851) );
  nnd2s1 U2907 ( .DIN1(n2853), .DIN2(n2854), .Q(\u0/N127 ) );
  nnd2s1 U2908 ( .DIN1(\key[83] ), .DIN2(ld), .Q(n2854) );
  nnd2s1 U2909 ( .DIN1(n1946), .DIN2(n1574), .Q(n2853) );
  xnr2s1 U2910 ( .DIN1(w1[19]), .DIN2(n1722), .Q(n1946) );
  xnr2s1 U2911 ( .DIN1(n1500), .DIN2(n2855), .Q(n1722) );
  nor4s1 U2912 ( .DIN1(n2856), .DIN2(n2857), .DIN3(n2858), .DIN4(n2859), 
        .Q(n2855) );
  nnd3s1 U2913 ( .DIN1(n2715), .DIN2(n2800), .DIN3(n2773), .Q(n2859) );
  nor4s1 U2914 ( .DIN1(n2860), .DIN2(n2861), .DIN3(n2862), .DIN4(n2863), 
        .Q(n2773) );
  nnd4s1 U2915 ( .DIN1(n2864), .DIN2(n2865), .DIN3(n2866), .DIN4(n2867), 
        .Q(n2863) );
  nor2s1 U2916 ( .DIN1(n2868), .DIN2(n2869), .Q(n2867) );
  nor2s1 U2917 ( .DIN1(n2870), .DIN2(n2823), .Q(n2869) );
  nor2s1 U2918 ( .DIN1(n2824), .DIN2(n2702), .Q(n2868) );
  nnd2s1 U2919 ( .DIN1(n2652), .DIN2(n2699), .Q(n2866) );
  nnd2s1 U2920 ( .DIN1(n2724), .DIN2(n2684), .Q(n2865) );
  nnd2s1 U2921 ( .DIN1(n2751), .DIN2(n2725), .Q(n2864) );
  nnd3s1 U2922 ( .DIN1(n2871), .DIN2(n2872), .DIN3(n2873), .Q(n2862) );
  nnd2s1 U2923 ( .DIN1(n2761), .DIN2(n2765), .Q(n2873) );
  nnd2s1 U2924 ( .DIN1(n2650), .DIN2(n2874), .Q(n2872) );
  nnd3s1 U2925 ( .DIN1(n2826), .DIN2(n2791), .DIN3(n2875), .Q(n2874) );
  nnd2s1 U2926 ( .DIN1(n2806), .DIN2(n2876), .Q(n2871) );
  nnd3s1 U2927 ( .DIN1(n2722), .DIN2(n2664), .DIN3(n2697), .Q(n2876) );
  nor2s1 U2928 ( .DIN1(n2722), .DIN2(n2668), .Q(n2861) );
  nor2s1 U2929 ( .DIN1(n2877), .DIN2(n2878), .Q(n2860) );
  nor4s1 U2930 ( .DIN1(n2879), .DIN2(n2880), .DIN3(n2881), .DIN4(n2882), 
        .Q(n2800) );
  nnd4s1 U2931 ( .DIN1(n2883), .DIN2(n2884), .DIN3(n2885), .DIN4(n2886), 
        .Q(n2882) );
  nor2s1 U2932 ( .DIN1(n2887), .DIN2(n2888), .Q(n2886) );
  nor2s1 U2933 ( .DIN1(n2875), .DIN2(n2878), .Q(n2888) );
  nor2s1 U2934 ( .DIN1(n2764), .DIN2(n2664), .Q(n2887) );
  nnd2s1 U2935 ( .DIN1(n2816), .DIN2(n2669), .Q(n2884) );
  nnd2s1 U2936 ( .DIN1(n2737), .DIN2(n2649), .Q(n2883) );
  nnd3s1 U2937 ( .DIN1(n2889), .DIN2(n2890), .DIN3(n2891), .Q(n2881) );
  nnd2s1 U2938 ( .DIN1(n2725), .DIN2(n2892), .Q(n2891) );
  nnd2s1 U2939 ( .DIN1(n2827), .DIN2(n2740), .Q(n2892) );
  nnd2s1 U2940 ( .DIN1(n2684), .DIN2(n2893), .Q(n2890) );
  nnd2s1 U2941 ( .DIN1(n2852), .DIN2(n2791), .Q(n2893) );
  nnd2s1 U2942 ( .DIN1(n2651), .DIN2(n2762), .Q(n2889) );
  nnd2s1 U2943 ( .DIN1(n2742), .DIN2(n2792), .Q(n2762) );
  nor2s1 U2944 ( .DIN1(n2894), .DIN2(n2702), .Q(n2880) );
  nor2s1 U2945 ( .DIN1(n2640), .DIN2(n2661), .Q(n2894) );
  nor2s1 U2946 ( .DIN1(n2895), .DIN2(n2824), .Q(n2879) );
  and2s1 U2947 ( .DIN1(n2722), .DIN2(n2896), .Q(n2895) );
  nor4s1 U2948 ( .DIN1(n2897), .DIN2(n2898), .DIN3(n2899), .DIN4(n2900), 
        .Q(n2715) );
  nnd4s1 U2949 ( .DIN1(n2901), .DIN2(n2902), .DIN3(n2903), .DIN4(n2904), 
        .Q(n2900) );
  nnd2s1 U2950 ( .DIN1(n2805), .DIN2(n2727), .Q(n2904) );
  nor2s1 U2951 ( .DIN1(n2905), .DIN2(n2906), .Q(n2903) );
  nor2s1 U2952 ( .DIN1(n2736), .DIN2(n2667), .Q(n2906) );
  nor2s1 U2953 ( .DIN1(n2702), .DIN2(n2907), .Q(n2905) );
  nnd2s1 U2954 ( .DIN1(n2726), .DIN2(n2734), .Q(n2902) );
  nnd2s1 U2955 ( .DIN1(n2724), .DIN2(n2657), .Q(n2901) );
  nnd3s1 U2956 ( .DIN1(n2908), .DIN2(n2909), .DIN3(n2910), .Q(n2899) );
  nnd2s1 U2957 ( .DIN1(n2649), .DIN2(n2911), .Q(n2910) );
  nnd2s1 U2958 ( .DIN1(n2665), .DIN2(n2912), .Q(n2909) );
  nnd2s1 U2959 ( .DIN1(n2824), .DIN2(n2791), .Q(n2912) );
  nnd2s1 U2960 ( .DIN1(n2806), .DIN2(n2913), .Q(n2908) );
  nnd3s1 U2961 ( .DIN1(n2795), .DIN2(n2878), .DIN3(n2914), .Q(n2913) );
  nor2s1 U2962 ( .DIN1(n2664), .DIN2(n2668), .Q(n2898) );
  nor2s1 U2963 ( .DIN1(n2704), .DIN2(n2660), .Q(n2897) );
  nnd3s1 U2964 ( .DIN1(n2915), .DIN2(n2916), .DIN3(n2683), .Q(n2858) );
  nor3s1 U2965 ( .DIN1(n2917), .DIN2(n2918), .DIN3(n2919), .Q(n2683) );
  nnd4s1 U2966 ( .DIN1(n2799), .DIN2(n2744), .DIN3(n2840), .DIN4(n2920), 
        .Q(n2919) );
  and3s1 U2967 ( .DIN1(n2921), .DIN2(n2922), .DIN3(n2923), .Q(n2920) );
  nnd2s1 U2968 ( .DIN1(n2724), .DIN2(n2648), .Q(n2923) );
  nnd2s1 U2969 ( .DIN1(n2639), .DIN2(n2699), .Q(n2921) );
  nor4s1 U2970 ( .DIN1(n2924), .DIN2(n2925), .DIN3(n2926), .DIN4(n2927), 
        .Q(n2840) );
  nnd4s1 U2971 ( .DIN1(n2928), .DIN2(n2929), .DIN3(n2930), .DIN4(n2931), 
        .Q(n2927) );
  nnd2s1 U2972 ( .DIN1(n2724), .DIN2(n2932), .Q(n2931) );
  nnd2s1 U2973 ( .DIN1(n2870), .DIN2(n2795), .Q(n2932) );
  nor2s1 U2974 ( .DIN1(n2933), .DIN2(n2934), .Q(n2930) );
  nor2s1 U2975 ( .DIN1(n2935), .DIN2(n2764), .Q(n2934) );
  nor2s1 U2976 ( .DIN1(n2639), .DIN2(n2706), .Q(n2935) );
  nor2s1 U2977 ( .DIN1(n2936), .DIN2(n2667), .Q(n2933) );
  nor2s1 U2978 ( .DIN1(n2937), .DIN2(n2737), .Q(n2936) );
  nnd2s1 U2979 ( .DIN1(n2657), .DIN2(n2938), .Q(n2929) );
  nnd3s1 U2980 ( .DIN1(n2668), .DIN2(n2823), .DIN3(n2907), .Q(n2938) );
  nnd2s1 U2981 ( .DIN1(n2806), .DIN2(n2937), .Q(n2928) );
  nnd3s1 U2982 ( .DIN1(n2939), .DIN2(n2940), .DIN3(n2941), .Q(n2926) );
  nnd2s1 U2983 ( .DIN1(n2942), .DIN2(n2761), .Q(n2941) );
  nnd2s1 U2984 ( .DIN1(n2647), .DIN2(n2650), .Q(n2940) );
  nnd2s1 U2985 ( .DIN1(n2651), .DIN2(n2684), .Q(n2939) );
  nor2s1 U2986 ( .DIN1(n2875), .DIN2(n2702), .Q(n2925) );
  nor2s1 U2987 ( .DIN1(n2878), .DIN2(n2852), .Q(n2924) );
  nor4s1 U2988 ( .DIN1(n2943), .DIN2(n2944), .DIN3(n2945), .DIN4(n2946), 
        .Q(n2744) );
  nnd4s1 U2989 ( .DIN1(n2947), .DIN2(n2948), .DIN3(n2949), .DIN4(n2950), 
        .Q(n2946) );
  nnd2s1 U2990 ( .DIN1(n2648), .DIN2(n2669), .Q(n2950) );
  nnd2s1 U2991 ( .DIN1(n2699), .DIN2(n2725), .Q(n2949) );
  nnd2s1 U2992 ( .DIN1(n2751), .DIN2(n2657), .Q(n2948) );
  nnd2s1 U2993 ( .DIN1(n2724), .DIN2(n2726), .Q(n2947) );
  nnd3s1 U2994 ( .DIN1(n2951), .DIN2(n2952), .DIN3(n2953), .Q(n2945) );
  nnd2s1 U2995 ( .DIN1(n2641), .DIN2(n2954), .Q(n2953) );
  nnd3s1 U2996 ( .DIN1(n2736), .DIN2(n2702), .DIN3(n2792), .Q(n2954) );
  nnd2s1 U2997 ( .DIN1(n2754), .DIN2(n2955), .Q(n2952) );
  nnd2s1 U2998 ( .DIN1(n2896), .DIN2(n2736), .Q(n2955) );
  nor2s1 U2999 ( .DIN1(n2942), .DIN2(n2937), .Q(n2896) );
  nnd2s1 U3000 ( .DIN1(n2805), .DIN2(n2956), .Q(n2951) );
  nnd2s1 U3001 ( .DIN1(n2957), .DIN2(n2852), .Q(n2956) );
  nor2s1 U3002 ( .DIN1(n2795), .DIN2(n2827), .Q(n2944) );
  nor2s1 U3003 ( .DIN1(n2743), .DIN2(n2824), .Q(n2943) );
  hi1s1 U3004 ( .DIN(n2670), .Q(n2743) );
  nor2s1 U3005 ( .DIN1(n2958), .DIN2(n2959), .Q(n2799) );
  nnd4s1 U3006 ( .DIN1(n2960), .DIN2(n2961), .DIN3(n2962), .DIN4(n2963), 
        .Q(n2959) );
  nnd2s1 U3007 ( .DIN1(n2648), .DIN2(n2964), .Q(n2963) );
  nnd3s1 U3008 ( .DIN1(n2824), .DIN2(n2875), .DIN3(n2907), .Q(n2964) );
  nnd2s1 U3009 ( .DIN1(n2647), .DIN2(n2737), .Q(n2961) );
  nnd4s1 U3010 ( .DIN1(n2965), .DIN2(n2966), .DIN3(n2967), .DIN4(n2968), 
        .Q(n2958) );
  nnd2s1 U3011 ( .DIN1(n2669), .DIN2(n2969), .Q(n2968) );
  nnd2s1 U3012 ( .DIN1(n2970), .DIN2(n2702), .Q(n2969) );
  nnd2s1 U3013 ( .DIN1(n2640), .DIN2(n2971), .Q(n2967) );
  nnd2s1 U3014 ( .DIN1(n2665), .DIN2(n2972), .Q(n2966) );
  nnd2s1 U3015 ( .DIN1(n2827), .DIN2(n2907), .Q(n2972) );
  nnd2s1 U3016 ( .DIN1(n2805), .DIN2(n2973), .Q(n2965) );
  nnd2s1 U3017 ( .DIN1(n2689), .DIN2(n2823), .Q(n2973) );
  nnd3s1 U3018 ( .DIN1(n2974), .DIN2(n2975), .DIN3(n2976), .Q(n2918) );
  nnd2s1 U3019 ( .DIN1(n2649), .DIN2(n2657), .Q(n2976) );
  nnd2s1 U3020 ( .DIN1(n2937), .DIN2(n2977), .Q(n2975) );
  nnd3s1 U3021 ( .DIN1(n2875), .DIN2(n2668), .DIN3(n2978), .Q(n2977) );
  or2s1 U3022 ( .DIN1(n2736), .DIN2(n2979), .Q(n2974) );
  nnd3s1 U3023 ( .DIN1(n2980), .DIN2(n2981), .DIN3(n2982), .Q(n2917) );
  nnd2s1 U3024 ( .DIN1(n2665), .DIN2(n2983), .Q(n2982) );
  nnd2s1 U3025 ( .DIN1(n2831), .DIN2(n2826), .Q(n2983) );
  nnd2s1 U3026 ( .DIN1(n2734), .DIN2(n2984), .Q(n2981) );
  or2s1 U3027 ( .DIN1(n2765), .DIN2(n2650), .Q(n2984) );
  nnd2s1 U3028 ( .DIN1(n2702), .DIN2(n2688), .Q(n2765) );
  nnd2s1 U3029 ( .DIN1(n2761), .DIN2(n2985), .Q(n2980) );
  nnd2s1 U3030 ( .DIN1(n2663), .DIN2(n2722), .Q(n2985) );
  nnd2s1 U3031 ( .DIN1(n2699), .DIN2(n2816), .Q(n2916) );
  nnd2s1 U3032 ( .DIN1(n2661), .DIN2(n2726), .Q(n2915) );
  nnd3s1 U3033 ( .DIN1(n2986), .DIN2(n2987), .DIN3(n2988), .Q(n2857) );
  nnd2s1 U3034 ( .DIN1(n2942), .DIN2(n2669), .Q(n2988) );
  nnd2s1 U3035 ( .DIN1(n2782), .DIN2(n2989), .Q(n2987) );
  nnd4s1 U3036 ( .DIN1(n2990), .DIN2(n2991), .DIN3(n2992), .DIN4(n2993), 
        .Q(n2856) );
  nnd2s1 U3037 ( .DIN1(n2754), .DIN2(n2994), .Q(n2993) );
  nnd2s1 U3038 ( .DIN1(n2704), .DIN2(n2760), .Q(n2994) );
  nor2s1 U3039 ( .DIN1(n2737), .DIN2(n2725), .Q(n2704) );
  nnd2s1 U3040 ( .DIN1(n2725), .DIN2(n2995), .Q(n2992) );
  nnd2s1 U3041 ( .DIN1(n2739), .DIN2(n2826), .Q(n2995) );
  nnd2s1 U3042 ( .DIN1(n2642), .DIN2(n2996), .Q(n2991) );
  nnd2s1 U3043 ( .DIN1(n2740), .DIN2(n2668), .Q(n2996) );
  nnd2s1 U3044 ( .DIN1(n2657), .DIN2(n2814), .Q(n2990) );
  nnd2s1 U3045 ( .DIN1(n2997), .DIN2(n2998), .Q(\u0/N126 ) );
  nnd2s1 U3046 ( .DIN1(\key[82] ), .DIN2(ld), .Q(n2998) );
  nnd2s1 U3047 ( .DIN1(n1949), .DIN2(n1567), .Q(n2997) );
  xnr2s1 U3048 ( .DIN1(w1[18]), .DIN2(n1725), .Q(n1949) );
  xnr2s1 U3049 ( .DIN1(n1465), .DIN2(n2999), .Q(n1725) );
  nor4s1 U3050 ( .DIN1(n3000), .DIN2(n3001), .DIN3(n3002), .DIN4(n3003), 
        .Q(n2999) );
  nnd3s1 U3051 ( .DIN1(n3004), .DIN2(n3005), .DIN3(n3006), .Q(n3003) );
  nnd3s1 U3052 ( .DIN1(n3007), .DIN2(n3008), .DIN3(n2635), .Q(n3002) );
  nor3s1 U3053 ( .DIN1(n3009), .DIN2(n3010), .DIN3(n3011), .Q(n2635) );
  nnd4s1 U3054 ( .DIN1(n3012), .DIN2(n3013), .DIN3(n3014), .DIN4(n3015), 
        .Q(n3011) );
  and3s1 U3055 ( .DIN1(n3016), .DIN2(n3017), .DIN3(n3018), .Q(n3015) );
  nnd2s1 U3056 ( .DIN1(n2695), .DIN2(n2642), .Q(n3018) );
  nnd2s1 U3057 ( .DIN1(n2647), .DIN2(n2726), .Q(n3017) );
  nnd2s1 U3058 ( .DIN1(n2661), .DIN2(n2725), .Q(n3016) );
  nnd3s1 U3059 ( .DIN1(n3019), .DIN2(n3020), .DIN3(n2962), .Q(n3010) );
  nnd2s1 U3060 ( .DIN1(n2724), .DIN2(n2937), .Q(n2962) );
  or2s1 U3061 ( .DIN1(n2667), .DIN2(n2970), .Q(n3020) );
  nor2s1 U3062 ( .DIN1(n2639), .DIN2(n2650), .Q(n2970) );
  nnd2s1 U3063 ( .DIN1(n2754), .DIN2(n2706), .Q(n3019) );
  nnd2s1 U3064 ( .DIN1(n2742), .DIN2(n2697), .Q(n2706) );
  nnd4s1 U3065 ( .DIN1(n3021), .DIN2(n3022), .DIN3(n3023), .DIN4(n3024), 
        .Q(n3009) );
  nnd2s1 U3066 ( .DIN1(n2782), .DIN2(n3025), .Q(n3024) );
  nnd2s1 U3067 ( .DIN1(n2641), .DIN2(n3026), .Q(n3023) );
  nnd2s1 U3068 ( .DIN1(n2697), .DIN2(n2760), .Q(n3026) );
  nnd2s1 U3069 ( .DIN1(n2737), .DIN2(n3027), .Q(n3022) );
  nnd2s1 U3070 ( .DIN1(n2740), .DIN2(n2660), .Q(n3027) );
  nnd2s1 U3071 ( .DIN1(n2665), .DIN2(n3028), .Q(n3021) );
  nnd2s1 U3072 ( .DIN1(n2978), .DIN2(n2875), .Q(n3028) );
  hi1s1 U3073 ( .DIN(n2753), .Q(n2978) );
  nnd2s1 U3074 ( .DIN1(n2823), .DIN2(n2764), .Q(n2753) );
  nnd2s1 U3075 ( .DIN1(n2661), .DIN2(n2652), .Q(n3008) );
  nnd2s1 U3076 ( .DIN1(n2657), .DIN2(n2727), .Q(n3007) );
  nnd3s1 U3077 ( .DIN1(n3029), .DIN2(n3030), .DIN3(n3031), .Q(n3001) );
  nnd2s1 U3078 ( .DIN1(n2726), .DIN2(n2649), .Q(n3031) );
  or2s1 U3079 ( .DIN1(n2663), .DIN2(n2659), .Q(n3030) );
  nor2s1 U3080 ( .DIN1(n2695), .DIN2(n2699), .Q(n2659) );
  nnd2s1 U3081 ( .DIN1(n2805), .DIN2(n2669), .Q(n3029) );
  nnd4s1 U3082 ( .DIN1(n3032), .DIN2(n3033), .DIN3(n3034), .DIN4(n3035), 
        .Q(n3000) );
  nnd2s1 U3083 ( .DIN1(n2942), .DIN2(n3036), .Q(n3035) );
  nnd2s1 U3084 ( .DIN1(n2979), .DIN2(n2823), .Q(n3036) );
  nnd2s1 U3085 ( .DIN1(n2640), .DIN2(n3037), .Q(n3034) );
  nnd2s1 U3086 ( .DIN1(n2789), .DIN2(n2698), .Q(n3037) );
  nor2s1 U3087 ( .DIN1(n2648), .DIN2(n2937), .Q(n2789) );
  nnd2s1 U3088 ( .DIN1(n2641), .DIN2(n3038), .Q(n3033) );
  nnd2s1 U3089 ( .DIN1(n2642), .DIN2(n3025), .Q(n3032) );
  nnd2s1 U3090 ( .DIN1(n2827), .DIN2(n2660), .Q(n3025) );
  nnd2s1 U3091 ( .DIN1(n3039), .DIN2(n3040), .Q(\u0/N125 ) );
  nnd2s1 U3092 ( .DIN1(\key[81] ), .DIN2(ld), .Q(n3040) );
  nnd2s1 U3093 ( .DIN1(n1952), .DIN2(n1567), .Q(n3039) );
  xnr2s1 U3094 ( .DIN1(w1[17]), .DIN2(n1728), .Q(n1952) );
  xnr2s1 U3095 ( .DIN1(n1501), .DIN2(n3041), .Q(n1728) );
  nor4s1 U3096 ( .DIN1(n3042), .DIN2(n3043), .DIN3(n3044), .DIN4(n3045), 
        .Q(n3041) );
  nnd3s1 U3097 ( .DIN1(n3006), .DIN2(n2632), .DIN3(n3046), .Q(n3045) );
  nor2s1 U3098 ( .DIN1(n3047), .DIN2(n3048), .Q(n2632) );
  nnd4s1 U3099 ( .DIN1(n3049), .DIN2(n3050), .DIN3(n3051), .DIN4(n3052), 
        .Q(n3048) );
  nnd2s1 U3100 ( .DIN1(n2652), .DIN2(n2814), .Q(n3052) );
  nnd2s1 U3101 ( .DIN1(n2740), .DIN2(n2667), .Q(n2814) );
  nnd2s1 U3102 ( .DIN1(n2648), .DIN2(n2649), .Q(n3051) );
  nnd2s1 U3103 ( .DIN1(n2641), .DIN2(n2737), .Q(n3050) );
  nnd2s1 U3104 ( .DIN1(n2805), .DIN2(n2761), .Q(n3049) );
  nnd4s1 U3105 ( .DIN1(n3053), .DIN2(n3054), .DIN3(n3055), .DIN4(n3056), 
        .Q(n3047) );
  nnd2s1 U3106 ( .DIN1(n2684), .DIN2(n3057), .Q(n3056) );
  or2s1 U3107 ( .DIN1(n2989), .DIN2(n2651), .Q(n3057) );
  nnd2s1 U3108 ( .DIN1(n2727), .DIN2(n3058), .Q(n3055) );
  nnd2s1 U3109 ( .DIN1(n2688), .DIN2(n2736), .Q(n3058) );
  nnd2s1 U3110 ( .DIN1(n2642), .DIN2(n3059), .Q(n3054) );
  nnd2s1 U3111 ( .DIN1(n2831), .DIN2(n2668), .Q(n3059) );
  nnd2s1 U3112 ( .DIN1(n2665), .DIN2(n3060), .Q(n3053) );
  nnd3s1 U3113 ( .DIN1(n2827), .DIN2(n2831), .DIN3(n3061), .Q(n3060) );
  nor4s1 U3114 ( .DIN1(n3062), .DIN2(n3063), .DIN3(n3064), .DIN4(n3065), 
        .Q(n3006) );
  nnd4s1 U3115 ( .DIN1(n3066), .DIN2(n2960), .DIN3(n3067), .DIN4(n3068), 
        .Q(n3065) );
  nnd2s1 U3116 ( .DIN1(n2751), .DIN2(n2670), .Q(n3068) );
  nnd2s1 U3117 ( .DIN1(n2754), .DIN2(n2642), .Q(n3067) );
  nnd2s1 U3118 ( .DIN1(n2651), .DIN2(n2942), .Q(n2960) );
  nnd2s1 U3119 ( .DIN1(n2695), .DIN2(n2782), .Q(n3066) );
  nnd3s1 U3120 ( .DIN1(n3069), .DIN2(n3070), .DIN3(n3071), .Q(n3064) );
  nnd2s1 U3121 ( .DIN1(n2657), .DIN2(n3072), .Q(n3071) );
  nnd2s1 U3122 ( .DIN1(n2647), .DIN2(n3073), .Q(n3070) );
  nnd2s1 U3123 ( .DIN1(n2701), .DIN2(n2698), .Q(n3073) );
  nnd2s1 U3124 ( .DIN1(n2816), .DIN2(n3074), .Q(n3069) );
  nnd2s1 U3125 ( .DIN1(n2689), .DIN2(n2667), .Q(n3074) );
  nor2s1 U3126 ( .DIN1(n2877), .DIN2(n2733), .Q(n3063) );
  nor2s1 U3127 ( .DIN1(n2761), .DIN2(n2754), .Q(n2877) );
  nor2s1 U3128 ( .DIN1(n3075), .DIN2(n2957), .Q(n3062) );
  nor2s1 U3129 ( .DIN1(n2737), .DIN2(n2726), .Q(n3075) );
  nnd3s1 U3130 ( .DIN1(n3076), .DIN2(n2838), .DIN3(n3013), .Q(n3044) );
  nor2s1 U3131 ( .DIN1(n3077), .DIN2(n3078), .Q(n3013) );
  nnd4s1 U3132 ( .DIN1(n3079), .DIN2(n3080), .DIN3(n2986), .DIN4(n3081), 
        .Q(n3078) );
  nnd2s1 U3133 ( .DIN1(n2816), .DIN2(n2691), .Q(n3081) );
  nnd2s1 U3134 ( .DIN1(n2852), .DIN2(n2668), .Q(n2691) );
  nnd2s1 U3135 ( .DIN1(n2695), .DIN2(n2650), .Q(n2986) );
  nnd2s1 U3136 ( .DIN1(n2806), .DIN2(n2782), .Q(n3080) );
  nnd2s1 U3137 ( .DIN1(n2642), .DIN2(n2699), .Q(n3079) );
  nnd4s1 U3138 ( .DIN1(n3082), .DIN2(n3083), .DIN3(n3084), .DIN4(n3085), 
        .Q(n3077) );
  nnd2s1 U3139 ( .DIN1(n2651), .DIN2(n3086), .Q(n3085) );
  nnd2s1 U3140 ( .DIN1(n2878), .DIN2(n2792), .Q(n3086) );
  nnd2s1 U3141 ( .DIN1(n2751), .DIN2(n3087), .Q(n3084) );
  nnd2s1 U3142 ( .DIN1(n2742), .DIN2(n2760), .Q(n3087) );
  nnd2s1 U3143 ( .DIN1(n2724), .DIN2(n3088), .Q(n3083) );
  nnd3s1 U3144 ( .DIN1(n2688), .DIN2(n2702), .DIN3(n2698), .Q(n3088) );
  nnd2s1 U3145 ( .DIN1(n2734), .DIN2(n3089), .Q(n3082) );
  nnd4s1 U3146 ( .DIN1(n2701), .DIN2(n2722), .DIN3(n2795), .DIN4(n2742), 
        .Q(n3089) );
  nnd2s1 U3147 ( .DIN1(n2652), .DIN2(n2751), .Q(n2838) );
  nnd2s1 U3148 ( .DIN1(n2806), .DIN2(n2665), .Q(n3076) );
  nnd3s1 U3149 ( .DIN1(n3090), .DIN2(n3091), .DIN3(n3092), .Q(n3043) );
  nnd2s1 U3150 ( .DIN1(n2695), .DIN2(n2725), .Q(n3092) );
  nnd2s1 U3151 ( .DIN1(n2651), .DIN2(n2648), .Q(n3091) );
  nnd2s1 U3152 ( .DIN1(n2782), .DIN2(n2640), .Q(n3090) );
  nnd4s1 U3153 ( .DIN1(n3093), .DIN2(n3094), .DIN3(n3095), .DIN4(n3096), 
        .Q(n3042) );
  nnd2s1 U3154 ( .DIN1(n2937), .DIN2(n3097), .Q(n3096) );
  nnd2s1 U3155 ( .DIN1(n2823), .DIN2(n2791), .Q(n3097) );
  nnd2s1 U3156 ( .DIN1(n2657), .DIN2(n3098), .Q(n3095) );
  nnd2s1 U3157 ( .DIN1(n2957), .DIN2(n2827), .Q(n3098) );
  nnd2s1 U3158 ( .DIN1(n2726), .DIN2(n3099), .Q(n3094) );
  nnd2s1 U3159 ( .DIN1(n2723), .DIN2(n2852), .Q(n3099) );
  nor2s1 U3160 ( .DIN1(n2641), .DIN2(n2754), .Q(n2723) );
  nnd2s1 U3161 ( .DIN1(n2737), .DIN2(n3100), .Q(n3093) );
  nnd3s1 U3162 ( .DIN1(n2824), .DIN2(n2826), .DIN3(n2689), .Q(n3100) );
  nor2s1 U3163 ( .DIN1(n2669), .DIN2(n2754), .Q(n2689) );
  nnd2s1 U3164 ( .DIN1(n3101), .DIN2(n3102), .Q(\u0/N124 ) );
  nnd2s1 U3165 ( .DIN1(\key[80] ), .DIN2(ld), .Q(n3102) );
  nnd2s1 U3166 ( .DIN1(n1955), .DIN2(n1567), .Q(n3101) );
  xnr2s1 U3167 ( .DIN1(w1[16]), .DIN2(n1731), .Q(n1955) );
  xnr2s1 U3168 ( .DIN1(n1466), .DIN2(n3103), .Q(n1731) );
  nor4s1 U3169 ( .DIN1(n3104), .DIN2(n3105), .DIN3(n3106), .DIN4(n3107), 
        .Q(n3103) );
  nnd3s1 U3170 ( .DIN1(n3005), .DIN2(n2634), .DIN3(n3046), .Q(n3107) );
  nor3s1 U3171 ( .DIN1(n3108), .DIN2(n3109), .DIN3(n3110), .Q(n3046) );
  nnd4s1 U3172 ( .DIN1(n2633), .DIN2(n3012), .DIN3(n3004), .DIN4(n3111), 
        .Q(n3110) );
  and3s1 U3173 ( .DIN1(n3112), .DIN2(n3113), .DIN3(n3114), .Q(n3111) );
  nnd2s1 U3174 ( .DIN1(n2726), .DIN2(n2751), .Q(n3114) );
  nnd2s1 U3175 ( .DIN1(n2642), .DIN2(n2734), .Q(n3113) );
  hi1s1 U3176 ( .DIN(n2702), .Q(n2642) );
  nnd2s1 U3177 ( .DIN1(n2806), .DIN2(n2657), .Q(n3112) );
  hi1s1 U3178 ( .DIN(n2742), .Q(n2657) );
  nor4s1 U3179 ( .DIN1(n3115), .DIN2(n3116), .DIN3(n3117), .DIN4(n3118), 
        .Q(n3004) );
  nnd4s1 U3180 ( .DIN1(n3119), .DIN2(n3120), .DIN3(n2885), .DIN4(n2780), 
        .Q(n3118) );
  nnd2s1 U3181 ( .DIN1(n2651), .DIN2(n2816), .Q(n2780) );
  nnd2s1 U3182 ( .DIN1(n2724), .DIN2(n2639), .Q(n2885) );
  nnd2s1 U3183 ( .DIN1(n2695), .DIN2(n2665), .Q(n3120) );
  nnd2s1 U3184 ( .DIN1(n2806), .DIN2(n2726), .Q(n3119) );
  nnd3s1 U3185 ( .DIN1(n3121), .DIN2(n3122), .DIN3(n3123), .Q(n3117) );
  nnd2s1 U3186 ( .DIN1(n2652), .DIN2(n3072), .Q(n3123) );
  nnd2s1 U3187 ( .DIN1(n2791), .DIN2(n2764), .Q(n3072) );
  nnd2s1 U3188 ( .DIN1(n2649), .DIN2(n3124), .Q(n3122) );
  nnd2s1 U3189 ( .DIN1(n2914), .DIN2(n2742), .Q(n3124) );
  nor2s1 U3190 ( .DIN1(n2805), .DIN2(n2782), .Q(n2914) );
  nnd2s1 U3191 ( .DIN1(n2942), .DIN2(n3125), .Q(n3121) );
  nnd2s1 U3192 ( .DIN1(n2827), .DIN2(n2667), .Q(n3125) );
  and2s1 U3193 ( .DIN1(n2727), .DIN2(n3126), .Q(n3116) );
  nnd3s1 U3194 ( .DIN1(n2664), .DIN2(n2702), .DIN3(n2698), .Q(n3126) );
  nor2s1 U3195 ( .DIN1(n3127), .DIN2(n2701), .Q(n3115) );
  nor2s1 U3196 ( .DIN1(n2651), .DIN2(n2695), .Q(n3127) );
  nor4s1 U3197 ( .DIN1(n3128), .DIN2(n3129), .DIN3(n3130), .DIN4(n3131), 
        .Q(n3012) );
  nnd4s1 U3198 ( .DIN1(n3132), .DIN2(n3133), .DIN3(n3134), .DIN4(n3135), 
        .Q(n3131) );
  and3s1 U3199 ( .DIN1(n3136), .DIN2(n3137), .DIN3(n3138), .Q(n3135) );
  nnd2s1 U3200 ( .DIN1(n2647), .DIN2(n2937), .Q(n3138) );
  nnd2s1 U3201 ( .DIN1(n2648), .DIN2(n3139), .Q(n3137) );
  nnd2s1 U3202 ( .DIN1(n2740), .DIN2(n2793), .Q(n3139) );
  nnd2s1 U3203 ( .DIN1(n2661), .DIN2(n3038), .Q(n3136) );
  nnd2s1 U3204 ( .DIN1(n2733), .DIN2(n2736), .Q(n3038) );
  nnd2s1 U3205 ( .DIN1(n2640), .DIN2(n3140), .Q(n3134) );
  nnd2s1 U3206 ( .DIN1(n2701), .DIN2(n2760), .Q(n3140) );
  nnd2s1 U3207 ( .DIN1(n2650), .DIN2(n3141), .Q(n3133) );
  nnd2s1 U3208 ( .DIN1(n2660), .DIN2(n2668), .Q(n3141) );
  nnd2s1 U3209 ( .DIN1(n2942), .DIN2(n3142), .Q(n3132) );
  nnd2s1 U3210 ( .DIN1(n2875), .DIN2(n2957), .Q(n3142) );
  nnd3s1 U3211 ( .DIN1(n3143), .DIN2(n3144), .DIN3(n3145), .Q(n3130) );
  nnd2s1 U3212 ( .DIN1(n2761), .DIN2(n2725), .Q(n3145) );
  nnd2s1 U3213 ( .DIN1(n2754), .DIN2(n2684), .Q(n3144) );
  nnd2s1 U3214 ( .DIN1(n2652), .DIN2(n2669), .Q(n3143) );
  nor2s1 U3215 ( .DIN1(n2824), .DIN2(n2870), .Q(n3129) );
  nor2s1 U3216 ( .DIN1(n2733), .DIN2(n2852), .Q(n3128) );
  nor4s1 U3217 ( .DIN1(n3146), .DIN2(n3147), .DIN3(n3148), .DIN4(n3149), 
        .Q(n2633) );
  nnd4s1 U3218 ( .DIN1(n3150), .DIN2(n3151), .DIN3(n3152), .DIN4(n3153), 
        .Q(n3149) );
  nnd2s1 U3219 ( .DIN1(n2754), .DIN2(n2648), .Q(n3153) );
  nnd2s1 U3220 ( .DIN1(n2641), .DIN2(n2650), .Q(n3152) );
  nnd2s1 U3221 ( .DIN1(n2684), .DIN2(n2669), .Q(n3151) );
  hi1s1 U3222 ( .DIN(n2760), .Q(n2684) );
  nnd2s1 U3223 ( .DIN1(n2639), .DIN2(n2649), .Q(n3150) );
  nnd3s1 U3224 ( .DIN1(n3154), .DIN2(n3155), .DIN3(n3156), .Q(n3148) );
  nnd2s1 U3225 ( .DIN1(n2726), .DIN2(n3157), .Q(n3156) );
  nnd3s1 U3226 ( .DIN1(n2793), .DIN2(n2764), .DIN3(n2824), .Q(n3157) );
  nnd2s1 U3227 ( .DIN1(n2652), .DIN2(n3158), .Q(n3155) );
  nnd2s1 U3228 ( .DIN1(n2823), .DIN2(n2907), .Q(n3158) );
  hi1s1 U3229 ( .DIN(n2688), .Q(n2652) );
  nnd2s1 U3230 ( .DIN1(n2751), .DIN2(n3159), .Q(n3154) );
  nnd2s1 U3231 ( .DIN1(n2663), .DIN2(n2792), .Q(n3159) );
  nor2s1 U3232 ( .DIN1(n2742), .DIN2(n2668), .Q(n3147) );
  and2s1 U3233 ( .DIN1(n2806), .DIN2(n3160), .Q(n3146) );
  nnd4s1 U3234 ( .DIN1(n2760), .DIN2(n2701), .DIN3(n2698), .DIN4(n2702), 
        .Q(n3160) );
  nnd3s1 U3235 ( .DIN1(n3161), .DIN2(n3162), .DIN3(n3163), .Q(n3109) );
  nnd2s1 U3236 ( .DIN1(n2695), .DIN2(n2648), .Q(n3163) );
  hi1s1 U3237 ( .DIN(n2664), .Q(n2648) );
  nnd2s1 U3238 ( .DIN1(n2942), .DIN2(n2647), .Q(n3162) );
  nnd2s1 U3239 ( .DIN1(n2724), .DIN2(n2816), .Q(n3161) );
  nnd4s1 U3240 ( .DIN1(n3164), .DIN2(n3165), .DIN3(n3166), .DIN4(n3167), 
        .Q(n3108) );
  nnd2s1 U3241 ( .DIN1(n2937), .DIN2(n3168), .Q(n3167) );
  nnd2s1 U3242 ( .DIN1(n2831), .DIN2(n2667), .Q(n3168) );
  nnd2s1 U3243 ( .DIN1(n2805), .DIN2(n3169), .Q(n3166) );
  nnd4s1 U3244 ( .DIN1(n2907), .DIN2(n2957), .DIN3(n2824), .DIN4(n2831), 
        .Q(n3169) );
  nnd2s1 U3245 ( .DIN1(n2761), .DIN2(n2911), .Q(n3165) );
  nnd2s1 U3246 ( .DIN1(n2878), .DIN2(n2664), .Q(n2911) );
  nnd2s1 U3247 ( .DIN1(n2649), .DIN2(n2815), .Q(n3164) );
  nnd2s1 U3248 ( .DIN1(n2688), .DIN2(n2697), .Q(n2815) );
  nor4s1 U3249 ( .DIN1(n3170), .DIN2(n3171), .DIN3(n3172), .DIN4(n3173), 
        .Q(n2634) );
  nnd4s1 U3250 ( .DIN1(n3174), .DIN2(n3175), .DIN3(n3176), .DIN4(n3177), 
        .Q(n3173) );
  nor2s1 U3251 ( .DIN1(n3178), .DIN2(n3179), .Q(n3177) );
  nor2s1 U3252 ( .DIN1(n2793), .DIN2(n2742), .Q(n3179) );
  nnd2s1 U3253 ( .DIN1(n3180), .DIN2(n3181), .Q(n2742) );
  nor2s1 U3254 ( .DIN1(n2979), .DIN2(n2792), .Q(n3178) );
  nor2s1 U3255 ( .DIN1(n2695), .DIN2(n2669), .Q(n2979) );
  nnd2s1 U3256 ( .DIN1(n2727), .DIN2(n2813), .Q(n3176) );
  nnd2s1 U3257 ( .DIN1(n2733), .DIN2(n2722), .Q(n2813) );
  nnd2s1 U3258 ( .DIN1(n2650), .DIN2(n3182), .Q(n3175) );
  nnd3s1 U3259 ( .DIN1(n2824), .DIN2(n2831), .DIN3(n2957), .Q(n3182) );
  nnd2s1 U3260 ( .DIN1(n2725), .DIN2(n3183), .Q(n3174) );
  nnd3s1 U3261 ( .DIN1(n2793), .DIN2(n2826), .DIN3(n2875), .Q(n3183) );
  nnd3s1 U3262 ( .DIN1(n3184), .DIN2(n2681), .DIN3(n3185), .Q(n3172) );
  nnd2s1 U3263 ( .DIN1(n2665), .DIN2(n2649), .Q(n3185) );
  nnd2s1 U3264 ( .DIN1(n2640), .DIN2(n2816), .Q(n2681) );
  nnd2s1 U3265 ( .DIN1(n2699), .DIN2(n2782), .Q(n3184) );
  nor2s1 U3266 ( .DIN1(n2663), .DIN2(n2823), .Q(n3171) );
  nor2s1 U3267 ( .DIN1(n2875), .DIN2(n2664), .Q(n3170) );
  nor4s1 U3268 ( .DIN1(n3186), .DIN2(n3187), .DIN3(n3188), .DIN4(n3189), 
        .Q(n3005) );
  nnd4s1 U3269 ( .DIN1(n3190), .DIN2(n3191), .DIN3(n3192), .DIN4(n3193), 
        .Q(n3189) );
  nor2s1 U3270 ( .DIN1(n3194), .DIN2(n3195), .Q(n3193) );
  nor2s1 U3271 ( .DIN1(n2824), .DIN2(n2697), .Q(n3195) );
  nor2s1 U3272 ( .DIN1(n2826), .DIN2(n2702), .Q(n3194) );
  nnd2s1 U3273 ( .DIN1(n2734), .DIN2(n2782), .Q(n3192) );
  or2s1 U3274 ( .DIN1(n2907), .DIN2(n2787), .Q(n3191) );
  nor2s1 U3275 ( .DIN1(n2665), .DIN2(n2782), .Q(n2787) );
  hi1s1 U3276 ( .DIN(n2736), .Q(n2782) );
  nnd2s1 U3277 ( .DIN1(n2639), .DIN2(n2647), .Q(n3190) );
  nnd3s1 U3278 ( .DIN1(n3196), .DIN2(n3197), .DIN3(n3198), .Q(n3188) );
  nnd2s1 U3279 ( .DIN1(n2640), .DIN2(n2850), .Q(n3198) );
  nnd2s1 U3280 ( .DIN1(n2697), .DIN2(n2795), .Q(n2850) );
  nnd2s1 U3281 ( .DIN1(n2816), .DIN2(n3199), .Q(n3197) );
  nnd2s1 U3282 ( .DIN1(n2875), .DIN2(n2740), .Q(n3199) );
  nnd2s1 U3283 ( .DIN1(n2725), .DIN2(n3200), .Q(n3196) );
  nnd2s1 U3284 ( .DIN1(n2660), .DIN2(n2907), .Q(n3200) );
  hi1s1 U3285 ( .DIN(n2698), .Q(n2725) );
  nor2s1 U3286 ( .DIN1(n3201), .DIN2(n2664), .Q(n3187) );
  nor2s1 U3287 ( .DIN1(n2641), .DIN2(n2724), .Q(n3201) );
  nor2s1 U3288 ( .DIN1(n3202), .DIN2(n2688), .Q(n3186) );
  nnd2s1 U3289 ( .DIN1(n3180), .DIN2(n3203), .Q(n2688) );
  nor2s1 U3290 ( .DIN1(n2647), .DIN2(n2695), .Q(n3202) );
  hi1s1 U3291 ( .DIN(n2852), .Q(n2695) );
  nnd3s1 U3292 ( .DIN1(w3[10]), .DIN2(n1361), .DIN3(n3204), .Q(n2852) );
  hi1s1 U3293 ( .DIN(n2668), .Q(n2647) );
  nnd4s1 U3294 ( .DIN1(n3014), .DIN2(n3205), .DIN3(n3206), .DIN4(n3207), 
        .Q(n3106) );
  nnd2s1 U3295 ( .DIN1(n2639), .DIN2(n2734), .Q(n3207) );
  hi1s1 U3296 ( .DIN(n2823), .Q(n2734) );
  hi1s1 U3297 ( .DIN(n2733), .Q(n2639) );
  nnd2s1 U3298 ( .DIN1(n2724), .DIN2(n2665), .Q(n3206) );
  nnd2s1 U3299 ( .DIN1(n2805), .DIN2(n2751), .Q(n3205) );
  hi1s1 U3300 ( .DIN(n2701), .Q(n2805) );
  nor4s1 U3301 ( .DIN1(n3208), .DIN2(n3209), .DIN3(n3210), .DIN4(n3211), 
        .Q(n3014) );
  nnd4s1 U3302 ( .DIN1(n3212), .DIN2(n2922), .DIN3(n3213), .DIN4(n3214), 
        .Q(n3211) );
  nnd2s1 U3303 ( .DIN1(n2754), .DIN2(n2937), .Q(n3214) );
  nnd2s1 U3304 ( .DIN1(n2649), .DIN2(n2816), .Q(n3213) );
  hi1s1 U3305 ( .DIN(n2722), .Q(n2816) );
  hi1s1 U3306 ( .DIN(n2826), .Q(n2649) );
  nnd3s1 U3307 ( .DIN1(n1553), .DIN2(n1361), .DIN3(n3204), .Q(n2826) );
  nnd2s1 U3308 ( .DIN1(n2661), .DIN2(n2942), .Q(n2922) );
  hi1s1 U3309 ( .DIN(n2697), .Q(n2942) );
  nnd2s1 U3310 ( .DIN1(n2641), .DIN2(n2665), .Q(n3212) );
  hi1s1 U3311 ( .DIN(n2870), .Q(n2665) );
  nnd2s1 U3312 ( .DIN1(n3180), .DIN2(n3215), .Q(n2870) );
  nnd3s1 U3313 ( .DIN1(n3216), .DIN2(n3217), .DIN3(n3218), .Q(n3210) );
  nnd2s1 U3314 ( .DIN1(n2751), .DIN2(n3219), .Q(n3218) );
  nnd2s1 U3315 ( .DIN1(n2702), .DIN2(n2733), .Q(n3219) );
  hi1s1 U3316 ( .DIN(n2875), .Q(n2751) );
  nnd2s1 U3317 ( .DIN1(n3220), .DIN2(n3221), .Q(n2875) );
  nnd2s1 U3318 ( .DIN1(n2640), .DIN2(n3222), .Q(n3217) );
  nnd2s1 U3319 ( .DIN1(n2663), .DIN2(n2702), .Q(n3222) );
  nnd2s1 U3320 ( .DIN1(n3181), .DIN2(n3223), .Q(n2702) );
  hi1s1 U3321 ( .DIN(n2764), .Q(n2640) );
  nnd2s1 U3322 ( .DIN1(n3224), .DIN2(n3220), .Q(n2764) );
  nnd2s1 U3323 ( .DIN1(n2724), .DIN2(n2971), .Q(n3216) );
  nnd2s1 U3324 ( .DIN1(n2736), .DIN2(n2760), .Q(n2971) );
  hi1s1 U3325 ( .DIN(n2957), .Q(n2724) );
  nnd3s1 U3326 ( .DIN1(w3[8]), .DIN2(n1413), .DIN3(n3224), .Q(n2957) );
  nor2s1 U3327 ( .DIN1(n3061), .DIN2(n2733), .Q(n3209) );
  nor2s1 U3328 ( .DIN1(n2651), .DIN2(n2669), .Q(n3061) );
  hi1s1 U3329 ( .DIN(n2793), .Q(n2669) );
  nnd3s1 U3330 ( .DIN1(n3221), .DIN2(n1413), .DIN3(w3[8]), .Q(n2793) );
  hi1s1 U3331 ( .DIN(n2660), .Q(n2651) );
  nnd3s1 U3332 ( .DIN1(w3[9]), .DIN2(n1553), .DIN3(n3225), .Q(n2660) );
  and2s1 U3333 ( .DIN1(n2699), .DIN2(n3226), .Q(n3208) );
  nnd3s1 U3334 ( .DIN1(n2701), .DIN2(n2664), .DIN3(n2760), .Q(n3226) );
  nnd2s1 U3335 ( .DIN1(n3203), .DIN2(n3223), .Q(n2664) );
  nnd2s1 U3336 ( .DIN1(n3215), .DIN2(n3227), .Q(n2701) );
  hi1s1 U3337 ( .DIN(n2667), .Q(n2699) );
  nnd3s1 U3338 ( .DIN1(w3[10]), .DIN2(w3[8]), .DIN3(n3204), .Q(n2667) );
  nnd4s1 U3339 ( .DIN1(n2839), .DIN2(n3228), .DIN3(n3229), .DIN4(n3230), 
        .Q(n3105) );
  nnd2s1 U3340 ( .DIN1(n2737), .DIN2(n2989), .Q(n3230) );
  nnd2s1 U3341 ( .DIN1(n2827), .DIN2(n2668), .Q(n2989) );
  nnd3s1 U3342 ( .DIN1(w3[9]), .DIN2(n3220), .DIN3(w3[10]), .Q(n2668) );
  hi1s1 U3343 ( .DIN(n2663), .Q(n2737) );
  nnd2s1 U3344 ( .DIN1(n3227), .DIN2(n3231), .Q(n2663) );
  nnd2s1 U3345 ( .DIN1(n2761), .DIN2(n2670), .Q(n3229) );
  nnd2s1 U3346 ( .DIN1(n2736), .DIN2(n2795), .Q(n2670) );
  nnd2s1 U3347 ( .DIN1(n3180), .DIN2(n3231), .Q(n2736) );
  nor2s1 U3348 ( .DIN1(n1393), .DIN2(w3[14]), .Q(n3180) );
  hi1s1 U3349 ( .DIN(n2827), .Q(n2761) );
  nnd3s1 U3350 ( .DIN1(n1413), .DIN2(n1361), .DIN3(n3224), .Q(n2827) );
  nnd2s1 U3351 ( .DIN1(n2937), .DIN2(n2727), .Q(n3228) );
  hi1s1 U3352 ( .DIN(n2792), .Q(n2937) );
  nnd2s1 U3353 ( .DIN1(n3215), .DIN2(n3232), .Q(n2792) );
  nnd2s1 U3354 ( .DIN1(n2754), .DIN2(n2650), .Q(n2839) );
  hi1s1 U3355 ( .DIN(n2795), .Q(n2650) );
  nnd2s1 U3356 ( .DIN1(n3223), .DIN2(n3231), .Q(n2795) );
  hi1s1 U3357 ( .DIN(n2907), .Q(n2754) );
  nnd3s1 U3358 ( .DIN1(w3[8]), .DIN2(n1553), .DIN3(n3204), .Q(n2907) );
  nor2s1 U3359 ( .DIN1(n1547), .DIN2(w3[11]), .Q(n3204) );
  nnd4s1 U3360 ( .DIN1(n3233), .DIN2(n3234), .DIN3(n3235), .DIN4(n3236), 
        .Q(n3104) );
  nnd2s1 U3361 ( .DIN1(n2641), .DIN2(n3237), .Q(n3236) );
  nnd2s1 U3362 ( .DIN1(n2698), .DIN2(n2722), .Q(n3237) );
  nnd2s1 U3363 ( .DIN1(n3181), .DIN2(n3232), .Q(n2722) );
  nnd2s1 U3364 ( .DIN1(n3232), .DIN2(n3231), .Q(n2698) );
  nor2s1 U3365 ( .DIN1(n1414), .DIN2(n1372), .Q(n3231) );
  hi1s1 U3366 ( .DIN(n2791), .Q(n2641) );
  nnd2s1 U3367 ( .DIN1(n3225), .DIN2(n3221), .Q(n2791) );
  nnd2s1 U3368 ( .DIN1(n2726), .DIN2(n3238), .Q(n3235) );
  nnd2s1 U3369 ( .DIN1(n2831), .DIN2(n2823), .Q(n3238) );
  nnd2s1 U3370 ( .DIN1(n3225), .DIN2(n3224), .Q(n2823) );
  nor2s1 U3371 ( .DIN1(n1553), .DIN2(w3[9]), .Q(n3224) );
  hi1s1 U3372 ( .DIN(n2878), .Q(n2726) );
  nnd2s1 U3373 ( .DIN1(n3215), .DIN2(n3223), .Q(n2878) );
  nor2s1 U3374 ( .DIN1(n1474), .DIN2(w3[12]), .Q(n3223) );
  nor2s1 U3375 ( .DIN1(w3[15]), .DIN2(w3[13]), .Q(n3215) );
  or2s1 U3376 ( .DIN1(n2760), .DIN2(n2739), .Q(n3234) );
  nor2s1 U3377 ( .DIN1(n2661), .DIN2(n2727), .Q(n2739) );
  hi1s1 U3378 ( .DIN(n2824), .Q(n2727) );
  nnd3s1 U3379 ( .DIN1(n3220), .DIN2(n1553), .DIN3(w3[9]), .Q(n2824) );
  nor2s1 U3380 ( .DIN1(n1361), .DIN2(n1413), .Q(n3220) );
  hi1s1 U3381 ( .DIN(n2831), .Q(n2661) );
  nnd3s1 U3382 ( .DIN1(n1413), .DIN2(n1361), .DIN3(n3221), .Q(n2831) );
  nor2s1 U3383 ( .DIN1(w3[9]), .DIN2(w3[10]), .Q(n3221) );
  nnd2s1 U3384 ( .DIN1(n3203), .DIN2(n3232), .Q(n2760) );
  nor2s1 U3385 ( .DIN1(n1393), .DIN2(n1474), .Q(n3232) );
  nnd2s1 U3386 ( .DIN1(n2806), .DIN2(n2752), .Q(n3233) );
  nnd2s1 U3387 ( .DIN1(n2733), .DIN2(n2697), .Q(n2752) );
  nnd2s1 U3388 ( .DIN1(n3227), .DIN2(n3181), .Q(n2697) );
  nor2s1 U3389 ( .DIN1(n1414), .DIN2(w3[13]), .Q(n3181) );
  nnd2s1 U3390 ( .DIN1(n3203), .DIN2(n3227), .Q(n2733) );
  nor2s1 U3391 ( .DIN1(w3[14]), .DIN2(w3[12]), .Q(n3227) );
  nor2s1 U3392 ( .DIN1(n1372), .DIN2(w3[15]), .Q(n3203) );
  hi1s1 U3393 ( .DIN(n2740), .Q(n2806) );
  nnd3s1 U3394 ( .DIN1(w3[10]), .DIN2(w3[9]), .DIN3(n3225), .Q(n2740) );
  nor2s1 U3395 ( .DIN1(n1413), .DIN2(w3[8]), .Q(n3225) );
  nnd2s1 U3396 ( .DIN1(n3239), .DIN2(n3240), .Q(\u0/N123 ) );
  nnd2s1 U3397 ( .DIN1(\key[79] ), .DIN2(ld), .Q(n3240) );
  nnd2s1 U3398 ( .DIN1(n1958), .DIN2(n1567), .Q(n3239) );
  xnr2s1 U3399 ( .DIN1(w1[15]), .DIN2(n1734), .Q(n1958) );
  xnr2s1 U3400 ( .DIN1(n1467), .DIN2(n3241), .Q(n1734) );
  nor4s1 U3401 ( .DIN1(n3242), .DIN2(n3243), .DIN3(n3244), .DIN4(n3245), 
        .Q(n3241) );
  nnd3s1 U3402 ( .DIN1(n3246), .DIN2(n3247), .DIN3(n3248), .Q(n3245) );
  nnd4s1 U3403 ( .DIN1(n3249), .DIN2(n3250), .DIN3(n3251), .DIN4(n3252), 
        .Q(n3244) );
  nnd2s1 U3404 ( .DIN1(n3253), .DIN2(n3254), .Q(n3251) );
  nnd2s1 U3405 ( .DIN1(n3255), .DIN2(n3256), .Q(n3250) );
  nnd4s1 U3406 ( .DIN1(n3257), .DIN2(n3258), .DIN3(n3259), .DIN4(n3260), 
        .Q(n3243) );
  nnd2s1 U3407 ( .DIN1(n3261), .DIN2(n3262), .Q(n3260) );
  nnd2s1 U3408 ( .DIN1(n3263), .DIN2(n3264), .Q(n3259) );
  nnd2s1 U3409 ( .DIN1(n3265), .DIN2(n3266), .Q(n3258) );
  nnd4s1 U3410 ( .DIN1(n3267), .DIN2(n3268), .DIN3(n3269), .DIN4(n3270), 
        .Q(n3242) );
  nnd2s1 U3411 ( .DIN1(n3271), .DIN2(n3272), .Q(n3270) );
  nnd2s1 U3412 ( .DIN1(n3273), .DIN2(n3274), .Q(n3272) );
  nnd2s1 U3413 ( .DIN1(n3275), .DIN2(n3276), .Q(n3269) );
  nnd2s1 U3414 ( .DIN1(n3277), .DIN2(n3278), .Q(n3276) );
  nnd2s1 U3415 ( .DIN1(n3279), .DIN2(n3280), .Q(n3268) );
  nnd2s1 U3416 ( .DIN1(n3281), .DIN2(n3282), .Q(n3280) );
  nnd2s1 U3417 ( .DIN1(n3283), .DIN2(n3284), .Q(n3267) );
  nnd2s1 U3418 ( .DIN1(n3285), .DIN2(n3286), .Q(\u0/N122 ) );
  nnd2s1 U3419 ( .DIN1(\key[78] ), .DIN2(ld), .Q(n3286) );
  nnd2s1 U3420 ( .DIN1(n1961), .DIN2(n1567), .Q(n3285) );
  xnr2s1 U3421 ( .DIN1(w1[14]), .DIN2(n1737), .Q(n1961) );
  xnr2s1 U3422 ( .DIN1(n1502), .DIN2(n3287), .Q(n1737) );
  nor4s1 U3423 ( .DIN1(n3288), .DIN2(n3289), .DIN3(n3290), .DIN4(n3291), 
        .Q(n3287) );
  nnd3s1 U3424 ( .DIN1(n3292), .DIN2(n3293), .DIN3(n3294), .Q(n3291) );
  nnd3s1 U3425 ( .DIN1(n3295), .DIN2(n3296), .DIN3(n3297), .Q(n3290) );
  nnd2s1 U3426 ( .DIN1(n3298), .DIN2(n3263), .Q(n3296) );
  nnd2s1 U3427 ( .DIN1(n3254), .DIN2(n3299), .Q(n3295) );
  nnd3s1 U3428 ( .DIN1(n3300), .DIN2(n3301), .DIN3(n3302), .Q(n3289) );
  or2s1 U3429 ( .DIN1(n3303), .DIN2(n3304), .Q(n3302) );
  or2s1 U3430 ( .DIN1(n3278), .DIN2(n3305), .Q(n3301) );
  nnd2s1 U3431 ( .DIN1(n3279), .DIN2(n3306), .Q(n3300) );
  nnd3s1 U3432 ( .DIN1(n3307), .DIN2(n3308), .DIN3(n3309), .Q(n3288) );
  nnd2s1 U3433 ( .DIN1(n3310), .DIN2(n3311), .Q(n3309) );
  nnd2s1 U3434 ( .DIN1(n3312), .DIN2(n3313), .Q(n3311) );
  nnd2s1 U3435 ( .DIN1(n3314), .DIN2(n3315), .Q(n3308) );
  nnd2s1 U3436 ( .DIN1(n3316), .DIN2(n3317), .Q(n3315) );
  nnd2s1 U3437 ( .DIN1(n3255), .DIN2(n3318), .Q(n3307) );
  nnd2s1 U3438 ( .DIN1(n3319), .DIN2(n3320), .Q(n3318) );
  hi1s1 U3439 ( .DIN(n3321), .Q(n3320) );
  nnd2s1 U3440 ( .DIN1(n3322), .DIN2(n3323), .Q(\u0/N121 ) );
  nnd2s1 U3441 ( .DIN1(\key[77] ), .DIN2(ld), .Q(n3323) );
  nnd2s1 U3442 ( .DIN1(n1964), .DIN2(n1568), .Q(n3322) );
  xnr2s1 U3443 ( .DIN1(w1[13]), .DIN2(n1740), .Q(n1964) );
  xnr2s1 U3444 ( .DIN1(n1468), .DIN2(n3324), .Q(n1740) );
  nor4s1 U3445 ( .DIN1(n3325), .DIN2(n3326), .DIN3(n3327), .DIN4(n3328), 
        .Q(n3324) );
  nnd3s1 U3446 ( .DIN1(n3329), .DIN2(n3293), .DIN3(n3330), .Q(n3328) );
  nor2s1 U3447 ( .DIN1(n3331), .DIN2(n3332), .Q(n3293) );
  nnd4s1 U3448 ( .DIN1(n3333), .DIN2(n3334), .DIN3(n3335), .DIN4(n3336), 
        .Q(n3332) );
  or2s1 U3449 ( .DIN1(n3337), .DIN2(n3338), .Q(n3336) );
  nnd2s1 U3450 ( .DIN1(n3339), .DIN2(n3340), .Q(n3335) );
  nnd2s1 U3451 ( .DIN1(n3341), .DIN2(n3254), .Q(n3334) );
  nnd2s1 U3452 ( .DIN1(n3266), .DIN2(n3342), .Q(n3333) );
  nnd4s1 U3453 ( .DIN1(n3343), .DIN2(n3344), .DIN3(n3345), .DIN4(n3346), 
        .Q(n3331) );
  nnd2s1 U3454 ( .DIN1(n3265), .DIN2(n3347), .Q(n3346) );
  nnd2s1 U3455 ( .DIN1(n3316), .DIN2(n3348), .Q(n3347) );
  nnd2s1 U3456 ( .DIN1(n3349), .DIN2(n3350), .Q(n3345) );
  nnd2s1 U3457 ( .DIN1(n3312), .DIN2(n3351), .Q(n3350) );
  nnd2s1 U3458 ( .DIN1(n3352), .DIN2(n3353), .Q(n3344) );
  nnd2s1 U3459 ( .DIN1(n3354), .DIN2(n3355), .Q(n3353) );
  nnd2s1 U3460 ( .DIN1(n3275), .DIN2(n3356), .Q(n3343) );
  nnd3s1 U3461 ( .DIN1(n3316), .DIN2(n3357), .DIN3(n3358), .Q(n3356) );
  nnd4s1 U3462 ( .DIN1(n3359), .DIN2(n3360), .DIN3(n3361), .DIN4(n3252), 
        .Q(n3327) );
  nnd2s1 U3463 ( .DIN1(n3341), .DIN2(n3314), .Q(n3252) );
  nnd2s1 U3464 ( .DIN1(n3310), .DIN2(n3352), .Q(n3361) );
  nnd2s1 U3465 ( .DIN1(n3339), .DIN2(n3256), .Q(n3360) );
  nnd4s1 U3466 ( .DIN1(n3362), .DIN2(n3363), .DIN3(n3364), .DIN4(n3365), 
        .Q(n3326) );
  nnd2s1 U3467 ( .DIN1(n3366), .DIN2(n3367), .Q(n3365) );
  nnd2s1 U3468 ( .DIN1(n3266), .DIN2(n3368), .Q(n3364) );
  nnd2s1 U3469 ( .DIN1(n3253), .DIN2(n3369), .Q(n3363) );
  nnd2s1 U3470 ( .DIN1(n3298), .DIN2(n3342), .Q(n3362) );
  nnd4s1 U3471 ( .DIN1(n3370), .DIN2(n3371), .DIN3(n3372), .DIN4(n3373), 
        .Q(n3325) );
  nnd2s1 U3472 ( .DIN1(n3283), .DIN2(n3374), .Q(n3373) );
  nnd2s1 U3473 ( .DIN1(n3313), .DIN2(n3375), .Q(n3374) );
  nnd2s1 U3474 ( .DIN1(n3376), .DIN2(n3377), .Q(n3372) );
  nnd2s1 U3475 ( .DIN1(n3279), .DIN2(n3378), .Q(n3371) );
  nnd2s1 U3476 ( .DIN1(n3379), .DIN2(n3274), .Q(n3378) );
  nnd2s1 U3477 ( .DIN1(n3263), .DIN2(n3380), .Q(n3370) );
  nnd2s1 U3478 ( .DIN1(n3381), .DIN2(n3382), .Q(\u0/N120 ) );
  nnd2s1 U3479 ( .DIN1(\key[76] ), .DIN2(ld), .Q(n3382) );
  nnd2s1 U3480 ( .DIN1(n1967), .DIN2(n1568), .Q(n3381) );
  xnr2s1 U3481 ( .DIN1(w1[12]), .DIN2(n1743), .Q(n1967) );
  xnr2s1 U3482 ( .DIN1(n1469), .DIN2(n3383), .Q(n1743) );
  nor4s1 U3483 ( .DIN1(n3384), .DIN2(n3385), .DIN3(n3386), .DIN4(n3387), 
        .Q(n3383) );
  nnd3s1 U3484 ( .DIN1(n3329), .DIN2(n3294), .DIN3(n3388), .Q(n3387) );
  and4s1 U3485 ( .DIN1(n3389), .DIN2(n3390), .DIN3(n3391), .DIN4(n3392), 
        .Q(n3294) );
  and4s1 U3486 ( .DIN1(n3393), .DIN2(n3394), .DIN3(n3395), .DIN4(n3396), 
        .Q(n3392) );
  nnd2s1 U3487 ( .DIN1(n3261), .DIN2(n3298), .Q(n3396) );
  nnd2s1 U3488 ( .DIN1(n3339), .DIN2(n3397), .Q(n3394) );
  nnd2s1 U3489 ( .DIN1(n3349), .DIN2(n3262), .Q(n3393) );
  and3s1 U3490 ( .DIN1(n3398), .DIN2(n3399), .DIN3(n3400), .Q(n3391) );
  nnd2s1 U3491 ( .DIN1(n3366), .DIN2(n3401), .Q(n3400) );
  nnd2s1 U3492 ( .DIN1(n3402), .DIN2(n3277), .Q(n3401) );
  nnd2s1 U3493 ( .DIN1(n3275), .DIN2(n3403), .Q(n3399) );
  nnd2s1 U3494 ( .DIN1(n3404), .DIN2(n3375), .Q(n3403) );
  nnd2s1 U3495 ( .DIN1(n3341), .DIN2(n3405), .Q(n3398) );
  nnd2s1 U3496 ( .DIN1(n3406), .DIN2(n3274), .Q(n3405) );
  nnd2s1 U3497 ( .DIN1(n3254), .DIN2(n3407), .Q(n3390) );
  nnd3s1 U3498 ( .DIN1(n3408), .DIN2(n3313), .DIN3(n3316), .Q(n3407) );
  nnd2s1 U3499 ( .DIN1(n3283), .DIN2(n3409), .Q(n3389) );
  nor3s1 U3500 ( .DIN1(n3410), .DIN2(n3411), .DIN3(n3412), .Q(n3329) );
  nnd4s1 U3501 ( .DIN1(n3292), .DIN2(n3413), .DIN3(n3414), .DIN4(n3415), 
        .Q(n3412) );
  and3s1 U3502 ( .DIN1(n3416), .DIN2(n3417), .DIN3(n3418), .Q(n3415) );
  nnd2s1 U3503 ( .DIN1(n3341), .DIN2(n3342), .Q(n3418) );
  nnd2s1 U3504 ( .DIN1(n3419), .DIN2(n3255), .Q(n3417) );
  nnd2s1 U3505 ( .DIN1(n3420), .DIN2(n3266), .Q(n3416) );
  nor2s1 U3506 ( .DIN1(n3421), .DIN2(n3422), .Q(n3292) );
  nnd4s1 U3507 ( .DIN1(n3423), .DIN2(n3424), .DIN3(n3425), .DIN4(n3426), 
        .Q(n3422) );
  nnd2s1 U3508 ( .DIN1(n3310), .DIN2(n3427), .Q(n3426) );
  nnd2s1 U3509 ( .DIN1(n3279), .DIN2(n3428), .Q(n3425) );
  nnd2s1 U3510 ( .DIN1(n3261), .DIN2(n3429), .Q(n3424) );
  nnd2s1 U3511 ( .DIN1(n3275), .DIN2(n3299), .Q(n3423) );
  nnd4s1 U3512 ( .DIN1(n3430), .DIN2(n3431), .DIN3(n3432), .DIN4(n3433), 
        .Q(n3421) );
  nnd2s1 U3513 ( .DIN1(n3298), .DIN2(n3428), .Q(n3433) );
  nnd2s1 U3514 ( .DIN1(n3265), .DIN2(n3434), .Q(n3432) );
  nnd2s1 U3515 ( .DIN1(n3317), .DIN2(n3351), .Q(n3434) );
  nnd2s1 U3516 ( .DIN1(n3253), .DIN2(n3435), .Q(n3431) );
  nnd2s1 U3517 ( .DIN1(n3436), .DIN2(n3437), .Q(n3435) );
  nnd2s1 U3518 ( .DIN1(n3419), .DIN2(n3438), .Q(n3430) );
  nnd3s1 U3519 ( .DIN1(n3282), .DIN2(n3439), .DIN3(n3440), .Q(n3438) );
  nnd3s1 U3520 ( .DIN1(n3441), .DIN2(n3442), .DIN3(n3257), .Q(n3411) );
  nnd2s1 U3521 ( .DIN1(n3349), .DIN2(n3340), .Q(n3257) );
  nnd2s1 U3522 ( .DIN1(n3253), .DIN2(n3443), .Q(n3442) );
  nnd3s1 U3523 ( .DIN1(n3355), .DIN2(n3444), .DIN3(n3305), .Q(n3443) );
  nor2s1 U3524 ( .DIN1(n3376), .DIN2(n3255), .Q(n3305) );
  nnd2s1 U3525 ( .DIN1(n3352), .DIN2(n3283), .Q(n3441) );
  nnd3s1 U3526 ( .DIN1(n3445), .DIN2(n3446), .DIN3(n3447), .Q(n3410) );
  nnd2s1 U3527 ( .DIN1(n3366), .DIN2(n3448), .Q(n3447) );
  nnd2s1 U3528 ( .DIN1(n3337), .DIN2(n3375), .Q(n3448) );
  nnd2s1 U3529 ( .DIN1(n3263), .DIN2(n3449), .Q(n3446) );
  nnd2s1 U3530 ( .DIN1(n3351), .DIN2(n3337), .Q(n3449) );
  nnd2s1 U3531 ( .DIN1(n3310), .DIN2(n3450), .Q(n3445) );
  nnd2s1 U3532 ( .DIN1(n3404), .DIN2(n3317), .Q(n3450) );
  nnd3s1 U3533 ( .DIN1(n3451), .DIN2(n3452), .DIN3(n3453), .Q(n3386) );
  nnd3s1 U3534 ( .DIN1(n3454), .DIN2(n3455), .DIN3(n3456), .Q(n3385) );
  nnd2s1 U3535 ( .DIN1(n3339), .DIN2(n3429), .Q(n3456) );
  nnd2s1 U3536 ( .DIN1(n3263), .DIN2(n3367), .Q(n3455) );
  nnd2s1 U3537 ( .DIN1(n3352), .DIN2(n3368), .Q(n3454) );
  nnd4s1 U3538 ( .DIN1(n3457), .DIN2(n3458), .DIN3(n3459), .DIN4(n3460), 
        .Q(n3384) );
  nnd2s1 U3539 ( .DIN1(n3261), .DIN2(n3461), .Q(n3460) );
  nnd2s1 U3540 ( .DIN1(n3348), .DIN2(n3313), .Q(n3461) );
  nnd2s1 U3541 ( .DIN1(n3298), .DIN2(n3462), .Q(n3459) );
  nnd2s1 U3542 ( .DIN1(n3440), .DIN2(n3436), .Q(n3462) );
  nnd2s1 U3543 ( .DIN1(n3314), .DIN2(n3463), .Q(n3458) );
  nnd2s1 U3544 ( .DIN1(n3271), .DIN2(n3464), .Q(n3457) );
  nnd2s1 U3545 ( .DIN1(n3465), .DIN2(n3437), .Q(n3464) );
  nnd2s1 U3546 ( .DIN1(n3466), .DIN2(n3467), .Q(\u0/N119 ) );
  nnd2s1 U3547 ( .DIN1(\key[75] ), .DIN2(ld), .Q(n3467) );
  nnd2s1 U3548 ( .DIN1(n1970), .DIN2(n1568), .Q(n3466) );
  xnr2s1 U3549 ( .DIN1(w1[11]), .DIN2(n1746), .Q(n1970) );
  xor2s1 U3550 ( .DIN1(w0[11]), .DIN2(n3468), .Q(n1746) );
  nor4s1 U3551 ( .DIN1(n3469), .DIN2(n3470), .DIN3(n3471), .DIN4(n3472), 
        .Q(n3468) );
  nnd3s1 U3552 ( .DIN1(n3330), .DIN2(n3414), .DIN3(n3388), .Q(n3472) );
  nor4s1 U3553 ( .DIN1(n3473), .DIN2(n3474), .DIN3(n3475), .DIN4(n3476), 
        .Q(n3388) );
  nnd4s1 U3554 ( .DIN1(n3477), .DIN2(n3478), .DIN3(n3479), .DIN4(n3480), 
        .Q(n3476) );
  nnd2s1 U3555 ( .DIN1(n3266), .DIN2(n3314), .Q(n3480) );
  nor2s1 U3556 ( .DIN1(n3481), .DIN2(n3482), .Q(n3479) );
  nor2s1 U3557 ( .DIN1(n3313), .DIN2(n3483), .Q(n3482) );
  nor2s1 U3558 ( .DIN1(n3375), .DIN2(n3484), .Q(n3481) );
  nnd2s1 U3559 ( .DIN1(n3256), .DIN2(n3342), .Q(n3478) );
  nnd2s1 U3560 ( .DIN1(n3349), .DIN2(n3279), .Q(n3477) );
  nnd3s1 U3561 ( .DIN1(n3485), .DIN2(n3486), .DIN3(n3487), .Q(n3475) );
  nnd2s1 U3562 ( .DIN1(n3376), .DIN2(n3380), .Q(n3487) );
  nnd2s1 U3563 ( .DIN1(n3264), .DIN2(n3488), .Q(n3486) );
  nnd3s1 U3564 ( .DIN1(n3439), .DIN2(n3406), .DIN3(n3483), .Q(n3488) );
  nnd2s1 U3565 ( .DIN1(n3420), .DIN2(n3489), .Q(n3485) );
  nnd3s1 U3566 ( .DIN1(n3337), .DIN2(n3278), .DIN3(n3312), .Q(n3489) );
  nor2s1 U3567 ( .DIN1(n3337), .DIN2(n3282), .Q(n3474) );
  nor2s1 U3568 ( .DIN1(n3490), .DIN2(n3491), .Q(n3473) );
  nor4s1 U3569 ( .DIN1(n3492), .DIN2(n3493), .DIN3(n3494), .DIN4(n3495), 
        .Q(n3414) );
  nnd4s1 U3570 ( .DIN1(n3496), .DIN2(n3497), .DIN3(n3498), .DIN4(n3499), 
        .Q(n3495) );
  nor2s1 U3571 ( .DIN1(n3500), .DIN2(n3501), .Q(n3499) );
  nor2s1 U3572 ( .DIN1(n3483), .DIN2(n3491), .Q(n3501) );
  nor2s1 U3573 ( .DIN1(n3379), .DIN2(n3278), .Q(n3500) );
  nnd2s1 U3574 ( .DIN1(n3299), .DIN2(n3283), .Q(n3497) );
  nnd2s1 U3575 ( .DIN1(n3352), .DIN2(n3263), .Q(n3496) );
  nnd3s1 U3576 ( .DIN1(n3502), .DIN2(n3503), .DIN3(n3504), .Q(n3494) );
  nnd2s1 U3577 ( .DIN1(n3340), .DIN2(n3505), .Q(n3504) );
  nnd2s1 U3578 ( .DIN1(n3440), .DIN2(n3355), .Q(n3505) );
  nnd2s1 U3579 ( .DIN1(n3298), .DIN2(n3506), .Q(n3503) );
  nnd2s1 U3580 ( .DIN1(n3465), .DIN2(n3406), .Q(n3506) );
  nnd2s1 U3581 ( .DIN1(n3265), .DIN2(n3377), .Q(n3502) );
  nnd2s1 U3582 ( .DIN1(n3357), .DIN2(n3507), .Q(n3377) );
  nor2s1 U3583 ( .DIN1(n3508), .DIN2(n3317), .Q(n3493) );
  nor2s1 U3584 ( .DIN1(n3254), .DIN2(n3275), .Q(n3508) );
  nor2s1 U3585 ( .DIN1(n3509), .DIN2(n3437), .Q(n3492) );
  and2s1 U3586 ( .DIN1(n3337), .DIN2(n3510), .Q(n3509) );
  nor4s1 U3587 ( .DIN1(n3511), .DIN2(n3512), .DIN3(n3513), .DIN4(n3514), 
        .Q(n3330) );
  nnd4s1 U3588 ( .DIN1(n3515), .DIN2(n3516), .DIN3(n3517), .DIN4(n3518), 
        .Q(n3514) );
  nnd2s1 U3589 ( .DIN1(n3419), .DIN2(n3342), .Q(n3518) );
  nor2s1 U3590 ( .DIN1(n3519), .DIN2(n3520), .Q(n3517) );
  nor2s1 U3591 ( .DIN1(n3317), .DIN2(n3521), .Q(n3519) );
  nnd2s1 U3592 ( .DIN1(n3341), .DIN2(n3349), .Q(n3516) );
  nnd2s1 U3593 ( .DIN1(n3339), .DIN2(n3271), .Q(n3515) );
  nnd3s1 U3594 ( .DIN1(n3522), .DIN2(n3523), .DIN3(n3524), .Q(n3513) );
  nnd2s1 U3595 ( .DIN1(n3263), .DIN2(n3525), .Q(n3524) );
  nnd2s1 U3596 ( .DIN1(n3279), .DIN2(n3526), .Q(n3523) );
  nnd2s1 U3597 ( .DIN1(n3437), .DIN2(n3406), .Q(n3526) );
  nnd2s1 U3598 ( .DIN1(n3420), .DIN2(n3527), .Q(n3522) );
  nnd3s1 U3599 ( .DIN1(n3408), .DIN2(n3491), .DIN3(n3528), .Q(n3527) );
  nor2s1 U3600 ( .DIN1(n3278), .DIN2(n3282), .Q(n3512) );
  nor2s1 U3601 ( .DIN1(n3319), .DIN2(n3274), .Q(n3511) );
  nnd3s1 U3602 ( .DIN1(n3529), .DIN2(n3530), .DIN3(n3297), .Q(n3471) );
  nor3s1 U3603 ( .DIN1(n3531), .DIN2(n3532), .DIN3(n3533), .Q(n3297) );
  nnd4s1 U3604 ( .DIN1(n3413), .DIN2(n3359), .DIN3(n3453), .DIN4(n3534), 
        .Q(n3533) );
  and3s1 U3605 ( .DIN1(n3535), .DIN2(n3536), .DIN3(n3537), .Q(n3534) );
  nnd2s1 U3606 ( .DIN1(n3339), .DIN2(n3262), .Q(n3537) );
  nnd2s1 U3607 ( .DIN1(n3253), .DIN2(n3314), .Q(n3535) );
  nor4s1 U3608 ( .DIN1(n3538), .DIN2(n3539), .DIN3(n3540), .DIN4(n3541), 
        .Q(n3453) );
  nnd4s1 U3609 ( .DIN1(n3542), .DIN2(n3543), .DIN3(n3544), .DIN4(n3545), 
        .Q(n3541) );
  nnd2s1 U3610 ( .DIN1(n3339), .DIN2(n3546), .Q(n3545) );
  nnd2s1 U3611 ( .DIN1(n3547), .DIN2(n3408), .Q(n3546) );
  nor2s1 U3612 ( .DIN1(n3548), .DIN2(n3549), .Q(n3544) );
  nor2s1 U3613 ( .DIN1(n3550), .DIN2(n3379), .Q(n3549) );
  nor2s1 U3614 ( .DIN1(n3253), .DIN2(n3321), .Q(n3550) );
  nor2s1 U3615 ( .DIN1(n3551), .DIN2(n3281), .Q(n3548) );
  nor2s1 U3616 ( .DIN1(n3409), .DIN2(n3352), .Q(n3551) );
  nnd2s1 U3617 ( .DIN1(n3271), .DIN2(n3552), .Q(n3543) );
  nnd3s1 U3618 ( .DIN1(n3282), .DIN2(n3436), .DIN3(n3521), .Q(n3552) );
  nnd2s1 U3619 ( .DIN1(n3420), .DIN2(n3409), .Q(n3542) );
  nnd3s1 U3620 ( .DIN1(n3553), .DIN2(n3554), .DIN3(n3555), .Q(n3540) );
  nnd2s1 U3621 ( .DIN1(n3556), .DIN2(n3376), .Q(n3555) );
  nnd2s1 U3622 ( .DIN1(n3261), .DIN2(n3264), .Q(n3554) );
  nnd2s1 U3623 ( .DIN1(n3265), .DIN2(n3298), .Q(n3553) );
  nor2s1 U3624 ( .DIN1(n3483), .DIN2(n3317), .Q(n3539) );
  nor2s1 U3625 ( .DIN1(n3491), .DIN2(n3465), .Q(n3538) );
  nor4s1 U3626 ( .DIN1(n3557), .DIN2(n3558), .DIN3(n3559), .DIN4(n3560), 
        .Q(n3359) );
  nnd4s1 U3627 ( .DIN1(n3561), .DIN2(n3562), .DIN3(n3563), .DIN4(n3564), 
        .Q(n3560) );
  nnd2s1 U3628 ( .DIN1(n3262), .DIN2(n3283), .Q(n3564) );
  nnd2s1 U3629 ( .DIN1(n3314), .DIN2(n3340), .Q(n3563) );
  nnd2s1 U3630 ( .DIN1(n3366), .DIN2(n3271), .Q(n3562) );
  nnd2s1 U3631 ( .DIN1(n3339), .DIN2(n3341), .Q(n3561) );
  nnd3s1 U3632 ( .DIN1(n3565), .DIN2(n3566), .DIN3(n3567), .Q(n3559) );
  nnd2s1 U3633 ( .DIN1(n3255), .DIN2(n3568), .Q(n3567) );
  nnd3s1 U3634 ( .DIN1(n3351), .DIN2(n3317), .DIN3(n3507), .Q(n3568) );
  nnd2s1 U3635 ( .DIN1(n3369), .DIN2(n3569), .Q(n3566) );
  nnd2s1 U3636 ( .DIN1(n3510), .DIN2(n3351), .Q(n3569) );
  nor2s1 U3637 ( .DIN1(n3556), .DIN2(n3409), .Q(n3510) );
  nnd2s1 U3638 ( .DIN1(n3419), .DIN2(n3570), .Q(n3565) );
  nnd2s1 U3639 ( .DIN1(n3484), .DIN2(n3465), .Q(n3570) );
  nor2s1 U3640 ( .DIN1(n3408), .DIN2(n3440), .Q(n3558) );
  nor2s1 U3641 ( .DIN1(n3358), .DIN2(n3437), .Q(n3557) );
  hi1s1 U3642 ( .DIN(n3284), .Q(n3358) );
  nor2s1 U3643 ( .DIN1(n3571), .DIN2(n3572), .Q(n3413) );
  nnd4s1 U3644 ( .DIN1(n3573), .DIN2(n3574), .DIN3(n3575), .DIN4(n3576), 
        .Q(n3572) );
  nnd2s1 U3645 ( .DIN1(n3262), .DIN2(n3577), .Q(n3576) );
  nnd3s1 U3646 ( .DIN1(n3437), .DIN2(n3483), .DIN3(n3521), .Q(n3577) );
  nnd2s1 U3647 ( .DIN1(n3261), .DIN2(n3352), .Q(n3574) );
  nnd4s1 U3648 ( .DIN1(n3578), .DIN2(n3579), .DIN3(n3580), .DIN4(n3581), 
        .Q(n3571) );
  nnd2s1 U3649 ( .DIN1(n3283), .DIN2(n3582), .Q(n3581) );
  nnd2s1 U3650 ( .DIN1(n3583), .DIN2(n3317), .Q(n3582) );
  nnd2s1 U3651 ( .DIN1(n3254), .DIN2(n3584), .Q(n3580) );
  nnd2s1 U3652 ( .DIN1(n3279), .DIN2(n3585), .Q(n3579) );
  nnd2s1 U3653 ( .DIN1(n3440), .DIN2(n3521), .Q(n3585) );
  nnd2s1 U3654 ( .DIN1(n3419), .DIN2(n3586), .Q(n3578) );
  nnd2s1 U3655 ( .DIN1(n3304), .DIN2(n3436), .Q(n3586) );
  nnd3s1 U3656 ( .DIN1(n3587), .DIN2(n3588), .DIN3(n3589), .Q(n3532) );
  nnd2s1 U3657 ( .DIN1(n3263), .DIN2(n3271), .Q(n3589) );
  nnd2s1 U3658 ( .DIN1(n3409), .DIN2(n3590), .Q(n3588) );
  nnd3s1 U3659 ( .DIN1(n3483), .DIN2(n3282), .DIN3(n3591), .Q(n3590) );
  or2s1 U3660 ( .DIN1(n3351), .DIN2(n3592), .Q(n3587) );
  nnd3s1 U3661 ( .DIN1(n3593), .DIN2(n3594), .DIN3(n3595), .Q(n3531) );
  nnd2s1 U3662 ( .DIN1(n3279), .DIN2(n3596), .Q(n3595) );
  nnd2s1 U3663 ( .DIN1(n3444), .DIN2(n3439), .Q(n3596) );
  nnd2s1 U3664 ( .DIN1(n3349), .DIN2(n3597), .Q(n3594) );
  or2s1 U3665 ( .DIN1(n3380), .DIN2(n3264), .Q(n3597) );
  nnd2s1 U3666 ( .DIN1(n3317), .DIN2(n3303), .Q(n3380) );
  nnd2s1 U3667 ( .DIN1(n3376), .DIN2(n3598), .Q(n3593) );
  nnd2s1 U3668 ( .DIN1(n3277), .DIN2(n3337), .Q(n3598) );
  nnd2s1 U3669 ( .DIN1(n3314), .DIN2(n3299), .Q(n3530) );
  nnd2s1 U3670 ( .DIN1(n3275), .DIN2(n3341), .Q(n3529) );
  nnd3s1 U3671 ( .DIN1(n3599), .DIN2(n3600), .DIN3(n3601), .Q(n3470) );
  nnd2s1 U3672 ( .DIN1(n3556), .DIN2(n3283), .Q(n3601) );
  nnd2s1 U3673 ( .DIN1(n3397), .DIN2(n3602), .Q(n3600) );
  nnd4s1 U3674 ( .DIN1(n3603), .DIN2(n3604), .DIN3(n3605), .DIN4(n3606), 
        .Q(n3469) );
  nnd2s1 U3675 ( .DIN1(n3369), .DIN2(n3607), .Q(n3606) );
  nnd2s1 U3676 ( .DIN1(n3319), .DIN2(n3375), .Q(n3607) );
  nor2s1 U3677 ( .DIN1(n3352), .DIN2(n3340), .Q(n3319) );
  nnd2s1 U3678 ( .DIN1(n3340), .DIN2(n3608), .Q(n3605) );
  nnd2s1 U3679 ( .DIN1(n3354), .DIN2(n3439), .Q(n3608) );
  nnd2s1 U3680 ( .DIN1(n3256), .DIN2(n3609), .Q(n3604) );
  nnd2s1 U3681 ( .DIN1(n3355), .DIN2(n3282), .Q(n3609) );
  nnd2s1 U3682 ( .DIN1(n3271), .DIN2(n3428), .Q(n3603) );
  nnd2s1 U3683 ( .DIN1(n3610), .DIN2(n3611), .Q(\u0/N118 ) );
  nnd2s1 U3684 ( .DIN1(\key[74] ), .DIN2(ld), .Q(n3611) );
  nnd2s1 U3685 ( .DIN1(n1973), .DIN2(n1568), .Q(n3610) );
  xnr2s1 U3686 ( .DIN1(w1[10]), .DIN2(n1749), .Q(n1973) );
  xnr2s1 U3687 ( .DIN1(n1499), .DIN2(n3612), .Q(n1749) );
  nor4s1 U3688 ( .DIN1(n3613), .DIN2(n3614), .DIN3(n3615), .DIN4(n3616), 
        .Q(n3612) );
  nnd3s1 U3689 ( .DIN1(n3617), .DIN2(n3618), .DIN3(n3619), .Q(n3616) );
  nnd3s1 U3690 ( .DIN1(n3620), .DIN2(n3621), .DIN3(n3249), .Q(n3615) );
  nor3s1 U3691 ( .DIN1(n3622), .DIN2(n3623), .DIN3(n3624), .Q(n3249) );
  nnd4s1 U3692 ( .DIN1(n3625), .DIN2(n3626), .DIN3(n3627), .DIN4(n3628), 
        .Q(n3624) );
  and3s1 U3693 ( .DIN1(n3629), .DIN2(n3630), .DIN3(n3631), .Q(n3628) );
  nnd2s1 U3694 ( .DIN1(n3310), .DIN2(n3256), .Q(n3631) );
  nnd2s1 U3695 ( .DIN1(n3261), .DIN2(n3341), .Q(n3630) );
  nnd2s1 U3696 ( .DIN1(n3275), .DIN2(n3340), .Q(n3629) );
  nnd3s1 U3697 ( .DIN1(n3632), .DIN2(n3633), .DIN3(n3575), .Q(n3623) );
  nnd2s1 U3698 ( .DIN1(n3339), .DIN2(n3409), .Q(n3575) );
  or2s1 U3699 ( .DIN1(n3281), .DIN2(n3583), .Q(n3633) );
  nor2s1 U3700 ( .DIN1(n3253), .DIN2(n3264), .Q(n3583) );
  nnd2s1 U3701 ( .DIN1(n3369), .DIN2(n3321), .Q(n3632) );
  nnd2s1 U3702 ( .DIN1(n3357), .DIN2(n3312), .Q(n3321) );
  nnd4s1 U3703 ( .DIN1(n3634), .DIN2(n3635), .DIN3(n3636), .DIN4(n3637), 
        .Q(n3622) );
  nnd2s1 U3704 ( .DIN1(n3397), .DIN2(n3638), .Q(n3637) );
  nnd2s1 U3705 ( .DIN1(n3255), .DIN2(n3639), .Q(n3636) );
  nnd2s1 U3706 ( .DIN1(n3312), .DIN2(n3375), .Q(n3639) );
  nnd2s1 U3707 ( .DIN1(n3352), .DIN2(n3640), .Q(n3635) );
  nnd2s1 U3708 ( .DIN1(n3355), .DIN2(n3274), .Q(n3640) );
  nnd2s1 U3709 ( .DIN1(n3279), .DIN2(n3641), .Q(n3634) );
  nnd2s1 U3710 ( .DIN1(n3591), .DIN2(n3483), .Q(n3641) );
  hi1s1 U3711 ( .DIN(n3368), .Q(n3591) );
  nnd2s1 U3712 ( .DIN1(n3436), .DIN2(n3379), .Q(n3368) );
  nnd2s1 U3713 ( .DIN1(n3275), .DIN2(n3266), .Q(n3621) );
  nnd2s1 U3714 ( .DIN1(n3271), .DIN2(n3342), .Q(n3620) );
  nnd3s1 U3715 ( .DIN1(n3642), .DIN2(n3643), .DIN3(n3644), .Q(n3614) );
  nnd2s1 U3716 ( .DIN1(n3341), .DIN2(n3263), .Q(n3644) );
  or2s1 U3717 ( .DIN1(n3277), .DIN2(n3273), .Q(n3643) );
  nor2s1 U3718 ( .DIN1(n3310), .DIN2(n3314), .Q(n3273) );
  nnd2s1 U3719 ( .DIN1(n3419), .DIN2(n3283), .Q(n3642) );
  nnd4s1 U3720 ( .DIN1(n3645), .DIN2(n3646), .DIN3(n3647), .DIN4(n3648), 
        .Q(n3613) );
  nnd2s1 U3721 ( .DIN1(n3556), .DIN2(n3649), .Q(n3648) );
  nnd2s1 U3722 ( .DIN1(n3592), .DIN2(n3436), .Q(n3649) );
  nnd2s1 U3723 ( .DIN1(n3254), .DIN2(n3650), .Q(n3647) );
  nnd2s1 U3724 ( .DIN1(n3404), .DIN2(n3313), .Q(n3650) );
  nor2s1 U3725 ( .DIN1(n3262), .DIN2(n3409), .Q(n3404) );
  nnd2s1 U3726 ( .DIN1(n3255), .DIN2(n3651), .Q(n3646) );
  nnd2s1 U3727 ( .DIN1(n3256), .DIN2(n3638), .Q(n3645) );
  nnd2s1 U3728 ( .DIN1(n3440), .DIN2(n3274), .Q(n3638) );
  nnd2s1 U3729 ( .DIN1(n3652), .DIN2(n3653), .Q(\u0/N117 ) );
  nnd2s1 U3730 ( .DIN1(\key[73] ), .DIN2(ld), .Q(n3653) );
  nnd2s1 U3731 ( .DIN1(n1976), .DIN2(n1568), .Q(n3652) );
  xnr2s1 U3732 ( .DIN1(w1[9]), .DIN2(n1752), .Q(n1976) );
  xnr2s1 U3733 ( .DIN1(n1503), .DIN2(n3654), .Q(n1752) );
  nor4s1 U3734 ( .DIN1(n3655), .DIN2(n3656), .DIN3(n3657), .DIN4(n3658), 
        .Q(n3654) );
  nnd3s1 U3735 ( .DIN1(n3619), .DIN2(n3246), .DIN3(n3659), .Q(n3658) );
  nor2s1 U3736 ( .DIN1(n3660), .DIN2(n3661), .Q(n3246) );
  nnd4s1 U3737 ( .DIN1(n3662), .DIN2(n3663), .DIN3(n3664), .DIN4(n3665), 
        .Q(n3661) );
  nnd2s1 U3738 ( .DIN1(n3266), .DIN2(n3428), .Q(n3665) );
  nnd2s1 U3739 ( .DIN1(n3355), .DIN2(n3281), .Q(n3428) );
  nnd2s1 U3740 ( .DIN1(n3262), .DIN2(n3263), .Q(n3664) );
  nnd2s1 U3741 ( .DIN1(n3255), .DIN2(n3352), .Q(n3663) );
  nnd2s1 U3742 ( .DIN1(n3419), .DIN2(n3376), .Q(n3662) );
  nnd4s1 U3743 ( .DIN1(n3666), .DIN2(n3667), .DIN3(n3668), .DIN4(n3669), 
        .Q(n3660) );
  nnd2s1 U3744 ( .DIN1(n3298), .DIN2(n3670), .Q(n3669) );
  or2s1 U3745 ( .DIN1(n3602), .DIN2(n3265), .Q(n3670) );
  nnd2s1 U3746 ( .DIN1(n3342), .DIN2(n3671), .Q(n3668) );
  nnd2s1 U3747 ( .DIN1(n3303), .DIN2(n3351), .Q(n3671) );
  nnd2s1 U3748 ( .DIN1(n3256), .DIN2(n3672), .Q(n3667) );
  nnd2s1 U3749 ( .DIN1(n3444), .DIN2(n3282), .Q(n3672) );
  nnd2s1 U3750 ( .DIN1(n3279), .DIN2(n3673), .Q(n3666) );
  nnd3s1 U3751 ( .DIN1(n3440), .DIN2(n3444), .DIN3(n3674), .Q(n3673) );
  nor4s1 U3752 ( .DIN1(n3675), .DIN2(n3676), .DIN3(n3677), .DIN4(n3678), 
        .Q(n3619) );
  nnd4s1 U3753 ( .DIN1(n3679), .DIN2(n3573), .DIN3(n3680), .DIN4(n3681), 
        .Q(n3678) );
  nnd2s1 U3754 ( .DIN1(n3366), .DIN2(n3284), .Q(n3681) );
  nnd2s1 U3755 ( .DIN1(n3369), .DIN2(n3256), .Q(n3680) );
  nnd2s1 U3756 ( .DIN1(n3265), .DIN2(n3556), .Q(n3573) );
  nnd2s1 U3757 ( .DIN1(n3310), .DIN2(n3397), .Q(n3679) );
  nnd3s1 U3758 ( .DIN1(n3682), .DIN2(n3683), .DIN3(n3684), .Q(n3677) );
  nnd2s1 U3759 ( .DIN1(n3271), .DIN2(n3685), .Q(n3684) );
  nnd2s1 U3760 ( .DIN1(n3261), .DIN2(n3686), .Q(n3683) );
  nnd2s1 U3761 ( .DIN1(n3316), .DIN2(n3313), .Q(n3686) );
  nnd2s1 U3762 ( .DIN1(n3299), .DIN2(n3687), .Q(n3682) );
  nnd2s1 U3763 ( .DIN1(n3304), .DIN2(n3281), .Q(n3687) );
  nor2s1 U3764 ( .DIN1(n3490), .DIN2(n3348), .Q(n3676) );
  nor2s1 U3765 ( .DIN1(n3376), .DIN2(n3369), .Q(n3490) );
  nor2s1 U3766 ( .DIN1(n3688), .DIN2(n3484), .Q(n3675) );
  nor2s1 U3767 ( .DIN1(n3352), .DIN2(n3341), .Q(n3688) );
  nnd3s1 U3768 ( .DIN1(n3689), .DIN2(n3451), .DIN3(n3626), .Q(n3657) );
  nor2s1 U3769 ( .DIN1(n3690), .DIN2(n3691), .Q(n3626) );
  nnd4s1 U3770 ( .DIN1(n3692), .DIN2(n3693), .DIN3(n3599), .DIN4(n3694), 
        .Q(n3691) );
  nnd2s1 U3771 ( .DIN1(n3299), .DIN2(n3306), .Q(n3694) );
  nnd2s1 U3772 ( .DIN1(n3465), .DIN2(n3282), .Q(n3306) );
  nnd2s1 U3773 ( .DIN1(n3310), .DIN2(n3264), .Q(n3599) );
  nnd2s1 U3774 ( .DIN1(n3420), .DIN2(n3397), .Q(n3693) );
  nnd2s1 U3775 ( .DIN1(n3256), .DIN2(n3314), .Q(n3692) );
  nnd4s1 U3776 ( .DIN1(n3695), .DIN2(n3696), .DIN3(n3697), .DIN4(n3698), 
        .Q(n3690) );
  nnd2s1 U3777 ( .DIN1(n3265), .DIN2(n3699), .Q(n3698) );
  nnd2s1 U3778 ( .DIN1(n3491), .DIN2(n3507), .Q(n3699) );
  nnd2s1 U3779 ( .DIN1(n3366), .DIN2(n3700), .Q(n3697) );
  nnd2s1 U3780 ( .DIN1(n3357), .DIN2(n3375), .Q(n3700) );
  nnd2s1 U3781 ( .DIN1(n3339), .DIN2(n3701), .Q(n3696) );
  nnd3s1 U3782 ( .DIN1(n3303), .DIN2(n3317), .DIN3(n3313), .Q(n3701) );
  nnd2s1 U3783 ( .DIN1(n3349), .DIN2(n3702), .Q(n3695) );
  nnd4s1 U3784 ( .DIN1(n3316), .DIN2(n3337), .DIN3(n3408), .DIN4(n3357), 
        .Q(n3702) );
  nnd2s1 U3785 ( .DIN1(n3266), .DIN2(n3366), .Q(n3451) );
  nnd2s1 U3786 ( .DIN1(n3420), .DIN2(n3279), .Q(n3689) );
  nnd3s1 U3787 ( .DIN1(n3703), .DIN2(n3704), .DIN3(n3705), .Q(n3656) );
  nnd2s1 U3788 ( .DIN1(n3310), .DIN2(n3340), .Q(n3705) );
  nnd2s1 U3789 ( .DIN1(n3265), .DIN2(n3262), .Q(n3704) );
  nnd2s1 U3790 ( .DIN1(n3397), .DIN2(n3254), .Q(n3703) );
  nnd4s1 U3791 ( .DIN1(n3706), .DIN2(n3707), .DIN3(n3708), .DIN4(n3709), 
        .Q(n3655) );
  nnd2s1 U3792 ( .DIN1(n3409), .DIN2(n3710), .Q(n3709) );
  nnd2s1 U3793 ( .DIN1(n3436), .DIN2(n3406), .Q(n3710) );
  nnd2s1 U3794 ( .DIN1(n3271), .DIN2(n3711), .Q(n3708) );
  nnd2s1 U3795 ( .DIN1(n3484), .DIN2(n3440), .Q(n3711) );
  nnd2s1 U3796 ( .DIN1(n3341), .DIN2(n3712), .Q(n3707) );
  nnd2s1 U3797 ( .DIN1(n3338), .DIN2(n3465), .Q(n3712) );
  nor2s1 U3798 ( .DIN1(n3255), .DIN2(n3369), .Q(n3338) );
  nnd2s1 U3799 ( .DIN1(n3352), .DIN2(n3713), .Q(n3706) );
  nnd3s1 U3800 ( .DIN1(n3437), .DIN2(n3439), .DIN3(n3304), .Q(n3713) );
  nor2s1 U3801 ( .DIN1(n3283), .DIN2(n3369), .Q(n3304) );
  nnd2s1 U3802 ( .DIN1(n3714), .DIN2(n3715), .Q(\u0/N116 ) );
  nnd2s1 U3803 ( .DIN1(\key[72] ), .DIN2(ld), .Q(n3715) );
  nnd2s1 U3804 ( .DIN1(n1979), .DIN2(n1568), .Q(n3714) );
  xnr2s1 U3805 ( .DIN1(w1[8]), .DIN2(n1755), .Q(n1979) );
  xnr2s1 U3806 ( .DIN1(n1470), .DIN2(n3716), .Q(n1755) );
  nor4s1 U3807 ( .DIN1(n3717), .DIN2(n3718), .DIN3(n3719), .DIN4(n3720), 
        .Q(n3716) );
  nnd3s1 U3808 ( .DIN1(n3618), .DIN2(n3248), .DIN3(n3659), .Q(n3720) );
  nor3s1 U3809 ( .DIN1(n3721), .DIN2(n3722), .DIN3(n3723), .Q(n3659) );
  nnd4s1 U3810 ( .DIN1(n3247), .DIN2(n3625), .DIN3(n3617), .DIN4(n3724), 
        .Q(n3723) );
  and3s1 U3811 ( .DIN1(n3725), .DIN2(n3726), .DIN3(n3727), .Q(n3724) );
  nnd2s1 U3812 ( .DIN1(n3341), .DIN2(n3366), .Q(n3727) );
  nnd2s1 U3813 ( .DIN1(n3256), .DIN2(n3349), .Q(n3726) );
  nnd2s1 U3814 ( .DIN1(n3420), .DIN2(n3271), .Q(n3725) );
  hi1s1 U3815 ( .DIN(n3357), .Q(n3271) );
  and4s1 U3816 ( .DIN1(n3728), .DIN2(n3729), .DIN3(n3730), .DIN4(n3731), 
        .Q(n3617) );
  and4s1 U3817 ( .DIN1(n3732), .DIN2(n3733), .DIN3(n3498), .DIN4(n3395), 
        .Q(n3731) );
  nnd2s1 U3818 ( .DIN1(n3265), .DIN2(n3299), .Q(n3395) );
  nnd2s1 U3819 ( .DIN1(n3339), .DIN2(n3253), .Q(n3498) );
  nnd2s1 U3820 ( .DIN1(n3310), .DIN2(n3279), .Q(n3733) );
  nnd2s1 U3821 ( .DIN1(n3420), .DIN2(n3341), .Q(n3732) );
  and3s1 U3822 ( .DIN1(n3734), .DIN2(n3735), .DIN3(n3736), .Q(n3730) );
  nnd2s1 U3823 ( .DIN1(n3266), .DIN2(n3685), .Q(n3736) );
  nnd2s1 U3824 ( .DIN1(n3406), .DIN2(n3379), .Q(n3685) );
  nnd2s1 U3825 ( .DIN1(n3263), .DIN2(n3737), .Q(n3735) );
  nnd2s1 U3826 ( .DIN1(n3528), .DIN2(n3357), .Q(n3737) );
  nor2s1 U3827 ( .DIN1(n3419), .DIN2(n3397), .Q(n3528) );
  nnd2s1 U3828 ( .DIN1(n3556), .DIN2(n3738), .Q(n3734) );
  nnd2s1 U3829 ( .DIN1(n3440), .DIN2(n3281), .Q(n3738) );
  nnd2s1 U3830 ( .DIN1(n3419), .DIN2(n3739), .Q(n3729) );
  nnd2s1 U3831 ( .DIN1(n3465), .DIN2(n3274), .Q(n3739) );
  nnd2s1 U3832 ( .DIN1(n3342), .DIN2(n3740), .Q(n3728) );
  nnd3s1 U3833 ( .DIN1(n3278), .DIN2(n3317), .DIN3(n3313), .Q(n3740) );
  nor4s1 U3834 ( .DIN1(n3741), .DIN2(n3742), .DIN3(n3743), .DIN4(n3744), 
        .Q(n3625) );
  nnd4s1 U3835 ( .DIN1(n3745), .DIN2(n3746), .DIN3(n3747), .DIN4(n3748), 
        .Q(n3744) );
  and3s1 U3836 ( .DIN1(n3749), .DIN2(n3750), .DIN3(n3751), .Q(n3748) );
  nnd2s1 U3837 ( .DIN1(n3261), .DIN2(n3409), .Q(n3751) );
  nnd2s1 U3838 ( .DIN1(n3262), .DIN2(n3752), .Q(n3750) );
  nnd2s1 U3839 ( .DIN1(n3355), .DIN2(n3753), .Q(n3752) );
  nnd2s1 U3840 ( .DIN1(n3275), .DIN2(n3651), .Q(n3749) );
  nnd2s1 U3841 ( .DIN1(n3348), .DIN2(n3351), .Q(n3651) );
  nnd2s1 U3842 ( .DIN1(n3254), .DIN2(n3754), .Q(n3747) );
  nnd2s1 U3843 ( .DIN1(n3316), .DIN2(n3375), .Q(n3754) );
  nnd2s1 U3844 ( .DIN1(n3264), .DIN2(n3755), .Q(n3746) );
  nnd2s1 U3845 ( .DIN1(n3274), .DIN2(n3282), .Q(n3755) );
  nnd2s1 U3846 ( .DIN1(n3556), .DIN2(n3756), .Q(n3745) );
  nnd2s1 U3847 ( .DIN1(n3483), .DIN2(n3484), .Q(n3756) );
  nnd3s1 U3848 ( .DIN1(n3757), .DIN2(n3758), .DIN3(n3759), .Q(n3743) );
  nnd2s1 U3849 ( .DIN1(n3376), .DIN2(n3340), .Q(n3759) );
  nnd2s1 U3850 ( .DIN1(n3369), .DIN2(n3298), .Q(n3758) );
  nnd2s1 U3851 ( .DIN1(n3266), .DIN2(n3283), .Q(n3757) );
  nor2s1 U3852 ( .DIN1(n3437), .DIN2(n3547), .Q(n3742) );
  nor2s1 U3853 ( .DIN1(n3348), .DIN2(n3465), .Q(n3741) );
  nor4s1 U3854 ( .DIN1(n3760), .DIN2(n3761), .DIN3(n3762), .DIN4(n3763), 
        .Q(n3247) );
  nnd4s1 U3855 ( .DIN1(n3764), .DIN2(n3765), .DIN3(n3766), .DIN4(n3767), 
        .Q(n3763) );
  nnd2s1 U3856 ( .DIN1(n3369), .DIN2(n3262), .Q(n3767) );
  nnd2s1 U3857 ( .DIN1(n3255), .DIN2(n3264), .Q(n3766) );
  nnd2s1 U3858 ( .DIN1(n3298), .DIN2(n3283), .Q(n3765) );
  hi1s1 U3859 ( .DIN(n3375), .Q(n3298) );
  nnd2s1 U3860 ( .DIN1(n3253), .DIN2(n3263), .Q(n3764) );
  nnd3s1 U3861 ( .DIN1(n3768), .DIN2(n3769), .DIN3(n3770), .Q(n3762) );
  nnd2s1 U3862 ( .DIN1(n3341), .DIN2(n3771), .Q(n3770) );
  nnd3s1 U3863 ( .DIN1(n3753), .DIN2(n3379), .DIN3(n3437), .Q(n3771) );
  nnd2s1 U3864 ( .DIN1(n3266), .DIN2(n3772), .Q(n3769) );
  nnd2s1 U3865 ( .DIN1(n3436), .DIN2(n3521), .Q(n3772) );
  hi1s1 U3866 ( .DIN(n3303), .Q(n3266) );
  nnd2s1 U3867 ( .DIN1(n3366), .DIN2(n3773), .Q(n3768) );
  nnd2s1 U3868 ( .DIN1(n3277), .DIN2(n3507), .Q(n3773) );
  nor2s1 U3869 ( .DIN1(n3357), .DIN2(n3282), .Q(n3761) );
  and2s1 U3870 ( .DIN1(n3420), .DIN2(n3774), .Q(n3760) );
  nnd4s1 U3871 ( .DIN1(n3375), .DIN2(n3316), .DIN3(n3313), .DIN4(n3317), 
        .Q(n3774) );
  nnd3s1 U3872 ( .DIN1(n3775), .DIN2(n3776), .DIN3(n3777), .Q(n3722) );
  nnd2s1 U3873 ( .DIN1(n3310), .DIN2(n3262), .Q(n3777) );
  nnd2s1 U3874 ( .DIN1(n3556), .DIN2(n3261), .Q(n3776) );
  nnd2s1 U3875 ( .DIN1(n3339), .DIN2(n3299), .Q(n3775) );
  nnd4s1 U3876 ( .DIN1(n3778), .DIN2(n3779), .DIN3(n3780), .DIN4(n3781), 
        .Q(n3721) );
  nnd2s1 U3877 ( .DIN1(n3409), .DIN2(n3782), .Q(n3781) );
  nnd2s1 U3878 ( .DIN1(n3444), .DIN2(n3281), .Q(n3782) );
  nnd2s1 U3879 ( .DIN1(n3419), .DIN2(n3783), .Q(n3780) );
  nnd4s1 U3880 ( .DIN1(n3521), .DIN2(n3484), .DIN3(n3437), .DIN4(n3444), 
        .Q(n3783) );
  nnd2s1 U3881 ( .DIN1(n3376), .DIN2(n3525), .Q(n3779) );
  nnd2s1 U3882 ( .DIN1(n3491), .DIN2(n3278), .Q(n3525) );
  nnd2s1 U3883 ( .DIN1(n3263), .DIN2(n3429), .Q(n3778) );
  nnd2s1 U3884 ( .DIN1(n3303), .DIN2(n3312), .Q(n3429) );
  nor4s1 U3885 ( .DIN1(n3784), .DIN2(n3785), .DIN3(n3786), .DIN4(n3787), 
        .Q(n3248) );
  nnd4s1 U3886 ( .DIN1(n3788), .DIN2(n3789), .DIN3(n3790), .DIN4(n3791), 
        .Q(n3787) );
  nnd2s1 U3887 ( .DIN1(n3279), .DIN2(n3263), .Q(n3791) );
  nor2s1 U3888 ( .DIN1(n3792), .DIN2(n3520), .Q(n3790) );
  nor2s1 U3889 ( .DIN1(n3351), .DIN2(n3281), .Q(n3520) );
  nor2s1 U3890 ( .DIN1(n3337), .DIN2(n3379), .Q(n3792) );
  nnd2s1 U3891 ( .DIN1(n3262), .DIN2(n3366), .Q(n3789) );
  hi1s1 U3892 ( .DIN(n3278), .Q(n3262) );
  nnd2s1 U3893 ( .DIN1(n3349), .DIN2(n3352), .Q(n3788) );
  nnd3s1 U3894 ( .DIN1(n3793), .DIN2(n3794), .DIN3(n3795), .Q(n3786) );
  nnd2s1 U3895 ( .DIN1(n3342), .DIN2(n3427), .Q(n3795) );
  nnd2s1 U3896 ( .DIN1(n3348), .DIN2(n3337), .Q(n3427) );
  nnd2s1 U3897 ( .DIN1(n3264), .DIN2(n3796), .Q(n3794) );
  nnd3s1 U3898 ( .DIN1(n3437), .DIN2(n3444), .DIN3(n3484), .Q(n3796) );
  nnd2s1 U3899 ( .DIN1(n3340), .DIN2(n3797), .Q(n3793) );
  nnd3s1 U3900 ( .DIN1(n3753), .DIN2(n3439), .DIN3(n3483), .Q(n3797) );
  nor2s1 U3901 ( .DIN1(n3753), .DIN2(n3357), .Q(n3785) );
  nnd2s1 U3902 ( .DIN1(n3798), .DIN2(n3799), .Q(n3357) );
  nor2s1 U3903 ( .DIN1(n3592), .DIN2(n3507), .Q(n3784) );
  nor2s1 U3904 ( .DIN1(n3310), .DIN2(n3283), .Q(n3592) );
  nor4s1 U3905 ( .DIN1(n3800), .DIN2(n3801), .DIN3(n3802), .DIN4(n3803), 
        .Q(n3618) );
  nnd4s1 U3906 ( .DIN1(n3804), .DIN2(n3805), .DIN3(n3806), .DIN4(n3807), 
        .Q(n3803) );
  nnd2s1 U3907 ( .DIN1(n3349), .DIN2(n3397), .Q(n3807) );
  nor2s1 U3908 ( .DIN1(n3808), .DIN2(n3809), .Q(n3806) );
  nor2s1 U3909 ( .DIN1(n3282), .DIN2(n3348), .Q(n3809) );
  nor2s1 U3910 ( .DIN1(n3402), .DIN2(n3521), .Q(n3808) );
  nor2s1 U3911 ( .DIN1(n3279), .DIN2(n3397), .Q(n3402) );
  hi1s1 U3912 ( .DIN(n3351), .Q(n3397) );
  nnd2s1 U3913 ( .DIN1(n3256), .DIN2(n3263), .Q(n3805) );
  hi1s1 U3914 ( .DIN(n3317), .Q(n3256) );
  nnd2s1 U3915 ( .DIN1(n3556), .DIN2(n3342), .Q(n3804) );
  nnd3s1 U3916 ( .DIN1(n3810), .DIN2(n3811), .DIN3(n3812), .Q(n3802) );
  nnd2s1 U3917 ( .DIN1(n3254), .DIN2(n3463), .Q(n3812) );
  nnd2s1 U3918 ( .DIN1(n3312), .DIN2(n3408), .Q(n3463) );
  nnd2s1 U3919 ( .DIN1(n3299), .DIN2(n3813), .Q(n3811) );
  nnd2s1 U3920 ( .DIN1(n3483), .DIN2(n3355), .Q(n3813) );
  nnd2s1 U3921 ( .DIN1(n3340), .DIN2(n3814), .Q(n3810) );
  nnd2s1 U3922 ( .DIN1(n3274), .DIN2(n3521), .Q(n3814) );
  hi1s1 U3923 ( .DIN(n3313), .Q(n3340) );
  nor2s1 U3924 ( .DIN1(n3815), .DIN2(n3278), .Q(n3801) );
  nor2s1 U3925 ( .DIN1(n3255), .DIN2(n3339), .Q(n3815) );
  nor2s1 U3926 ( .DIN1(n3816), .DIN2(n3303), .Q(n3800) );
  nnd2s1 U3927 ( .DIN1(n3798), .DIN2(n3817), .Q(n3303) );
  nor2s1 U3928 ( .DIN1(n3261), .DIN2(n3310), .Q(n3816) );
  hi1s1 U3929 ( .DIN(n3465), .Q(n3310) );
  nnd3s1 U3930 ( .DIN1(w3[2]), .DIN2(n1556), .DIN3(n3818), .Q(n3465) );
  hi1s1 U3931 ( .DIN(n3282), .Q(n3261) );
  nnd4s1 U3932 ( .DIN1(n3627), .DIN2(n3819), .DIN3(n3820), .DIN4(n3821), 
        .Q(n3719) );
  nnd2s1 U3933 ( .DIN1(n3253), .DIN2(n3349), .Q(n3821) );
  hi1s1 U3934 ( .DIN(n3436), .Q(n3349) );
  hi1s1 U3935 ( .DIN(n3348), .Q(n3253) );
  nnd2s1 U3936 ( .DIN1(n3339), .DIN2(n3279), .Q(n3820) );
  nnd2s1 U3937 ( .DIN1(n3419), .DIN2(n3366), .Q(n3819) );
  hi1s1 U3938 ( .DIN(n3316), .Q(n3419) );
  and4s1 U3939 ( .DIN1(n3822), .DIN2(n3823), .DIN3(n3824), .DIN4(n3825), 
        .Q(n3627) );
  and4s1 U3940 ( .DIN1(n3826), .DIN2(n3536), .DIN3(n3827), .DIN4(n3828), 
        .Q(n3825) );
  nnd2s1 U3941 ( .DIN1(n3369), .DIN2(n3409), .Q(n3828) );
  nnd2s1 U3942 ( .DIN1(n3263), .DIN2(n3299), .Q(n3827) );
  hi1s1 U3943 ( .DIN(n3337), .Q(n3299) );
  hi1s1 U3944 ( .DIN(n3439), .Q(n3263) );
  nnd3s1 U3945 ( .DIN1(n1556), .DIN2(n1369), .DIN3(n3818), .Q(n3439) );
  nnd2s1 U3946 ( .DIN1(n3275), .DIN2(n3556), .Q(n3536) );
  hi1s1 U3947 ( .DIN(n3312), .Q(n3556) );
  nnd2s1 U3948 ( .DIN1(n3255), .DIN2(n3279), .Q(n3826) );
  hi1s1 U3949 ( .DIN(n3547), .Q(n3279) );
  nnd2s1 U3950 ( .DIN1(n3798), .DIN2(n3829), .Q(n3547) );
  and3s1 U3951 ( .DIN1(n3830), .DIN2(n3831), .DIN3(n3832), .Q(n3824) );
  nnd2s1 U3952 ( .DIN1(n3366), .DIN2(n3833), .Q(n3832) );
  nnd2s1 U3953 ( .DIN1(n3317), .DIN2(n3348), .Q(n3833) );
  hi1s1 U3954 ( .DIN(n3483), .Q(n3366) );
  nnd3s1 U3955 ( .DIN1(n3834), .DIN2(n1411), .DIN3(w3[0]), .Q(n3483) );
  nnd2s1 U3956 ( .DIN1(n3254), .DIN2(n3835), .Q(n3831) );
  nnd2s1 U3957 ( .DIN1(n3277), .DIN2(n3317), .Q(n3835) );
  nnd2s1 U3958 ( .DIN1(n3799), .DIN2(n3836), .Q(n3317) );
  hi1s1 U3959 ( .DIN(n3379), .Q(n3254) );
  nnd3s1 U3960 ( .DIN1(w3[0]), .DIN2(n1411), .DIN3(n3837), .Q(n3379) );
  nnd2s1 U3961 ( .DIN1(n3339), .DIN2(n3584), .Q(n3830) );
  nnd2s1 U3962 ( .DIN1(n3351), .DIN2(n3375), .Q(n3584) );
  hi1s1 U3963 ( .DIN(n3484), .Q(n3339) );
  nnd3s1 U3964 ( .DIN1(w3[0]), .DIN2(n3838), .DIN3(w3[2]), .Q(n3484) );
  nnd2s1 U3965 ( .DIN1(n3314), .DIN2(n3839), .Q(n3823) );
  nnd3s1 U3966 ( .DIN1(n3316), .DIN2(n3278), .DIN3(n3375), .Q(n3839) );
  nnd2s1 U3967 ( .DIN1(n3817), .DIN2(n3836), .Q(n3278) );
  nnd2s1 U3968 ( .DIN1(n3829), .DIN2(n3840), .Q(n3316) );
  hi1s1 U3969 ( .DIN(n3281), .Q(n3314) );
  nnd3s1 U3970 ( .DIN1(w3[2]), .DIN2(w3[0]), .DIN3(n3818), .Q(n3281) );
  or2s1 U3971 ( .DIN1(n3348), .DIN2(n3674), .Q(n3822) );
  nor2s1 U3972 ( .DIN1(n3265), .DIN2(n3283), .Q(n3674) );
  hi1s1 U3973 ( .DIN(n3753), .Q(n3283) );
  nnd3s1 U3974 ( .DIN1(n3838), .DIN2(n1369), .DIN3(w3[0]), .Q(n3753) );
  hi1s1 U3975 ( .DIN(n3274), .Q(n3265) );
  nnd3s1 U3976 ( .DIN1(n3834), .DIN2(n1556), .DIN3(w3[1]), .Q(n3274) );
  nnd4s1 U3977 ( .DIN1(n3452), .DIN2(n3841), .DIN3(n3842), .DIN4(n3843), 
        .Q(n3718) );
  nnd2s1 U3978 ( .DIN1(n3352), .DIN2(n3602), .Q(n3843) );
  nnd2s1 U3979 ( .DIN1(n3440), .DIN2(n3282), .Q(n3602) );
  nnd3s1 U3980 ( .DIN1(w3[1]), .DIN2(w3[0]), .DIN3(n3837), .Q(n3282) );
  hi1s1 U3981 ( .DIN(n3277), .Q(n3352) );
  nnd2s1 U3982 ( .DIN1(n3840), .DIN2(n3844), .Q(n3277) );
  nnd2s1 U3983 ( .DIN1(n3376), .DIN2(n3284), .Q(n3842) );
  nnd2s1 U3984 ( .DIN1(n3351), .DIN2(n3408), .Q(n3284) );
  nnd2s1 U3985 ( .DIN1(n3798), .DIN2(n3844), .Q(n3351) );
  nor2s1 U3986 ( .DIN1(n1441), .DIN2(w3[6]), .Q(n3798) );
  hi1s1 U3987 ( .DIN(n3440), .Q(n3376) );
  nnd3s1 U3988 ( .DIN1(n3838), .DIN2(n1556), .DIN3(w3[2]), .Q(n3440) );
  nnd2s1 U3989 ( .DIN1(n3409), .DIN2(n3342), .Q(n3841) );
  hi1s1 U3990 ( .DIN(n3507), .Q(n3409) );
  nnd2s1 U3991 ( .DIN1(n3829), .DIN2(n3845), .Q(n3507) );
  nnd2s1 U3992 ( .DIN1(n3369), .DIN2(n3264), .Q(n3452) );
  hi1s1 U3993 ( .DIN(n3408), .Q(n3264) );
  nnd2s1 U3994 ( .DIN1(n3836), .DIN2(n3844), .Q(n3408) );
  hi1s1 U3995 ( .DIN(n3521), .Q(n3369) );
  nnd3s1 U3996 ( .DIN1(w3[0]), .DIN2(n1369), .DIN3(n3818), .Q(n3521) );
  nor2s1 U3997 ( .DIN1(n1411), .DIN2(w3[3]), .Q(n3818) );
  nnd4s1 U3998 ( .DIN1(n3846), .DIN2(n3847), .DIN3(n3848), .DIN4(n3849), 
        .Q(n3717) );
  nnd2s1 U3999 ( .DIN1(n3255), .DIN2(n3850), .Q(n3849) );
  nnd2s1 U4000 ( .DIN1(n3313), .DIN2(n3337), .Q(n3850) );
  nnd2s1 U4001 ( .DIN1(n3799), .DIN2(n3845), .Q(n3337) );
  nnd2s1 U4002 ( .DIN1(n3845), .DIN2(n3844), .Q(n3313) );
  nor2s1 U4003 ( .DIN1(n1442), .DIN2(n1375), .Q(n3844) );
  hi1s1 U4004 ( .DIN(n3406), .Q(n3255) );
  nnd3s1 U4005 ( .DIN1(n1556), .DIN2(n1411), .DIN3(n3834), .Q(n3406) );
  nnd2s1 U4006 ( .DIN1(n3341), .DIN2(n3851), .Q(n3848) );
  nnd2s1 U4007 ( .DIN1(n3444), .DIN2(n3436), .Q(n3851) );
  nnd3s1 U4008 ( .DIN1(n1556), .DIN2(n1411), .DIN3(n3837), .Q(n3436) );
  hi1s1 U4009 ( .DIN(n3491), .Q(n3341) );
  nnd2s1 U4010 ( .DIN1(n3829), .DIN2(n3836), .Q(n3491) );
  nor2s1 U4011 ( .DIN1(n1391), .DIN2(w3[4]), .Q(n3836) );
  nor2s1 U4012 ( .DIN1(w3[7]), .DIN2(w3[5]), .Q(n3829) );
  or2s1 U4013 ( .DIN1(n3375), .DIN2(n3354), .Q(n3847) );
  nor2s1 U4014 ( .DIN1(n3275), .DIN2(n3342), .Q(n3354) );
  hi1s1 U4015 ( .DIN(n3437), .Q(n3342) );
  nnd3s1 U4016 ( .DIN1(w3[0]), .DIN2(n3834), .DIN3(w3[1]), .Q(n3437) );
  nor2s1 U4017 ( .DIN1(n1440), .DIN2(w3[2]), .Q(n3834) );
  hi1s1 U4018 ( .DIN(n3444), .Q(n3275) );
  nnd3s1 U4019 ( .DIN1(n1556), .DIN2(n1369), .DIN3(n3838), .Q(n3444) );
  nor2s1 U4020 ( .DIN1(w3[3]), .DIN2(w3[1]), .Q(n3838) );
  nnd2s1 U4021 ( .DIN1(n3817), .DIN2(n3845), .Q(n3375) );
  nor2s1 U4022 ( .DIN1(n1441), .DIN2(n1391), .Q(n3845) );
  nnd2s1 U4023 ( .DIN1(n3420), .DIN2(n3367), .Q(n3846) );
  nnd2s1 U4024 ( .DIN1(n3348), .DIN2(n3312), .Q(n3367) );
  nnd2s1 U4025 ( .DIN1(n3840), .DIN2(n3799), .Q(n3312) );
  nor2s1 U4026 ( .DIN1(n1442), .DIN2(w3[5]), .Q(n3799) );
  nnd2s1 U4027 ( .DIN1(n3817), .DIN2(n3840), .Q(n3348) );
  nor2s1 U4028 ( .DIN1(w3[6]), .DIN2(w3[4]), .Q(n3840) );
  nor2s1 U4029 ( .DIN1(n1375), .DIN2(w3[7]), .Q(n3817) );
  hi1s1 U4030 ( .DIN(n3355), .Q(n3420) );
  nnd3s1 U4031 ( .DIN1(w3[1]), .DIN2(n1556), .DIN3(n3837), .Q(n3355) );
  nor2s1 U4032 ( .DIN1(n1369), .DIN2(n1440), .Q(n3837) );
  nnd2s1 U4033 ( .DIN1(n3852), .DIN2(n3853), .Q(\u0/N115 ) );
  nnd2s1 U4034 ( .DIN1(\key[71] ), .DIN2(ld), .Q(n3853) );
  nnd2s1 U4035 ( .DIN1(n1982), .DIN2(n1568), .Q(n3852) );
  xnr2s1 U4036 ( .DIN1(w1[7]), .DIN2(n1758), .Q(n1982) );
  xor2s1 U4037 ( .DIN1(w0[7]), .DIN2(n3854), .Q(n1758) );
  nor4s1 U4038 ( .DIN1(n3855), .DIN2(n3856), .DIN3(n3857), .DIN4(n3858), 
        .Q(n3854) );
  nnd3s1 U4039 ( .DIN1(n3859), .DIN2(n3860), .DIN3(n3861), .Q(n3858) );
  nnd4s1 U4040 ( .DIN1(n3862), .DIN2(n3863), .DIN3(n3864), .DIN4(n3865), 
        .Q(n3857) );
  nnd2s1 U4041 ( .DIN1(n3866), .DIN2(n3867), .Q(n3864) );
  nnd2s1 U4042 ( .DIN1(n3868), .DIN2(n3869), .Q(n3863) );
  nnd4s1 U4043 ( .DIN1(n3870), .DIN2(n3871), .DIN3(n3872), .DIN4(n3873), 
        .Q(n3856) );
  nnd2s1 U4044 ( .DIN1(n3874), .DIN2(n3875), .Q(n3873) );
  nnd2s1 U4045 ( .DIN1(n3876), .DIN2(n3877), .Q(n3872) );
  nnd2s1 U4046 ( .DIN1(n3878), .DIN2(n3879), .Q(n3871) );
  nnd4s1 U4047 ( .DIN1(n3880), .DIN2(n3881), .DIN3(n3882), .DIN4(n3883), 
        .Q(n3855) );
  nnd2s1 U4048 ( .DIN1(n3884), .DIN2(n3885), .Q(n3883) );
  nnd2s1 U4049 ( .DIN1(n3886), .DIN2(n3887), .Q(n3885) );
  nnd2s1 U4050 ( .DIN1(n3888), .DIN2(n3889), .Q(n3882) );
  nnd2s1 U4051 ( .DIN1(n3890), .DIN2(n3891), .Q(n3889) );
  nnd2s1 U4052 ( .DIN1(n3892), .DIN2(n3893), .Q(n3881) );
  nnd2s1 U4053 ( .DIN1(n3894), .DIN2(n3895), .Q(n3893) );
  nnd2s1 U4054 ( .DIN1(n3896), .DIN2(n3897), .Q(n3880) );
  nnd2s1 U4055 ( .DIN1(n3898), .DIN2(n3899), .Q(\u0/N114 ) );
  nnd2s1 U4056 ( .DIN1(\key[70] ), .DIN2(ld), .Q(n3899) );
  nnd2s1 U4057 ( .DIN1(n1985), .DIN2(n1569), .Q(n3898) );
  xnr2s1 U4058 ( .DIN1(w1[6]), .DIN2(n1761), .Q(n1985) );
  xnr2s1 U4059 ( .DIN1(n1504), .DIN2(n3900), .Q(n1761) );
  nor4s1 U4060 ( .DIN1(n3901), .DIN2(n3902), .DIN3(n3903), .DIN4(n3904), 
        .Q(n3900) );
  nnd3s1 U4061 ( .DIN1(n3905), .DIN2(n3906), .DIN3(n3907), .Q(n3904) );
  nnd3s1 U4062 ( .DIN1(n3908), .DIN2(n3909), .DIN3(n3910), .Q(n3903) );
  nnd2s1 U4063 ( .DIN1(n3911), .DIN2(n3876), .Q(n3909) );
  nnd2s1 U4064 ( .DIN1(n3867), .DIN2(n3912), .Q(n3908) );
  nnd3s1 U4065 ( .DIN1(n3913), .DIN2(n3914), .DIN3(n3915), .Q(n3902) );
  or2s1 U4066 ( .DIN1(n3916), .DIN2(n3917), .Q(n3915) );
  or2s1 U4067 ( .DIN1(n3891), .DIN2(n3918), .Q(n3914) );
  nnd2s1 U4068 ( .DIN1(n3892), .DIN2(n3919), .Q(n3913) );
  nnd3s1 U4069 ( .DIN1(n3920), .DIN2(n3921), .DIN3(n3922), .Q(n3901) );
  nnd2s1 U4070 ( .DIN1(n3923), .DIN2(n3924), .Q(n3922) );
  nnd2s1 U4071 ( .DIN1(n3925), .DIN2(n3926), .Q(n3924) );
  nnd2s1 U4072 ( .DIN1(n3927), .DIN2(n3928), .Q(n3921) );
  nnd2s1 U4073 ( .DIN1(n3929), .DIN2(n3930), .Q(n3928) );
  nnd2s1 U4074 ( .DIN1(n3868), .DIN2(n3931), .Q(n3920) );
  nnd2s1 U4075 ( .DIN1(n3932), .DIN2(n3933), .Q(n3931) );
  hi1s1 U4076 ( .DIN(n3934), .Q(n3933) );
  nnd2s1 U4077 ( .DIN1(n3935), .DIN2(n3936), .Q(\u0/N113 ) );
  nnd2s1 U4078 ( .DIN1(\key[69] ), .DIN2(ld), .Q(n3936) );
  nnd2s1 U4079 ( .DIN1(n1988), .DIN2(n1569), .Q(n3935) );
  xnr2s1 U4080 ( .DIN1(w1[5]), .DIN2(n1764), .Q(n1988) );
  xnr2s1 U4081 ( .DIN1(n1471), .DIN2(n3937), .Q(n1764) );
  nor4s1 U4082 ( .DIN1(n3938), .DIN2(n3939), .DIN3(n3940), .DIN4(n3941), 
        .Q(n3937) );
  nnd3s1 U4083 ( .DIN1(n3942), .DIN2(n3906), .DIN3(n3943), .Q(n3941) );
  nor2s1 U4084 ( .DIN1(n3944), .DIN2(n3945), .Q(n3906) );
  nnd4s1 U4085 ( .DIN1(n3946), .DIN2(n3947), .DIN3(n3948), .DIN4(n3949), 
        .Q(n3945) );
  or2s1 U4086 ( .DIN1(n3950), .DIN2(n3951), .Q(n3949) );
  nnd2s1 U4087 ( .DIN1(n3952), .DIN2(n3953), .Q(n3948) );
  nnd2s1 U4088 ( .DIN1(n3954), .DIN2(n3867), .Q(n3947) );
  nnd2s1 U4089 ( .DIN1(n3879), .DIN2(n3955), .Q(n3946) );
  nnd4s1 U4090 ( .DIN1(n3956), .DIN2(n3957), .DIN3(n3958), .DIN4(n3959), 
        .Q(n3944) );
  nnd2s1 U4091 ( .DIN1(n3878), .DIN2(n3960), .Q(n3959) );
  nnd2s1 U4092 ( .DIN1(n3929), .DIN2(n3961), .Q(n3960) );
  nnd2s1 U4093 ( .DIN1(n3962), .DIN2(n3963), .Q(n3958) );
  nnd2s1 U4094 ( .DIN1(n3925), .DIN2(n3964), .Q(n3963) );
  nnd2s1 U4095 ( .DIN1(n3965), .DIN2(n3966), .Q(n3957) );
  nnd2s1 U4096 ( .DIN1(n3967), .DIN2(n3968), .Q(n3966) );
  nnd2s1 U4097 ( .DIN1(n3888), .DIN2(n3969), .Q(n3956) );
  nnd3s1 U4098 ( .DIN1(n3929), .DIN2(n3970), .DIN3(n3971), .Q(n3969) );
  nnd4s1 U4099 ( .DIN1(n3972), .DIN2(n3973), .DIN3(n3974), .DIN4(n3865), 
        .Q(n3940) );
  nnd2s1 U4100 ( .DIN1(n3954), .DIN2(n3927), .Q(n3865) );
  nnd2s1 U4101 ( .DIN1(n3923), .DIN2(n3965), .Q(n3974) );
  nnd2s1 U4102 ( .DIN1(n3952), .DIN2(n3869), .Q(n3973) );
  nnd4s1 U4103 ( .DIN1(n3975), .DIN2(n3976), .DIN3(n3977), .DIN4(n3978), 
        .Q(n3939) );
  nnd2s1 U4104 ( .DIN1(n3979), .DIN2(n3980), .Q(n3978) );
  nnd2s1 U4105 ( .DIN1(n3879), .DIN2(n3981), .Q(n3977) );
  nnd2s1 U4106 ( .DIN1(n3866), .DIN2(n3982), .Q(n3976) );
  nnd2s1 U4107 ( .DIN1(n3911), .DIN2(n3955), .Q(n3975) );
  nnd4s1 U4108 ( .DIN1(n3983), .DIN2(n3984), .DIN3(n3985), .DIN4(n3986), 
        .Q(n3938) );
  nnd2s1 U4109 ( .DIN1(n3896), .DIN2(n3987), .Q(n3986) );
  nnd2s1 U4110 ( .DIN1(n3926), .DIN2(n3988), .Q(n3987) );
  nnd2s1 U4111 ( .DIN1(n3989), .DIN2(n3990), .Q(n3985) );
  nnd2s1 U4112 ( .DIN1(n3892), .DIN2(n3991), .Q(n3984) );
  nnd2s1 U4113 ( .DIN1(n3992), .DIN2(n3887), .Q(n3991) );
  nnd2s1 U4114 ( .DIN1(n3876), .DIN2(n3993), .Q(n3983) );
  nnd2s1 U4115 ( .DIN1(n3994), .DIN2(n3995), .Q(\u0/N112 ) );
  nnd2s1 U4116 ( .DIN1(\key[68] ), .DIN2(ld), .Q(n3995) );
  nnd2s1 U4117 ( .DIN1(n1991), .DIN2(n1569), .Q(n3994) );
  xnr2s1 U4118 ( .DIN1(w1[4]), .DIN2(n1767), .Q(n1991) );
  xnr2s1 U4119 ( .DIN1(n1472), .DIN2(n3996), .Q(n1767) );
  nor4s1 U4120 ( .DIN1(n3997), .DIN2(n3998), .DIN3(n3999), .DIN4(n4000), 
        .Q(n3996) );
  nnd3s1 U4121 ( .DIN1(n3942), .DIN2(n3907), .DIN3(n4001), .Q(n4000) );
  and4s1 U4122 ( .DIN1(n4002), .DIN2(n4003), .DIN3(n4004), .DIN4(n4005), 
        .Q(n3907) );
  and4s1 U4123 ( .DIN1(n4006), .DIN2(n4007), .DIN3(n4008), .DIN4(n4009), 
        .Q(n4005) );
  nnd2s1 U4124 ( .DIN1(n3874), .DIN2(n3911), .Q(n4009) );
  nnd2s1 U4125 ( .DIN1(n3952), .DIN2(n4010), .Q(n4007) );
  nnd2s1 U4126 ( .DIN1(n3962), .DIN2(n3875), .Q(n4006) );
  and3s1 U4127 ( .DIN1(n4011), .DIN2(n4012), .DIN3(n4013), .Q(n4004) );
  nnd2s1 U4128 ( .DIN1(n3979), .DIN2(n4014), .Q(n4013) );
  nnd2s1 U4129 ( .DIN1(n4015), .DIN2(n3890), .Q(n4014) );
  nnd2s1 U4130 ( .DIN1(n3888), .DIN2(n4016), .Q(n4012) );
  nnd2s1 U4131 ( .DIN1(n4017), .DIN2(n3988), .Q(n4016) );
  nnd2s1 U4132 ( .DIN1(n3954), .DIN2(n4018), .Q(n4011) );
  nnd2s1 U4133 ( .DIN1(n4019), .DIN2(n3887), .Q(n4018) );
  nnd2s1 U4134 ( .DIN1(n3867), .DIN2(n4020), .Q(n4003) );
  nnd3s1 U4135 ( .DIN1(n4021), .DIN2(n3926), .DIN3(n3929), .Q(n4020) );
  nnd2s1 U4136 ( .DIN1(n3896), .DIN2(n4022), .Q(n4002) );
  nor3s1 U4137 ( .DIN1(n4023), .DIN2(n4024), .DIN3(n4025), .Q(n3942) );
  nnd4s1 U4138 ( .DIN1(n3905), .DIN2(n4026), .DIN3(n4027), .DIN4(n4028), 
        .Q(n4025) );
  and3s1 U4139 ( .DIN1(n4029), .DIN2(n4030), .DIN3(n4031), .Q(n4028) );
  nnd2s1 U4140 ( .DIN1(n3954), .DIN2(n3955), .Q(n4031) );
  nnd2s1 U4141 ( .DIN1(n4032), .DIN2(n3868), .Q(n4030) );
  nnd2s1 U4142 ( .DIN1(n4033), .DIN2(n3879), .Q(n4029) );
  nor2s1 U4143 ( .DIN1(n4034), .DIN2(n4035), .Q(n3905) );
  nnd4s1 U4144 ( .DIN1(n4036), .DIN2(n4037), .DIN3(n4038), .DIN4(n4039), 
        .Q(n4035) );
  nnd2s1 U4145 ( .DIN1(n3923), .DIN2(n4040), .Q(n4039) );
  nnd2s1 U4146 ( .DIN1(n3892), .DIN2(n4041), .Q(n4038) );
  nnd2s1 U4147 ( .DIN1(n3874), .DIN2(n4042), .Q(n4037) );
  nnd2s1 U4148 ( .DIN1(n3888), .DIN2(n3912), .Q(n4036) );
  nnd4s1 U4149 ( .DIN1(n4043), .DIN2(n4044), .DIN3(n4045), .DIN4(n4046), 
        .Q(n4034) );
  nnd2s1 U4150 ( .DIN1(n3911), .DIN2(n4041), .Q(n4046) );
  nnd2s1 U4151 ( .DIN1(n3878), .DIN2(n4047), .Q(n4045) );
  nnd2s1 U4152 ( .DIN1(n3930), .DIN2(n3964), .Q(n4047) );
  nnd2s1 U4153 ( .DIN1(n3866), .DIN2(n4048), .Q(n4044) );
  nnd2s1 U4154 ( .DIN1(n4049), .DIN2(n4050), .Q(n4048) );
  nnd2s1 U4155 ( .DIN1(n4032), .DIN2(n4051), .Q(n4043) );
  nnd3s1 U4156 ( .DIN1(n3895), .DIN2(n4052), .DIN3(n4053), .Q(n4051) );
  nnd3s1 U4157 ( .DIN1(n4054), .DIN2(n4055), .DIN3(n3870), .Q(n4024) );
  nnd2s1 U4158 ( .DIN1(n3962), .DIN2(n3953), .Q(n3870) );
  nnd2s1 U4159 ( .DIN1(n3866), .DIN2(n4056), .Q(n4055) );
  nnd3s1 U4160 ( .DIN1(n3968), .DIN2(n4057), .DIN3(n3918), .Q(n4056) );
  nor2s1 U4161 ( .DIN1(n3989), .DIN2(n3868), .Q(n3918) );
  nnd2s1 U4162 ( .DIN1(n3965), .DIN2(n3896), .Q(n4054) );
  nnd3s1 U4163 ( .DIN1(n4058), .DIN2(n4059), .DIN3(n4060), .Q(n4023) );
  nnd2s1 U4164 ( .DIN1(n3979), .DIN2(n4061), .Q(n4060) );
  nnd2s1 U4165 ( .DIN1(n3950), .DIN2(n3988), .Q(n4061) );
  nnd2s1 U4166 ( .DIN1(n3876), .DIN2(n4062), .Q(n4059) );
  nnd2s1 U4167 ( .DIN1(n3964), .DIN2(n3950), .Q(n4062) );
  nnd2s1 U4168 ( .DIN1(n3923), .DIN2(n4063), .Q(n4058) );
  nnd2s1 U4169 ( .DIN1(n4017), .DIN2(n3930), .Q(n4063) );
  nnd3s1 U4170 ( .DIN1(n4064), .DIN2(n4065), .DIN3(n4066), .Q(n3999) );
  nnd3s1 U4171 ( .DIN1(n4067), .DIN2(n4068), .DIN3(n4069), .Q(n3998) );
  nnd2s1 U4172 ( .DIN1(n3952), .DIN2(n4042), .Q(n4069) );
  nnd2s1 U4173 ( .DIN1(n3876), .DIN2(n3980), .Q(n4068) );
  nnd2s1 U4174 ( .DIN1(n3965), .DIN2(n3981), .Q(n4067) );
  nnd4s1 U4175 ( .DIN1(n4070), .DIN2(n4071), .DIN3(n4072), .DIN4(n4073), 
        .Q(n3997) );
  nnd2s1 U4176 ( .DIN1(n3874), .DIN2(n4074), .Q(n4073) );
  nnd2s1 U4177 ( .DIN1(n3961), .DIN2(n3926), .Q(n4074) );
  nnd2s1 U4178 ( .DIN1(n3911), .DIN2(n4075), .Q(n4072) );
  nnd2s1 U4179 ( .DIN1(n4053), .DIN2(n4049), .Q(n4075) );
  nnd2s1 U4180 ( .DIN1(n3927), .DIN2(n4076), .Q(n4071) );
  nnd2s1 U4181 ( .DIN1(n3884), .DIN2(n4077), .Q(n4070) );
  nnd2s1 U4182 ( .DIN1(n4078), .DIN2(n4050), .Q(n4077) );
  nnd2s1 U4183 ( .DIN1(n4079), .DIN2(n4080), .Q(\u0/N111 ) );
  nnd2s1 U4184 ( .DIN1(\key[67] ), .DIN2(ld), .Q(n4080) );
  nnd2s1 U4185 ( .DIN1(n1994), .DIN2(n1569), .Q(n4079) );
  xnr2s1 U4186 ( .DIN1(w1[3]), .DIN2(n1770), .Q(n1994) );
  xnr2s1 U4187 ( .DIN1(n1505), .DIN2(n4081), .Q(n1770) );
  nor4s1 U4188 ( .DIN1(n4082), .DIN2(n4083), .DIN3(n4084), .DIN4(n4085), 
        .Q(n4081) );
  nnd3s1 U4189 ( .DIN1(n3943), .DIN2(n4027), .DIN3(n4001), .Q(n4085) );
  nor4s1 U4190 ( .DIN1(n4086), .DIN2(n4087), .DIN3(n4088), .DIN4(n4089), 
        .Q(n4001) );
  nnd4s1 U4191 ( .DIN1(n4090), .DIN2(n4091), .DIN3(n4092), .DIN4(n4093), 
        .Q(n4089) );
  nnd2s1 U4192 ( .DIN1(n3879), .DIN2(n3927), .Q(n4093) );
  nor2s1 U4193 ( .DIN1(n4094), .DIN2(n4095), .Q(n4092) );
  nor2s1 U4194 ( .DIN1(n3926), .DIN2(n4096), .Q(n4095) );
  nor2s1 U4195 ( .DIN1(n3988), .DIN2(n4097), .Q(n4094) );
  nnd2s1 U4196 ( .DIN1(n3869), .DIN2(n3955), .Q(n4091) );
  nnd2s1 U4197 ( .DIN1(n3962), .DIN2(n3892), .Q(n4090) );
  nnd3s1 U4198 ( .DIN1(n4098), .DIN2(n4099), .DIN3(n4100), .Q(n4088) );
  nnd2s1 U4199 ( .DIN1(n3989), .DIN2(n3993), .Q(n4100) );
  nnd2s1 U4200 ( .DIN1(n3877), .DIN2(n4101), .Q(n4099) );
  nnd3s1 U4201 ( .DIN1(n4052), .DIN2(n4019), .DIN3(n4096), .Q(n4101) );
  nnd2s1 U4202 ( .DIN1(n4033), .DIN2(n4102), .Q(n4098) );
  nnd3s1 U4203 ( .DIN1(n3950), .DIN2(n3891), .DIN3(n3925), .Q(n4102) );
  nor2s1 U4204 ( .DIN1(n3950), .DIN2(n3895), .Q(n4087) );
  nor2s1 U4205 ( .DIN1(n4103), .DIN2(n4104), .Q(n4086) );
  nor4s1 U4206 ( .DIN1(n4105), .DIN2(n4106), .DIN3(n4107), .DIN4(n4108), 
        .Q(n4027) );
  nnd4s1 U4207 ( .DIN1(n4109), .DIN2(n4110), .DIN3(n4111), .DIN4(n4112), 
        .Q(n4108) );
  nor2s1 U4208 ( .DIN1(n4113), .DIN2(n4114), .Q(n4112) );
  nor2s1 U4209 ( .DIN1(n4096), .DIN2(n4104), .Q(n4114) );
  nor2s1 U4210 ( .DIN1(n3992), .DIN2(n3891), .Q(n4113) );
  nnd2s1 U4211 ( .DIN1(n3912), .DIN2(n3896), .Q(n4110) );
  nnd2s1 U4212 ( .DIN1(n3965), .DIN2(n3876), .Q(n4109) );
  nnd3s1 U4213 ( .DIN1(n4115), .DIN2(n4116), .DIN3(n4117), .Q(n4107) );
  nnd2s1 U4214 ( .DIN1(n3953), .DIN2(n4118), .Q(n4117) );
  nnd2s1 U4215 ( .DIN1(n4053), .DIN2(n3968), .Q(n4118) );
  nnd2s1 U4216 ( .DIN1(n3911), .DIN2(n4119), .Q(n4116) );
  nnd2s1 U4217 ( .DIN1(n4078), .DIN2(n4019), .Q(n4119) );
  nnd2s1 U4218 ( .DIN1(n3878), .DIN2(n3990), .Q(n4115) );
  nnd2s1 U4219 ( .DIN1(n3970), .DIN2(n4120), .Q(n3990) );
  nor2s1 U4220 ( .DIN1(n4121), .DIN2(n3930), .Q(n4106) );
  nor2s1 U4221 ( .DIN1(n3867), .DIN2(n3888), .Q(n4121) );
  nor2s1 U4222 ( .DIN1(n4122), .DIN2(n4050), .Q(n4105) );
  and2s1 U4223 ( .DIN1(n3950), .DIN2(n4123), .Q(n4122) );
  nor4s1 U4224 ( .DIN1(n4124), .DIN2(n4125), .DIN3(n4126), .DIN4(n4127), 
        .Q(n3943) );
  nnd4s1 U4225 ( .DIN1(n4128), .DIN2(n4129), .DIN3(n4130), .DIN4(n4131), 
        .Q(n4127) );
  nnd2s1 U4226 ( .DIN1(n4032), .DIN2(n3955), .Q(n4131) );
  nor2s1 U4227 ( .DIN1(n4132), .DIN2(n4133), .Q(n4130) );
  nor2s1 U4228 ( .DIN1(n3930), .DIN2(n4134), .Q(n4132) );
  nnd2s1 U4229 ( .DIN1(n3954), .DIN2(n3962), .Q(n4129) );
  nnd2s1 U4230 ( .DIN1(n3952), .DIN2(n3884), .Q(n4128) );
  nnd3s1 U4231 ( .DIN1(n4135), .DIN2(n4136), .DIN3(n4137), .Q(n4126) );
  nnd2s1 U4232 ( .DIN1(n3876), .DIN2(n4138), .Q(n4137) );
  nnd2s1 U4233 ( .DIN1(n3892), .DIN2(n4139), .Q(n4136) );
  nnd2s1 U4234 ( .DIN1(n4050), .DIN2(n4019), .Q(n4139) );
  nnd2s1 U4235 ( .DIN1(n4033), .DIN2(n4140), .Q(n4135) );
  nnd3s1 U4236 ( .DIN1(n4021), .DIN2(n4104), .DIN3(n4141), .Q(n4140) );
  nor2s1 U4237 ( .DIN1(n3891), .DIN2(n3895), .Q(n4125) );
  nor2s1 U4238 ( .DIN1(n3932), .DIN2(n3887), .Q(n4124) );
  nnd3s1 U4239 ( .DIN1(n4142), .DIN2(n4143), .DIN3(n3910), .Q(n4084) );
  nor3s1 U4240 ( .DIN1(n4144), .DIN2(n4145), .DIN3(n4146), .Q(n3910) );
  nnd4s1 U4241 ( .DIN1(n4026), .DIN2(n3972), .DIN3(n4066), .DIN4(n4147), 
        .Q(n4146) );
  and3s1 U4242 ( .DIN1(n4148), .DIN2(n4149), .DIN3(n4150), .Q(n4147) );
  nnd2s1 U4243 ( .DIN1(n3952), .DIN2(n3875), .Q(n4150) );
  nnd2s1 U4244 ( .DIN1(n3866), .DIN2(n3927), .Q(n4148) );
  nor4s1 U4245 ( .DIN1(n4151), .DIN2(n4152), .DIN3(n4153), .DIN4(n4154), 
        .Q(n4066) );
  nnd4s1 U4246 ( .DIN1(n4155), .DIN2(n4156), .DIN3(n4157), .DIN4(n4158), 
        .Q(n4154) );
  nnd2s1 U4247 ( .DIN1(n3952), .DIN2(n4159), .Q(n4158) );
  nnd2s1 U4248 ( .DIN1(n4160), .DIN2(n4021), .Q(n4159) );
  nor2s1 U4249 ( .DIN1(n4161), .DIN2(n4162), .Q(n4157) );
  nor2s1 U4250 ( .DIN1(n4163), .DIN2(n3992), .Q(n4162) );
  nor2s1 U4251 ( .DIN1(n3866), .DIN2(n3934), .Q(n4163) );
  nor2s1 U4252 ( .DIN1(n4164), .DIN2(n3894), .Q(n4161) );
  nor2s1 U4253 ( .DIN1(n4022), .DIN2(n3965), .Q(n4164) );
  nnd2s1 U4254 ( .DIN1(n3884), .DIN2(n4165), .Q(n4156) );
  nnd3s1 U4255 ( .DIN1(n3895), .DIN2(n4049), .DIN3(n4134), .Q(n4165) );
  nnd2s1 U4256 ( .DIN1(n4033), .DIN2(n4022), .Q(n4155) );
  nnd3s1 U4257 ( .DIN1(n4166), .DIN2(n4167), .DIN3(n4168), .Q(n4153) );
  nnd2s1 U4258 ( .DIN1(n4169), .DIN2(n3989), .Q(n4168) );
  nnd2s1 U4259 ( .DIN1(n3874), .DIN2(n3877), .Q(n4167) );
  nnd2s1 U4260 ( .DIN1(n3878), .DIN2(n3911), .Q(n4166) );
  nor2s1 U4261 ( .DIN1(n4096), .DIN2(n3930), .Q(n4152) );
  nor2s1 U4262 ( .DIN1(n4104), .DIN2(n4078), .Q(n4151) );
  nor4s1 U4263 ( .DIN1(n4170), .DIN2(n4171), .DIN3(n4172), .DIN4(n4173), 
        .Q(n3972) );
  nnd4s1 U4264 ( .DIN1(n4174), .DIN2(n4175), .DIN3(n4176), .DIN4(n4177), 
        .Q(n4173) );
  nnd2s1 U4265 ( .DIN1(n3875), .DIN2(n3896), .Q(n4177) );
  nnd2s1 U4266 ( .DIN1(n3927), .DIN2(n3953), .Q(n4176) );
  nnd2s1 U4267 ( .DIN1(n3979), .DIN2(n3884), .Q(n4175) );
  nnd2s1 U4268 ( .DIN1(n3952), .DIN2(n3954), .Q(n4174) );
  nnd3s1 U4269 ( .DIN1(n4178), .DIN2(n4179), .DIN3(n4180), .Q(n4172) );
  nnd2s1 U4270 ( .DIN1(n3868), .DIN2(n4181), .Q(n4180) );
  nnd3s1 U4271 ( .DIN1(n3964), .DIN2(n3930), .DIN3(n4120), .Q(n4181) );
  nnd2s1 U4272 ( .DIN1(n3982), .DIN2(n4182), .Q(n4179) );
  nnd2s1 U4273 ( .DIN1(n4123), .DIN2(n3964), .Q(n4182) );
  nor2s1 U4274 ( .DIN1(n4169), .DIN2(n4022), .Q(n4123) );
  nnd2s1 U4275 ( .DIN1(n4032), .DIN2(n4183), .Q(n4178) );
  nnd2s1 U4276 ( .DIN1(n4097), .DIN2(n4078), .Q(n4183) );
  nor2s1 U4277 ( .DIN1(n4021), .DIN2(n4053), .Q(n4171) );
  nor2s1 U4278 ( .DIN1(n3971), .DIN2(n4050), .Q(n4170) );
  hi1s1 U4279 ( .DIN(n3897), .Q(n3971) );
  nor2s1 U4280 ( .DIN1(n4184), .DIN2(n4185), .Q(n4026) );
  nnd4s1 U4281 ( .DIN1(n4186), .DIN2(n4187), .DIN3(n4188), .DIN4(n4189), 
        .Q(n4185) );
  nnd2s1 U4282 ( .DIN1(n3875), .DIN2(n4190), .Q(n4189) );
  nnd3s1 U4283 ( .DIN1(n4050), .DIN2(n4096), .DIN3(n4134), .Q(n4190) );
  nnd2s1 U4284 ( .DIN1(n3874), .DIN2(n3965), .Q(n4187) );
  nnd4s1 U4285 ( .DIN1(n4191), .DIN2(n4192), .DIN3(n4193), .DIN4(n4194), 
        .Q(n4184) );
  nnd2s1 U4286 ( .DIN1(n3896), .DIN2(n4195), .Q(n4194) );
  nnd2s1 U4287 ( .DIN1(n4196), .DIN2(n3930), .Q(n4195) );
  nnd2s1 U4288 ( .DIN1(n3867), .DIN2(n4197), .Q(n4193) );
  nnd2s1 U4289 ( .DIN1(n3892), .DIN2(n4198), .Q(n4192) );
  nnd2s1 U4290 ( .DIN1(n4053), .DIN2(n4134), .Q(n4198) );
  nnd2s1 U4291 ( .DIN1(n4032), .DIN2(n4199), .Q(n4191) );
  nnd2s1 U4292 ( .DIN1(n3917), .DIN2(n4049), .Q(n4199) );
  nnd3s1 U4293 ( .DIN1(n4200), .DIN2(n4201), .DIN3(n4202), .Q(n4145) );
  nnd2s1 U4294 ( .DIN1(n3876), .DIN2(n3884), .Q(n4202) );
  nnd2s1 U4295 ( .DIN1(n4022), .DIN2(n4203), .Q(n4201) );
  nnd3s1 U4296 ( .DIN1(n4096), .DIN2(n3895), .DIN3(n4204), .Q(n4203) );
  or2s1 U4297 ( .DIN1(n3964), .DIN2(n4205), .Q(n4200) );
  nnd3s1 U4298 ( .DIN1(n4206), .DIN2(n4207), .DIN3(n4208), .Q(n4144) );
  nnd2s1 U4299 ( .DIN1(n3892), .DIN2(n4209), .Q(n4208) );
  nnd2s1 U4300 ( .DIN1(n4057), .DIN2(n4052), .Q(n4209) );
  nnd2s1 U4301 ( .DIN1(n3962), .DIN2(n4210), .Q(n4207) );
  or2s1 U4302 ( .DIN1(n3993), .DIN2(n3877), .Q(n4210) );
  nnd2s1 U4303 ( .DIN1(n3930), .DIN2(n3916), .Q(n3993) );
  nnd2s1 U4304 ( .DIN1(n3989), .DIN2(n4211), .Q(n4206) );
  nnd2s1 U4305 ( .DIN1(n3890), .DIN2(n3950), .Q(n4211) );
  nnd2s1 U4306 ( .DIN1(n3927), .DIN2(n3912), .Q(n4143) );
  nnd2s1 U4307 ( .DIN1(n3888), .DIN2(n3954), .Q(n4142) );
  nnd3s1 U4308 ( .DIN1(n4212), .DIN2(n4213), .DIN3(n4214), .Q(n4083) );
  nnd2s1 U4309 ( .DIN1(n4169), .DIN2(n3896), .Q(n4214) );
  nnd2s1 U4310 ( .DIN1(n4010), .DIN2(n4215), .Q(n4213) );
  nnd4s1 U4311 ( .DIN1(n4216), .DIN2(n4217), .DIN3(n4218), .DIN4(n4219), 
        .Q(n4082) );
  nnd2s1 U4312 ( .DIN1(n3982), .DIN2(n4220), .Q(n4219) );
  nnd2s1 U4313 ( .DIN1(n3932), .DIN2(n3988), .Q(n4220) );
  nor2s1 U4314 ( .DIN1(n3965), .DIN2(n3953), .Q(n3932) );
  nnd2s1 U4315 ( .DIN1(n3953), .DIN2(n4221), .Q(n4218) );
  nnd2s1 U4316 ( .DIN1(n3967), .DIN2(n4052), .Q(n4221) );
  nnd2s1 U4317 ( .DIN1(n3869), .DIN2(n4222), .Q(n4217) );
  nnd2s1 U4318 ( .DIN1(n3968), .DIN2(n3895), .Q(n4222) );
  nnd2s1 U4319 ( .DIN1(n3884), .DIN2(n4041), .Q(n4216) );
  nnd2s1 U4320 ( .DIN1(n4223), .DIN2(n4224), .Q(\u0/N110 ) );
  nnd2s1 U4321 ( .DIN1(\key[66] ), .DIN2(ld), .Q(n4224) );
  nnd2s1 U4322 ( .DIN1(n1997), .DIN2(n1569), .Q(n4223) );
  xnr2s1 U4323 ( .DIN1(w1[2]), .DIN2(n1773), .Q(n1997) );
  xor2s1 U4324 ( .DIN1(w0[2]), .DIN2(n4225), .Q(n1773) );
  nor4s1 U4325 ( .DIN1(n4226), .DIN2(n4227), .DIN3(n4228), .DIN4(n4229), 
        .Q(n4225) );
  nnd3s1 U4326 ( .DIN1(n4230), .DIN2(n4231), .DIN3(n4232), .Q(n4229) );
  nnd3s1 U4327 ( .DIN1(n4233), .DIN2(n4234), .DIN3(n3862), .Q(n4228) );
  nor3s1 U4328 ( .DIN1(n4235), .DIN2(n4236), .DIN3(n4237), .Q(n3862) );
  nnd4s1 U4329 ( .DIN1(n4238), .DIN2(n4239), .DIN3(n4240), .DIN4(n4241), 
        .Q(n4237) );
  and3s1 U4330 ( .DIN1(n4242), .DIN2(n4243), .DIN3(n4244), .Q(n4241) );
  nnd2s1 U4331 ( .DIN1(n3923), .DIN2(n3869), .Q(n4244) );
  nnd2s1 U4332 ( .DIN1(n3874), .DIN2(n3954), .Q(n4243) );
  nnd2s1 U4333 ( .DIN1(n3888), .DIN2(n3953), .Q(n4242) );
  nnd3s1 U4334 ( .DIN1(n4245), .DIN2(n4246), .DIN3(n4188), .Q(n4236) );
  nnd2s1 U4335 ( .DIN1(n3952), .DIN2(n4022), .Q(n4188) );
  or2s1 U4336 ( .DIN1(n3894), .DIN2(n4196), .Q(n4246) );
  nor2s1 U4337 ( .DIN1(n3866), .DIN2(n3877), .Q(n4196) );
  nnd2s1 U4338 ( .DIN1(n3982), .DIN2(n3934), .Q(n4245) );
  nnd2s1 U4339 ( .DIN1(n3970), .DIN2(n3925), .Q(n3934) );
  nnd4s1 U4340 ( .DIN1(n4247), .DIN2(n4248), .DIN3(n4249), .DIN4(n4250), 
        .Q(n4235) );
  nnd2s1 U4341 ( .DIN1(n4010), .DIN2(n4251), .Q(n4250) );
  nnd2s1 U4342 ( .DIN1(n3868), .DIN2(n4252), .Q(n4249) );
  nnd2s1 U4343 ( .DIN1(n3925), .DIN2(n3988), .Q(n4252) );
  nnd2s1 U4344 ( .DIN1(n3965), .DIN2(n4253), .Q(n4248) );
  nnd2s1 U4345 ( .DIN1(n3968), .DIN2(n3887), .Q(n4253) );
  nnd2s1 U4346 ( .DIN1(n3892), .DIN2(n4254), .Q(n4247) );
  nnd2s1 U4347 ( .DIN1(n4204), .DIN2(n4096), .Q(n4254) );
  hi1s1 U4348 ( .DIN(n3981), .Q(n4204) );
  nnd2s1 U4349 ( .DIN1(n4049), .DIN2(n3992), .Q(n3981) );
  nnd2s1 U4350 ( .DIN1(n3888), .DIN2(n3879), .Q(n4234) );
  nnd2s1 U4351 ( .DIN1(n3884), .DIN2(n3955), .Q(n4233) );
  nnd3s1 U4352 ( .DIN1(n4255), .DIN2(n4256), .DIN3(n4257), .Q(n4227) );
  nnd2s1 U4353 ( .DIN1(n3954), .DIN2(n3876), .Q(n4257) );
  or2s1 U4354 ( .DIN1(n3890), .DIN2(n3886), .Q(n4256) );
  nor2s1 U4355 ( .DIN1(n3923), .DIN2(n3927), .Q(n3886) );
  nnd2s1 U4356 ( .DIN1(n4032), .DIN2(n3896), .Q(n4255) );
  nnd4s1 U4357 ( .DIN1(n4258), .DIN2(n4259), .DIN3(n4260), .DIN4(n4261), 
        .Q(n4226) );
  nnd2s1 U4358 ( .DIN1(n4169), .DIN2(n4262), .Q(n4261) );
  nnd2s1 U4359 ( .DIN1(n4205), .DIN2(n4049), .Q(n4262) );
  nnd2s1 U4360 ( .DIN1(n3867), .DIN2(n4263), .Q(n4260) );
  nnd2s1 U4361 ( .DIN1(n4017), .DIN2(n3926), .Q(n4263) );
  nor2s1 U4362 ( .DIN1(n3875), .DIN2(n4022), .Q(n4017) );
  nnd2s1 U4363 ( .DIN1(n3868), .DIN2(n4264), .Q(n4259) );
  nnd2s1 U4364 ( .DIN1(n3869), .DIN2(n4251), .Q(n4258) );
  nnd2s1 U4365 ( .DIN1(n4053), .DIN2(n3887), .Q(n4251) );
  nnd2s1 U4366 ( .DIN1(n4265), .DIN2(n4266), .Q(\u0/N109 ) );
  nnd2s1 U4367 ( .DIN1(\key[65] ), .DIN2(ld), .Q(n4266) );
  nnd2s1 U4368 ( .DIN1(n2000), .DIN2(n1569), .Q(n4265) );
  xnr2s1 U4369 ( .DIN1(w1[1]), .DIN2(n1776), .Q(n2000) );
  xor2s1 U4370 ( .DIN1(w0[1]), .DIN2(n4267), .Q(n1776) );
  nor4s1 U4371 ( .DIN1(n4268), .DIN2(n4269), .DIN3(n4270), .DIN4(n4271), 
        .Q(n4267) );
  nnd3s1 U4372 ( .DIN1(n4232), .DIN2(n3859), .DIN3(n4272), .Q(n4271) );
  nor2s1 U4373 ( .DIN1(n4273), .DIN2(n4274), .Q(n3859) );
  nnd4s1 U4374 ( .DIN1(n4275), .DIN2(n4276), .DIN3(n4277), .DIN4(n4278), 
        .Q(n4274) );
  nnd2s1 U4375 ( .DIN1(n3879), .DIN2(n4041), .Q(n4278) );
  nnd2s1 U4376 ( .DIN1(n3968), .DIN2(n3894), .Q(n4041) );
  nnd2s1 U4377 ( .DIN1(n3875), .DIN2(n3876), .Q(n4277) );
  nnd2s1 U4378 ( .DIN1(n3868), .DIN2(n3965), .Q(n4276) );
  nnd2s1 U4379 ( .DIN1(n4032), .DIN2(n3989), .Q(n4275) );
  nnd4s1 U4380 ( .DIN1(n4279), .DIN2(n4280), .DIN3(n4281), .DIN4(n4282), 
        .Q(n4273) );
  nnd2s1 U4381 ( .DIN1(n3911), .DIN2(n4283), .Q(n4282) );
  or2s1 U4382 ( .DIN1(n4215), .DIN2(n3878), .Q(n4283) );
  nnd2s1 U4383 ( .DIN1(n3955), .DIN2(n4284), .Q(n4281) );
  nnd2s1 U4384 ( .DIN1(n3916), .DIN2(n3964), .Q(n4284) );
  nnd2s1 U4385 ( .DIN1(n3869), .DIN2(n4285), .Q(n4280) );
  nnd2s1 U4386 ( .DIN1(n4057), .DIN2(n3895), .Q(n4285) );
  nnd2s1 U4387 ( .DIN1(n3892), .DIN2(n4286), .Q(n4279) );
  nnd3s1 U4388 ( .DIN1(n4053), .DIN2(n4057), .DIN3(n4287), .Q(n4286) );
  nor4s1 U4389 ( .DIN1(n4288), .DIN2(n4289), .DIN3(n4290), .DIN4(n4291), 
        .Q(n4232) );
  nnd4s1 U4390 ( .DIN1(n4292), .DIN2(n4186), .DIN3(n4293), .DIN4(n4294), 
        .Q(n4291) );
  nnd2s1 U4391 ( .DIN1(n3979), .DIN2(n3897), .Q(n4294) );
  nnd2s1 U4392 ( .DIN1(n3982), .DIN2(n3869), .Q(n4293) );
  nnd2s1 U4393 ( .DIN1(n3878), .DIN2(n4169), .Q(n4186) );
  nnd2s1 U4394 ( .DIN1(n3923), .DIN2(n4010), .Q(n4292) );
  nnd3s1 U4395 ( .DIN1(n4295), .DIN2(n4296), .DIN3(n4297), .Q(n4290) );
  nnd2s1 U4396 ( .DIN1(n3884), .DIN2(n4298), .Q(n4297) );
  nnd2s1 U4397 ( .DIN1(n3874), .DIN2(n4299), .Q(n4296) );
  nnd2s1 U4398 ( .DIN1(n3929), .DIN2(n3926), .Q(n4299) );
  nnd2s1 U4399 ( .DIN1(n3912), .DIN2(n4300), .Q(n4295) );
  nnd2s1 U4400 ( .DIN1(n3917), .DIN2(n3894), .Q(n4300) );
  nor2s1 U4401 ( .DIN1(n4103), .DIN2(n3961), .Q(n4289) );
  nor2s1 U4402 ( .DIN1(n3989), .DIN2(n3982), .Q(n4103) );
  nor2s1 U4403 ( .DIN1(n4301), .DIN2(n4097), .Q(n4288) );
  nor2s1 U4404 ( .DIN1(n3965), .DIN2(n3954), .Q(n4301) );
  nnd3s1 U4405 ( .DIN1(n4302), .DIN2(n4064), .DIN3(n4239), .Q(n4270) );
  nor2s1 U4406 ( .DIN1(n4303), .DIN2(n4304), .Q(n4239) );
  nnd4s1 U4407 ( .DIN1(n4305), .DIN2(n4306), .DIN3(n4212), .DIN4(n4307), 
        .Q(n4304) );
  nnd2s1 U4408 ( .DIN1(n3912), .DIN2(n3919), .Q(n4307) );
  nnd2s1 U4409 ( .DIN1(n4078), .DIN2(n3895), .Q(n3919) );
  nnd2s1 U4410 ( .DIN1(n3923), .DIN2(n3877), .Q(n4212) );
  nnd2s1 U4411 ( .DIN1(n4033), .DIN2(n4010), .Q(n4306) );
  nnd2s1 U4412 ( .DIN1(n3869), .DIN2(n3927), .Q(n4305) );
  nnd4s1 U4413 ( .DIN1(n4308), .DIN2(n4309), .DIN3(n4310), .DIN4(n4311), 
        .Q(n4303) );
  nnd2s1 U4414 ( .DIN1(n3878), .DIN2(n4312), .Q(n4311) );
  nnd2s1 U4415 ( .DIN1(n4104), .DIN2(n4120), .Q(n4312) );
  nnd2s1 U4416 ( .DIN1(n3979), .DIN2(n4313), .Q(n4310) );
  nnd2s1 U4417 ( .DIN1(n3970), .DIN2(n3988), .Q(n4313) );
  nnd2s1 U4418 ( .DIN1(n3952), .DIN2(n4314), .Q(n4309) );
  nnd3s1 U4419 ( .DIN1(n3916), .DIN2(n3930), .DIN3(n3926), .Q(n4314) );
  nnd2s1 U4420 ( .DIN1(n3962), .DIN2(n4315), .Q(n4308) );
  nnd4s1 U4421 ( .DIN1(n3929), .DIN2(n3950), .DIN3(n4021), .DIN4(n3970), 
        .Q(n4315) );
  nnd2s1 U4422 ( .DIN1(n3879), .DIN2(n3979), .Q(n4064) );
  nnd2s1 U4423 ( .DIN1(n4033), .DIN2(n3892), .Q(n4302) );
  nnd3s1 U4424 ( .DIN1(n4316), .DIN2(n4317), .DIN3(n4318), .Q(n4269) );
  nnd2s1 U4425 ( .DIN1(n3923), .DIN2(n3953), .Q(n4318) );
  nnd2s1 U4426 ( .DIN1(n3878), .DIN2(n3875), .Q(n4317) );
  nnd2s1 U4427 ( .DIN1(n4010), .DIN2(n3867), .Q(n4316) );
  nnd4s1 U4428 ( .DIN1(n4319), .DIN2(n4320), .DIN3(n4321), .DIN4(n4322), 
        .Q(n4268) );
  nnd2s1 U4429 ( .DIN1(n4022), .DIN2(n4323), .Q(n4322) );
  nnd2s1 U4430 ( .DIN1(n4049), .DIN2(n4019), .Q(n4323) );
  nnd2s1 U4431 ( .DIN1(n3884), .DIN2(n4324), .Q(n4321) );
  nnd2s1 U4432 ( .DIN1(n4097), .DIN2(n4053), .Q(n4324) );
  nnd2s1 U4433 ( .DIN1(n3954), .DIN2(n4325), .Q(n4320) );
  nnd2s1 U4434 ( .DIN1(n3951), .DIN2(n4078), .Q(n4325) );
  nor2s1 U4435 ( .DIN1(n3868), .DIN2(n3982), .Q(n3951) );
  nnd2s1 U4436 ( .DIN1(n3965), .DIN2(n4326), .Q(n4319) );
  nnd3s1 U4437 ( .DIN1(n4050), .DIN2(n4052), .DIN3(n3917), .Q(n4326) );
  nor2s1 U4438 ( .DIN1(n3896), .DIN2(n3982), .Q(n3917) );
  nnd2s1 U4439 ( .DIN1(n4327), .DIN2(n4328), .Q(\u0/N108 ) );
  nnd2s1 U4440 ( .DIN1(\key[64] ), .DIN2(ld), .Q(n4328) );
  nnd2s1 U4441 ( .DIN1(n2003), .DIN2(n1569), .Q(n4327) );
  xnr2s1 U4442 ( .DIN1(w1[0]), .DIN2(n1779), .Q(n2003) );
  xnr2s1 U4443 ( .DIN1(n1473), .DIN2(n4329), .Q(n1779) );
  nor4s1 U4444 ( .DIN1(n4330), .DIN2(n4331), .DIN3(n4332), .DIN4(n4333), 
        .Q(n4329) );
  nnd3s1 U4445 ( .DIN1(n4231), .DIN2(n3861), .DIN3(n4272), .Q(n4333) );
  nor3s1 U4446 ( .DIN1(n4334), .DIN2(n4335), .DIN3(n4336), .Q(n4272) );
  nnd4s1 U4447 ( .DIN1(n3860), .DIN2(n4238), .DIN3(n4230), .DIN4(n4337), 
        .Q(n4336) );
  and3s1 U4448 ( .DIN1(n4338), .DIN2(n4339), .DIN3(n4340), .Q(n4337) );
  nnd2s1 U4449 ( .DIN1(n3954), .DIN2(n3979), .Q(n4340) );
  nnd2s1 U4450 ( .DIN1(n3869), .DIN2(n3962), .Q(n4339) );
  nnd2s1 U4451 ( .DIN1(n4033), .DIN2(n3884), .Q(n4338) );
  hi1s1 U4452 ( .DIN(n3970), .Q(n3884) );
  and4s1 U4453 ( .DIN1(n4341), .DIN2(n4342), .DIN3(n4343), .DIN4(n4344), 
        .Q(n4230) );
  and4s1 U4454 ( .DIN1(n4345), .DIN2(n4346), .DIN3(n4111), .DIN4(n4008), 
        .Q(n4344) );
  nnd2s1 U4455 ( .DIN1(n3878), .DIN2(n3912), .Q(n4008) );
  nnd2s1 U4456 ( .DIN1(n3952), .DIN2(n3866), .Q(n4111) );
  nnd2s1 U4457 ( .DIN1(n3923), .DIN2(n3892), .Q(n4346) );
  nnd2s1 U4458 ( .DIN1(n4033), .DIN2(n3954), .Q(n4345) );
  and3s1 U4459 ( .DIN1(n4347), .DIN2(n4348), .DIN3(n4349), .Q(n4343) );
  nnd2s1 U4460 ( .DIN1(n3879), .DIN2(n4298), .Q(n4349) );
  nnd2s1 U4461 ( .DIN1(n4019), .DIN2(n3992), .Q(n4298) );
  nnd2s1 U4462 ( .DIN1(n3876), .DIN2(n4350), .Q(n4348) );
  nnd2s1 U4463 ( .DIN1(n4141), .DIN2(n3970), .Q(n4350) );
  nor2s1 U4464 ( .DIN1(n4032), .DIN2(n4010), .Q(n4141) );
  nnd2s1 U4465 ( .DIN1(n4169), .DIN2(n4351), .Q(n4347) );
  nnd2s1 U4466 ( .DIN1(n4053), .DIN2(n3894), .Q(n4351) );
  nnd2s1 U4467 ( .DIN1(n4032), .DIN2(n4352), .Q(n4342) );
  nnd2s1 U4468 ( .DIN1(n4078), .DIN2(n3887), .Q(n4352) );
  nnd2s1 U4469 ( .DIN1(n3955), .DIN2(n4353), .Q(n4341) );
  nnd3s1 U4470 ( .DIN1(n3891), .DIN2(n3930), .DIN3(n3926), .Q(n4353) );
  nor4s1 U4471 ( .DIN1(n4354), .DIN2(n4355), .DIN3(n4356), .DIN4(n4357), 
        .Q(n4238) );
  nnd4s1 U4472 ( .DIN1(n4358), .DIN2(n4359), .DIN3(n4360), .DIN4(n4361), 
        .Q(n4357) );
  and3s1 U4473 ( .DIN1(n4362), .DIN2(n4363), .DIN3(n4364), .Q(n4361) );
  nnd2s1 U4474 ( .DIN1(n3874), .DIN2(n4022), .Q(n4364) );
  nnd2s1 U4475 ( .DIN1(n3875), .DIN2(n4365), .Q(n4363) );
  nnd2s1 U4476 ( .DIN1(n3968), .DIN2(n4366), .Q(n4365) );
  nnd2s1 U4477 ( .DIN1(n3888), .DIN2(n4264), .Q(n4362) );
  nnd2s1 U4478 ( .DIN1(n3961), .DIN2(n3964), .Q(n4264) );
  nnd2s1 U4479 ( .DIN1(n3867), .DIN2(n4367), .Q(n4360) );
  nnd2s1 U4480 ( .DIN1(n3929), .DIN2(n3988), .Q(n4367) );
  nnd2s1 U4481 ( .DIN1(n3877), .DIN2(n4368), .Q(n4359) );
  nnd2s1 U4482 ( .DIN1(n3887), .DIN2(n3895), .Q(n4368) );
  nnd2s1 U4483 ( .DIN1(n4169), .DIN2(n4369), .Q(n4358) );
  nnd2s1 U4484 ( .DIN1(n4096), .DIN2(n4097), .Q(n4369) );
  nnd3s1 U4485 ( .DIN1(n4370), .DIN2(n4371), .DIN3(n4372), .Q(n4356) );
  nnd2s1 U4486 ( .DIN1(n3989), .DIN2(n3953), .Q(n4372) );
  nnd2s1 U4487 ( .DIN1(n3982), .DIN2(n3911), .Q(n4371) );
  nnd2s1 U4488 ( .DIN1(n3879), .DIN2(n3896), .Q(n4370) );
  nor2s1 U4489 ( .DIN1(n4050), .DIN2(n4160), .Q(n4355) );
  nor2s1 U4490 ( .DIN1(n3961), .DIN2(n4078), .Q(n4354) );
  nor4s1 U4491 ( .DIN1(n4373), .DIN2(n4374), .DIN3(n4375), .DIN4(n4376), 
        .Q(n3860) );
  nnd4s1 U4492 ( .DIN1(n4377), .DIN2(n4378), .DIN3(n4379), .DIN4(n4380), 
        .Q(n4376) );
  nnd2s1 U4493 ( .DIN1(n3982), .DIN2(n3875), .Q(n4380) );
  nnd2s1 U4494 ( .DIN1(n3868), .DIN2(n3877), .Q(n4379) );
  nnd2s1 U4495 ( .DIN1(n3911), .DIN2(n3896), .Q(n4378) );
  hi1s1 U4496 ( .DIN(n3988), .Q(n3911) );
  nnd2s1 U4497 ( .DIN1(n3866), .DIN2(n3876), .Q(n4377) );
  nnd3s1 U4498 ( .DIN1(n4381), .DIN2(n4382), .DIN3(n4383), .Q(n4375) );
  nnd2s1 U4499 ( .DIN1(n3954), .DIN2(n4384), .Q(n4383) );
  nnd3s1 U4500 ( .DIN1(n4366), .DIN2(n3992), .DIN3(n4050), .Q(n4384) );
  nnd2s1 U4501 ( .DIN1(n3879), .DIN2(n4385), .Q(n4382) );
  nnd2s1 U4502 ( .DIN1(n4049), .DIN2(n4134), .Q(n4385) );
  hi1s1 U4503 ( .DIN(n3916), .Q(n3879) );
  nnd2s1 U4504 ( .DIN1(n3979), .DIN2(n4386), .Q(n4381) );
  nnd2s1 U4505 ( .DIN1(n3890), .DIN2(n4120), .Q(n4386) );
  nor2s1 U4506 ( .DIN1(n3970), .DIN2(n3895), .Q(n4374) );
  and2s1 U4507 ( .DIN1(n4033), .DIN2(n4387), .Q(n4373) );
  nnd4s1 U4508 ( .DIN1(n3988), .DIN2(n3929), .DIN3(n3926), .DIN4(n3930), 
        .Q(n4387) );
  nnd3s1 U4509 ( .DIN1(n4388), .DIN2(n4389), .DIN3(n4390), .Q(n4335) );
  nnd2s1 U4510 ( .DIN1(n3923), .DIN2(n3875), .Q(n4390) );
  nnd2s1 U4511 ( .DIN1(n4169), .DIN2(n3874), .Q(n4389) );
  nnd2s1 U4512 ( .DIN1(n3952), .DIN2(n3912), .Q(n4388) );
  nnd4s1 U4513 ( .DIN1(n4391), .DIN2(n4392), .DIN3(n4393), .DIN4(n4394), 
        .Q(n4334) );
  nnd2s1 U4514 ( .DIN1(n4022), .DIN2(n4395), .Q(n4394) );
  nnd2s1 U4515 ( .DIN1(n4057), .DIN2(n3894), .Q(n4395) );
  nnd2s1 U4516 ( .DIN1(n4032), .DIN2(n4396), .Q(n4393) );
  nnd4s1 U4517 ( .DIN1(n4134), .DIN2(n4097), .DIN3(n4050), .DIN4(n4057), 
        .Q(n4396) );
  nnd2s1 U4518 ( .DIN1(n3989), .DIN2(n4138), .Q(n4392) );
  nnd2s1 U4519 ( .DIN1(n4104), .DIN2(n3891), .Q(n4138) );
  nnd2s1 U4520 ( .DIN1(n3876), .DIN2(n4042), .Q(n4391) );
  nnd2s1 U4521 ( .DIN1(n3916), .DIN2(n3925), .Q(n4042) );
  nor4s1 U4522 ( .DIN1(n4397), .DIN2(n4398), .DIN3(n4399), .DIN4(n4400), 
        .Q(n3861) );
  nnd4s1 U4523 ( .DIN1(n4401), .DIN2(n4402), .DIN3(n4403), .DIN4(n4404), 
        .Q(n4400) );
  nnd2s1 U4524 ( .DIN1(n3892), .DIN2(n3876), .Q(n4404) );
  nor2s1 U4525 ( .DIN1(n4405), .DIN2(n4133), .Q(n4403) );
  nor2s1 U4526 ( .DIN1(n3964), .DIN2(n3894), .Q(n4133) );
  nor2s1 U4527 ( .DIN1(n3950), .DIN2(n3992), .Q(n4405) );
  nnd2s1 U4528 ( .DIN1(n3875), .DIN2(n3979), .Q(n4402) );
  hi1s1 U4529 ( .DIN(n3891), .Q(n3875) );
  nnd2s1 U4530 ( .DIN1(n3962), .DIN2(n3965), .Q(n4401) );
  nnd3s1 U4531 ( .DIN1(n4406), .DIN2(n4407), .DIN3(n4408), .Q(n4399) );
  nnd2s1 U4532 ( .DIN1(n3955), .DIN2(n4040), .Q(n4408) );
  nnd2s1 U4533 ( .DIN1(n3961), .DIN2(n3950), .Q(n4040) );
  nnd2s1 U4534 ( .DIN1(n3877), .DIN2(n4409), .Q(n4407) );
  nnd3s1 U4535 ( .DIN1(n4050), .DIN2(n4057), .DIN3(n4097), .Q(n4409) );
  nnd2s1 U4536 ( .DIN1(n3953), .DIN2(n4410), .Q(n4406) );
  nnd3s1 U4537 ( .DIN1(n4366), .DIN2(n4052), .DIN3(n4096), .Q(n4410) );
  nor2s1 U4538 ( .DIN1(n4366), .DIN2(n3970), .Q(n4398) );
  nnd2s1 U4539 ( .DIN1(n4411), .DIN2(n4412), .Q(n3970) );
  nor2s1 U4540 ( .DIN1(n4205), .DIN2(n4120), .Q(n4397) );
  nor2s1 U4541 ( .DIN1(n3923), .DIN2(n3896), .Q(n4205) );
  nor4s1 U4542 ( .DIN1(n4413), .DIN2(n4414), .DIN3(n4415), .DIN4(n4416), 
        .Q(n4231) );
  nnd4s1 U4543 ( .DIN1(n4417), .DIN2(n4418), .DIN3(n4419), .DIN4(n4420), 
        .Q(n4416) );
  nnd2s1 U4544 ( .DIN1(n3962), .DIN2(n4010), .Q(n4420) );
  nor2s1 U4545 ( .DIN1(n4421), .DIN2(n4422), .Q(n4419) );
  nor2s1 U4546 ( .DIN1(n3895), .DIN2(n3961), .Q(n4422) );
  nor2s1 U4547 ( .DIN1(n4015), .DIN2(n4134), .Q(n4421) );
  nor2s1 U4548 ( .DIN1(n3892), .DIN2(n4010), .Q(n4015) );
  hi1s1 U4549 ( .DIN(n3964), .Q(n4010) );
  nnd2s1 U4550 ( .DIN1(n3869), .DIN2(n3876), .Q(n4418) );
  hi1s1 U4551 ( .DIN(n3930), .Q(n3869) );
  nnd2s1 U4552 ( .DIN1(n4169), .DIN2(n3955), .Q(n4417) );
  nnd3s1 U4553 ( .DIN1(n4423), .DIN2(n4424), .DIN3(n4425), .Q(n4415) );
  nnd2s1 U4554 ( .DIN1(n3867), .DIN2(n4076), .Q(n4425) );
  nnd2s1 U4555 ( .DIN1(n3925), .DIN2(n4021), .Q(n4076) );
  nnd2s1 U4556 ( .DIN1(n3912), .DIN2(n4426), .Q(n4424) );
  nnd2s1 U4557 ( .DIN1(n4096), .DIN2(n3968), .Q(n4426) );
  nnd2s1 U4558 ( .DIN1(n3953), .DIN2(n4427), .Q(n4423) );
  nnd2s1 U4559 ( .DIN1(n3887), .DIN2(n4134), .Q(n4427) );
  hi1s1 U4560 ( .DIN(n3926), .Q(n3953) );
  nor2s1 U4561 ( .DIN1(n4428), .DIN2(n3891), .Q(n4414) );
  nor2s1 U4562 ( .DIN1(n3868), .DIN2(n3952), .Q(n4428) );
  nor2s1 U4563 ( .DIN1(n4429), .DIN2(n3916), .Q(n4413) );
  nnd2s1 U4564 ( .DIN1(n4411), .DIN2(n4430), .Q(n3916) );
  nor2s1 U4565 ( .DIN1(n3874), .DIN2(n3923), .Q(n4429) );
  hi1s1 U4566 ( .DIN(n4078), .Q(n3923) );
  nnd3s1 U4567 ( .DIN1(w3[26]), .DIN2(n1554), .DIN3(n4431), .Q(n4078) );
  hi1s1 U4568 ( .DIN(n3895), .Q(n3874) );
  nnd4s1 U4569 ( .DIN1(n4240), .DIN2(n4432), .DIN3(n4433), .DIN4(n4434), 
        .Q(n4332) );
  nnd2s1 U4570 ( .DIN1(n3866), .DIN2(n3962), .Q(n4434) );
  hi1s1 U4571 ( .DIN(n4049), .Q(n3962) );
  hi1s1 U4572 ( .DIN(n3961), .Q(n3866) );
  nnd2s1 U4573 ( .DIN1(n3952), .DIN2(n3892), .Q(n4433) );
  nnd2s1 U4574 ( .DIN1(n4032), .DIN2(n3979), .Q(n4432) );
  hi1s1 U4575 ( .DIN(n3929), .Q(n4032) );
  and4s1 U4576 ( .DIN1(n4435), .DIN2(n4436), .DIN3(n4437), .DIN4(n4438), 
        .Q(n4240) );
  and4s1 U4577 ( .DIN1(n4439), .DIN2(n4149), .DIN3(n4440), .DIN4(n4441), 
        .Q(n4438) );
  nnd2s1 U4578 ( .DIN1(n3982), .DIN2(n4022), .Q(n4441) );
  nnd2s1 U4579 ( .DIN1(n3876), .DIN2(n3912), .Q(n4440) );
  hi1s1 U4580 ( .DIN(n3950), .Q(n3912) );
  hi1s1 U4581 ( .DIN(n4052), .Q(n3876) );
  nnd3s1 U4582 ( .DIN1(n1554), .DIN2(n1548), .DIN3(n4431), .Q(n4052) );
  nnd2s1 U4583 ( .DIN1(n3888), .DIN2(n4169), .Q(n4149) );
  hi1s1 U4584 ( .DIN(n3925), .Q(n4169) );
  nnd2s1 U4585 ( .DIN1(n3868), .DIN2(n3892), .Q(n4439) );
  hi1s1 U4586 ( .DIN(n4160), .Q(n3892) );
  nnd2s1 U4587 ( .DIN1(n4411), .DIN2(n4442), .Q(n4160) );
  and3s1 U4588 ( .DIN1(n4443), .DIN2(n4444), .DIN3(n4445), .Q(n4437) );
  nnd2s1 U4589 ( .DIN1(n3979), .DIN2(n4446), .Q(n4445) );
  nnd2s1 U4590 ( .DIN1(n3930), .DIN2(n3961), .Q(n4446) );
  hi1s1 U4591 ( .DIN(n4096), .Q(n3979) );
  nnd3s1 U4592 ( .DIN1(n4447), .DIN2(n1410), .DIN3(w3[24]), .Q(n4096) );
  nnd2s1 U4593 ( .DIN1(n3867), .DIN2(n4448), .Q(n4444) );
  nnd2s1 U4594 ( .DIN1(n3890), .DIN2(n3930), .Q(n4448) );
  nnd2s1 U4595 ( .DIN1(n4412), .DIN2(n4449), .Q(n3930) );
  hi1s1 U4596 ( .DIN(n3992), .Q(n3867) );
  nnd3s1 U4597 ( .DIN1(w3[24]), .DIN2(n1410), .DIN3(n4450), .Q(n3992) );
  nnd2s1 U4598 ( .DIN1(n3952), .DIN2(n4197), .Q(n4443) );
  nnd2s1 U4599 ( .DIN1(n3964), .DIN2(n3988), .Q(n4197) );
  hi1s1 U4600 ( .DIN(n4097), .Q(n3952) );
  nnd3s1 U4601 ( .DIN1(w3[24]), .DIN2(n4451), .DIN3(w3[26]), .Q(n4097) );
  nnd2s1 U4602 ( .DIN1(n3927), .DIN2(n4452), .Q(n4436) );
  nnd3s1 U4603 ( .DIN1(n3929), .DIN2(n3891), .DIN3(n3988), .Q(n4452) );
  nnd2s1 U4604 ( .DIN1(n4430), .DIN2(n4449), .Q(n3891) );
  nnd2s1 U4605 ( .DIN1(n4442), .DIN2(n4453), .Q(n3929) );
  hi1s1 U4606 ( .DIN(n3894), .Q(n3927) );
  nnd3s1 U4607 ( .DIN1(w3[26]), .DIN2(w3[24]), .DIN3(n4431), .Q(n3894) );
  or2s1 U4608 ( .DIN1(n3961), .DIN2(n4287), .Q(n4435) );
  nor2s1 U4609 ( .DIN1(n3878), .DIN2(n3896), .Q(n4287) );
  hi1s1 U4610 ( .DIN(n4366), .Q(n3896) );
  nnd3s1 U4611 ( .DIN1(n4451), .DIN2(n1548), .DIN3(w3[24]), .Q(n4366) );
  hi1s1 U4612 ( .DIN(n3887), .Q(n3878) );
  nnd3s1 U4613 ( .DIN1(n4447), .DIN2(n1554), .DIN3(w3[25]), .Q(n3887) );
  nnd4s1 U4614 ( .DIN1(n4065), .DIN2(n4454), .DIN3(n4455), .DIN4(n4456), 
        .Q(n4331) );
  nnd2s1 U4615 ( .DIN1(n3965), .DIN2(n4215), .Q(n4456) );
  nnd2s1 U4616 ( .DIN1(n4053), .DIN2(n3895), .Q(n4215) );
  nnd3s1 U4617 ( .DIN1(w3[25]), .DIN2(w3[24]), .DIN3(n4450), .Q(n3895) );
  hi1s1 U4618 ( .DIN(n3890), .Q(n3965) );
  nnd2s1 U4619 ( .DIN1(n4453), .DIN2(n4457), .Q(n3890) );
  nnd2s1 U4620 ( .DIN1(n3989), .DIN2(n3897), .Q(n4455) );
  nnd2s1 U4621 ( .DIN1(n3964), .DIN2(n4021), .Q(n3897) );
  nnd2s1 U4622 ( .DIN1(n4411), .DIN2(n4457), .Q(n3964) );
  nor2s1 U4623 ( .DIN1(n1392), .DIN2(w3[30]), .Q(n4411) );
  hi1s1 U4624 ( .DIN(n4053), .Q(n3989) );
  nnd3s1 U4625 ( .DIN1(n4451), .DIN2(n1554), .DIN3(w3[26]), .Q(n4053) );
  nnd2s1 U4626 ( .DIN1(n4022), .DIN2(n3955), .Q(n4454) );
  hi1s1 U4627 ( .DIN(n4120), .Q(n4022) );
  nnd2s1 U4628 ( .DIN1(n4442), .DIN2(n4458), .Q(n4120) );
  nnd2s1 U4629 ( .DIN1(n3982), .DIN2(n3877), .Q(n4065) );
  hi1s1 U4630 ( .DIN(n4021), .Q(n3877) );
  nnd2s1 U4631 ( .DIN1(n4449), .DIN2(n4457), .Q(n4021) );
  hi1s1 U4632 ( .DIN(n4134), .Q(n3982) );
  nnd3s1 U4633 ( .DIN1(w3[24]), .DIN2(n1548), .DIN3(n4431), .Q(n4134) );
  nor2s1 U4634 ( .DIN1(n1410), .DIN2(w3[27]), .Q(n4431) );
  nnd4s1 U4635 ( .DIN1(n4459), .DIN2(n4460), .DIN3(n4461), .DIN4(n4462), 
        .Q(n4330) );
  nnd2s1 U4636 ( .DIN1(n3868), .DIN2(n4463), .Q(n4462) );
  nnd2s1 U4637 ( .DIN1(n3926), .DIN2(n3950), .Q(n4463) );
  nnd2s1 U4638 ( .DIN1(n4412), .DIN2(n4458), .Q(n3950) );
  nnd2s1 U4639 ( .DIN1(n4458), .DIN2(n4457), .Q(n3926) );
  nor2s1 U4640 ( .DIN1(n1416), .DIN2(n1374), .Q(n4457) );
  hi1s1 U4641 ( .DIN(n4019), .Q(n3868) );
  nnd3s1 U4642 ( .DIN1(n1554), .DIN2(n1410), .DIN3(n4447), .Q(n4019) );
  nnd2s1 U4643 ( .DIN1(n3954), .DIN2(n4464), .Q(n4461) );
  nnd2s1 U4644 ( .DIN1(n4057), .DIN2(n4049), .Q(n4464) );
  nnd3s1 U4645 ( .DIN1(n1554), .DIN2(n1410), .DIN3(n4450), .Q(n4049) );
  hi1s1 U4646 ( .DIN(n4104), .Q(n3954) );
  nnd2s1 U4647 ( .DIN1(n4442), .DIN2(n4449), .Q(n4104) );
  nor2s1 U4648 ( .DIN1(n1475), .DIN2(w3[28]), .Q(n4449) );
  nor2s1 U4649 ( .DIN1(w3[31]), .DIN2(w3[29]), .Q(n4442) );
  or2s1 U4650 ( .DIN1(n3988), .DIN2(n3967), .Q(n4460) );
  nor2s1 U4651 ( .DIN1(n3888), .DIN2(n3955), .Q(n3967) );
  hi1s1 U4652 ( .DIN(n4050), .Q(n3955) );
  nnd3s1 U4653 ( .DIN1(w3[24]), .DIN2(n4447), .DIN3(w3[25]), .Q(n4050) );
  nor2s1 U4654 ( .DIN1(n1476), .DIN2(w3[26]), .Q(n4447) );
  hi1s1 U4655 ( .DIN(n4057), .Q(n3888) );
  nnd3s1 U4656 ( .DIN1(n1554), .DIN2(n1548), .DIN3(n4451), .Q(n4057) );
  nor2s1 U4657 ( .DIN1(w3[27]), .DIN2(w3[25]), .Q(n4451) );
  nnd2s1 U4658 ( .DIN1(n4430), .DIN2(n4458), .Q(n3988) );
  nor2s1 U4659 ( .DIN1(n1392), .DIN2(n1475), .Q(n4458) );
  nnd2s1 U4660 ( .DIN1(n4033), .DIN2(n3980), .Q(n4459) );
  nnd2s1 U4661 ( .DIN1(n3961), .DIN2(n3925), .Q(n3980) );
  nnd2s1 U4662 ( .DIN1(n4453), .DIN2(n4412), .Q(n3925) );
  nor2s1 U4663 ( .DIN1(n1416), .DIN2(w3[29]), .Q(n4412) );
  nnd2s1 U4664 ( .DIN1(n4430), .DIN2(n4453), .Q(n3961) );
  nor2s1 U4665 ( .DIN1(w3[30]), .DIN2(w3[28]), .Q(n4453) );
  nor2s1 U4666 ( .DIN1(n1374), .DIN2(w3[31]), .Q(n4430) );
  hi1s1 U4667 ( .DIN(n3968), .Q(n4033) );
  nnd3s1 U4668 ( .DIN1(w3[25]), .DIN2(n1554), .DIN3(n4450), .Q(n3968) );
  nor2s1 U4669 ( .DIN1(n1548), .DIN2(n1476), .Q(n4450) );
  nnd2s1 U4670 ( .DIN1(n4465), .DIN2(n4466), .Q(n1354) );
  nnd2s1 U4671 ( .DIN1(n4467), .DIN2(n1449), .Q(n4466) );
  nnd2s1 U4672 ( .DIN1(n4465), .DIN2(n4468), .Q(n1353) );
  nnd3s1 U4673 ( .DIN1(n4467), .DIN2(n4469), .DIN3(n15578), .Q(n4468) );
  nnd2s1 U4674 ( .DIN1(n4465), .DIN2(n4470), .Q(n1352) );
  nnd2s1 U4675 ( .DIN1(n4471), .DIN2(n4467), .Q(n4470) );
  hi1s1 U4676 ( .DIN(n4472), .Q(n4467) );
  xor2s1 U4677 ( .DIN1(n1449), .DIN2(n15577), .Q(n4471) );
  nnd2s1 U4678 ( .DIN1(rst), .DIN2(ld), .Q(n4465) );
  nor2s1 U4679 ( .DIN1(n4473), .DIN2(n4472), .Q(n1351) );
  nnd3s1 U4680 ( .DIN1(n4474), .DIN2(n1560), .DIN3(rst), .Q(n4472) );
  nnd2s1 U4681 ( .DIN1(n4475), .DIN2(n1526), .Q(n4474) );
  nor2s1 U4682 ( .DIN1(n4476), .DIN2(n4475), .Q(n4473) );
  hi1s1 U4683 ( .DIN(n4469), .Q(n4475) );
  nnd3s1 U4684 ( .DIN1(n1360), .DIN2(n1409), .DIN3(n1449), .Q(n4469) );
  nor2s1 U4685 ( .DIN1(n4477), .DIN2(n1360), .Q(n4476) );
  nor2s1 U4686 ( .DIN1(n15579), .DIN2(n15577), .Q(n4477) );
  nnd2s1 U4687 ( .DIN1(n4478), .DIN2(n4479), .Q(n1346) );
  nnd2s1 U4688 ( .DIN1(text_in_r[127]), .DIN2(n1570), .Q(n4479) );
  nnd2s1 U4689 ( .DIN1(\text_in[127] ), .DIN2(ld), .Q(n4478) );
  nnd2s1 U4690 ( .DIN1(n4480), .DIN2(n4481), .Q(n1345) );
  nnd2s1 U4691 ( .DIN1(text_in_r[126]), .DIN2(n1570), .Q(n4481) );
  nnd2s1 U4692 ( .DIN1(\text_in[126] ), .DIN2(ld), .Q(n4480) );
  nnd2s1 U4693 ( .DIN1(n4482), .DIN2(n4483), .Q(n1344) );
  nnd2s1 U4694 ( .DIN1(text_in_r[125]), .DIN2(n1570), .Q(n4483) );
  nnd2s1 U4695 ( .DIN1(\text_in[125] ), .DIN2(ld), .Q(n4482) );
  nnd2s1 U4696 ( .DIN1(n4484), .DIN2(n4485), .Q(n1343) );
  nnd2s1 U4697 ( .DIN1(text_in_r[124]), .DIN2(n1570), .Q(n4485) );
  nnd2s1 U4698 ( .DIN1(\text_in[124] ), .DIN2(ld), .Q(n4484) );
  nnd2s1 U4699 ( .DIN1(n4486), .DIN2(n4487), .Q(n1342) );
  nnd2s1 U4700 ( .DIN1(text_in_r[123]), .DIN2(n1570), .Q(n4487) );
  nnd2s1 U4701 ( .DIN1(\text_in[123] ), .DIN2(ld), .Q(n4486) );
  nnd2s1 U4702 ( .DIN1(n4488), .DIN2(n4489), .Q(n1341) );
  nnd2s1 U4703 ( .DIN1(text_in_r[122]), .DIN2(n1570), .Q(n4489) );
  nnd2s1 U4704 ( .DIN1(\text_in[122] ), .DIN2(ld), .Q(n4488) );
  nnd2s1 U4705 ( .DIN1(n4490), .DIN2(n4491), .Q(n1340) );
  nnd2s1 U4706 ( .DIN1(text_in_r[121]), .DIN2(n1570), .Q(n4491) );
  nnd2s1 U4707 ( .DIN1(\text_in[121] ), .DIN2(ld), .Q(n4490) );
  nnd2s1 U4708 ( .DIN1(n4492), .DIN2(n4493), .Q(n1339) );
  nnd2s1 U4709 ( .DIN1(text_in_r[120]), .DIN2(n1571), .Q(n4493) );
  nnd2s1 U4710 ( .DIN1(\text_in[120] ), .DIN2(ld), .Q(n4492) );
  nnd2s1 U4711 ( .DIN1(n4494), .DIN2(n4495), .Q(n1338) );
  nnd2s1 U4712 ( .DIN1(text_in_r[119]), .DIN2(n1571), .Q(n4495) );
  nnd2s1 U4713 ( .DIN1(\text_in[119] ), .DIN2(ld), .Q(n4494) );
  nnd2s1 U4714 ( .DIN1(n4496), .DIN2(n4497), .Q(n1337) );
  nnd2s1 U4715 ( .DIN1(text_in_r[118]), .DIN2(n1571), .Q(n4497) );
  nnd2s1 U4716 ( .DIN1(\text_in[118] ), .DIN2(ld), .Q(n4496) );
  nnd2s1 U4717 ( .DIN1(n4498), .DIN2(n4499), .Q(n1336) );
  nnd2s1 U4718 ( .DIN1(text_in_r[117]), .DIN2(n1571), .Q(n4499) );
  nnd2s1 U4719 ( .DIN1(\text_in[117] ), .DIN2(ld), .Q(n4498) );
  nnd2s1 U4720 ( .DIN1(n4500), .DIN2(n4501), .Q(n1335) );
  nnd2s1 U4721 ( .DIN1(text_in_r[116]), .DIN2(n1571), .Q(n4501) );
  nnd2s1 U4722 ( .DIN1(\text_in[116] ), .DIN2(ld), .Q(n4500) );
  nnd2s1 U4723 ( .DIN1(n4502), .DIN2(n4503), .Q(n1334) );
  nnd2s1 U4724 ( .DIN1(text_in_r[115]), .DIN2(n1571), .Q(n4503) );
  nnd2s1 U4725 ( .DIN1(\text_in[115] ), .DIN2(ld), .Q(n4502) );
  nnd2s1 U4726 ( .DIN1(n4504), .DIN2(n4505), .Q(n1333) );
  nnd2s1 U4727 ( .DIN1(text_in_r[114]), .DIN2(n1571), .Q(n4505) );
  nnd2s1 U4728 ( .DIN1(\text_in[114] ), .DIN2(ld), .Q(n4504) );
  nnd2s1 U4729 ( .DIN1(n4506), .DIN2(n4507), .Q(n1332) );
  nnd2s1 U4730 ( .DIN1(text_in_r[113]), .DIN2(n1572), .Q(n4507) );
  nnd2s1 U4731 ( .DIN1(\text_in[113] ), .DIN2(ld), .Q(n4506) );
  nnd2s1 U4732 ( .DIN1(n4508), .DIN2(n4509), .Q(n1331) );
  nnd2s1 U4733 ( .DIN1(text_in_r[112]), .DIN2(n1572), .Q(n4509) );
  nnd2s1 U4734 ( .DIN1(\text_in[112] ), .DIN2(ld), .Q(n4508) );
  nnd2s1 U4735 ( .DIN1(n4510), .DIN2(n4511), .Q(n1330) );
  nnd2s1 U4736 ( .DIN1(text_in_r[111]), .DIN2(n1572), .Q(n4511) );
  nnd2s1 U4737 ( .DIN1(\text_in[111] ), .DIN2(ld), .Q(n4510) );
  nnd2s1 U4738 ( .DIN1(n4512), .DIN2(n4513), .Q(n1329) );
  nnd2s1 U4739 ( .DIN1(text_in_r[110]), .DIN2(n1572), .Q(n4513) );
  nnd2s1 U4740 ( .DIN1(\text_in[110] ), .DIN2(ld), .Q(n4512) );
  nnd2s1 U4741 ( .DIN1(n4514), .DIN2(n4515), .Q(n1328) );
  nnd2s1 U4742 ( .DIN1(text_in_r[109]), .DIN2(n1572), .Q(n4515) );
  nnd2s1 U4743 ( .DIN1(\text_in[109] ), .DIN2(ld), .Q(n4514) );
  nnd2s1 U4744 ( .DIN1(n4516), .DIN2(n4517), .Q(n1327) );
  nnd2s1 U4745 ( .DIN1(text_in_r[108]), .DIN2(n1572), .Q(n4517) );
  nnd2s1 U4746 ( .DIN1(\text_in[108] ), .DIN2(ld), .Q(n4516) );
  nnd2s1 U4747 ( .DIN1(n4518), .DIN2(n4519), .Q(n1326) );
  nnd2s1 U4748 ( .DIN1(text_in_r[107]), .DIN2(n1572), .Q(n4519) );
  nnd2s1 U4749 ( .DIN1(\text_in[107] ), .DIN2(ld), .Q(n4518) );
  nnd2s1 U4750 ( .DIN1(n4520), .DIN2(n4521), .Q(n1325) );
  nnd2s1 U4751 ( .DIN1(text_in_r[106]), .DIN2(n1573), .Q(n4521) );
  nnd2s1 U4752 ( .DIN1(\text_in[106] ), .DIN2(ld), .Q(n4520) );
  nnd2s1 U4753 ( .DIN1(n4522), .DIN2(n4523), .Q(n1324) );
  nnd2s1 U4754 ( .DIN1(text_in_r[105]), .DIN2(n1573), .Q(n4523) );
  nnd2s1 U4755 ( .DIN1(\text_in[105] ), .DIN2(ld), .Q(n4522) );
  nnd2s1 U4756 ( .DIN1(n4524), .DIN2(n4525), .Q(n1323) );
  nnd2s1 U4757 ( .DIN1(text_in_r[104]), .DIN2(n1573), .Q(n4525) );
  nnd2s1 U4758 ( .DIN1(\text_in[104] ), .DIN2(ld), .Q(n4524) );
  nnd2s1 U4759 ( .DIN1(n4526), .DIN2(n4527), .Q(n1322) );
  nnd2s1 U4760 ( .DIN1(text_in_r[103]), .DIN2(n1573), .Q(n4527) );
  nnd2s1 U4761 ( .DIN1(\text_in[103] ), .DIN2(ld), .Q(n4526) );
  nnd2s1 U4762 ( .DIN1(n4528), .DIN2(n4529), .Q(n1321) );
  nnd2s1 U4763 ( .DIN1(text_in_r[102]), .DIN2(n1573), .Q(n4529) );
  nnd2s1 U4764 ( .DIN1(\text_in[102] ), .DIN2(ld), .Q(n4528) );
  nnd2s1 U4765 ( .DIN1(n4530), .DIN2(n4531), .Q(n1320) );
  nnd2s1 U4766 ( .DIN1(text_in_r[101]), .DIN2(n1573), .Q(n4531) );
  nnd2s1 U4767 ( .DIN1(\text_in[101] ), .DIN2(ld), .Q(n4530) );
  nnd2s1 U4768 ( .DIN1(n4532), .DIN2(n4533), .Q(n1319) );
  nnd2s1 U4769 ( .DIN1(text_in_r[100]), .DIN2(n1573), .Q(n4533) );
  nnd2s1 U4770 ( .DIN1(\text_in[100] ), .DIN2(ld), .Q(n4532) );
  nnd2s1 U4771 ( .DIN1(n4534), .DIN2(n4535), .Q(n1318) );
  nnd2s1 U4772 ( .DIN1(text_in_r[99]), .DIN2(n1574), .Q(n4535) );
  nnd2s1 U4773 ( .DIN1(\text_in[99] ), .DIN2(ld), .Q(n4534) );
  nnd2s1 U4774 ( .DIN1(n4536), .DIN2(n4537), .Q(n1317) );
  nnd2s1 U4775 ( .DIN1(text_in_r[98]), .DIN2(n1574), .Q(n4537) );
  nnd2s1 U4776 ( .DIN1(\text_in[98] ), .DIN2(ld), .Q(n4536) );
  nnd2s1 U4777 ( .DIN1(n4538), .DIN2(n4539), .Q(n1316) );
  nnd2s1 U4778 ( .DIN1(text_in_r[97]), .DIN2(n1574), .Q(n4539) );
  nnd2s1 U4779 ( .DIN1(\text_in[97] ), .DIN2(ld), .Q(n4538) );
  nnd2s1 U4780 ( .DIN1(n4540), .DIN2(n4541), .Q(n1315) );
  nnd2s1 U4781 ( .DIN1(text_in_r[96]), .DIN2(n1574), .Q(n4541) );
  nnd2s1 U4782 ( .DIN1(\text_in[96] ), .DIN2(ld), .Q(n4540) );
  nnd2s1 U4783 ( .DIN1(n4542), .DIN2(n4543), .Q(n1314) );
  nnd2s1 U4784 ( .DIN1(text_in_r[95]), .DIN2(n1574), .Q(n4543) );
  nnd2s1 U4785 ( .DIN1(\text_in[95] ), .DIN2(ld), .Q(n4542) );
  nnd2s1 U4786 ( .DIN1(n4544), .DIN2(n4545), .Q(n1313) );
  nnd2s1 U4787 ( .DIN1(text_in_r[94]), .DIN2(n1574), .Q(n4545) );
  nnd2s1 U4788 ( .DIN1(\text_in[94] ), .DIN2(ld), .Q(n4544) );
  nnd2s1 U4789 ( .DIN1(n4546), .DIN2(n4547), .Q(n1312) );
  nnd2s1 U4790 ( .DIN1(text_in_r[93]), .DIN2(n1575), .Q(n4547) );
  nnd2s1 U4791 ( .DIN1(\text_in[93] ), .DIN2(ld), .Q(n4546) );
  nnd2s1 U4792 ( .DIN1(n4548), .DIN2(n4549), .Q(n1311) );
  nnd2s1 U4793 ( .DIN1(text_in_r[92]), .DIN2(n1575), .Q(n4549) );
  nnd2s1 U4794 ( .DIN1(\text_in[92] ), .DIN2(ld), .Q(n4548) );
  nnd2s1 U4795 ( .DIN1(n4550), .DIN2(n4551), .Q(n1310) );
  nnd2s1 U4796 ( .DIN1(text_in_r[91]), .DIN2(n1575), .Q(n4551) );
  nnd2s1 U4797 ( .DIN1(\text_in[91] ), .DIN2(ld), .Q(n4550) );
  nnd2s1 U4798 ( .DIN1(n4552), .DIN2(n4553), .Q(n1309) );
  nnd2s1 U4799 ( .DIN1(text_in_r[90]), .DIN2(n1575), .Q(n4553) );
  nnd2s1 U4800 ( .DIN1(\text_in[90] ), .DIN2(ld), .Q(n4552) );
  nnd2s1 U4801 ( .DIN1(n4554), .DIN2(n4555), .Q(n1308) );
  nnd2s1 U4802 ( .DIN1(text_in_r[89]), .DIN2(n1575), .Q(n4555) );
  nnd2s1 U4803 ( .DIN1(\text_in[89] ), .DIN2(ld), .Q(n4554) );
  nnd2s1 U4804 ( .DIN1(n4556), .DIN2(n4557), .Q(n1307) );
  nnd2s1 U4805 ( .DIN1(text_in_r[88]), .DIN2(n1575), .Q(n4557) );
  nnd2s1 U4806 ( .DIN1(\text_in[88] ), .DIN2(ld), .Q(n4556) );
  nnd2s1 U4807 ( .DIN1(n4558), .DIN2(n4559), .Q(n1306) );
  nnd2s1 U4808 ( .DIN1(text_in_r[87]), .DIN2(n1575), .Q(n4559) );
  nnd2s1 U4809 ( .DIN1(\text_in[87] ), .DIN2(ld), .Q(n4558) );
  nnd2s1 U4810 ( .DIN1(n4560), .DIN2(n4561), .Q(n1305) );
  nnd2s1 U4811 ( .DIN1(text_in_r[86]), .DIN2(n1576), .Q(n4561) );
  nnd2s1 U4812 ( .DIN1(\text_in[86] ), .DIN2(ld), .Q(n4560) );
  nnd2s1 U4813 ( .DIN1(n4562), .DIN2(n4563), .Q(n1304) );
  nnd2s1 U4814 ( .DIN1(text_in_r[85]), .DIN2(n1576), .Q(n4563) );
  nnd2s1 U4815 ( .DIN1(\text_in[85] ), .DIN2(ld), .Q(n4562) );
  nnd2s1 U4816 ( .DIN1(n4564), .DIN2(n4565), .Q(n1303) );
  nnd2s1 U4817 ( .DIN1(text_in_r[84]), .DIN2(n1576), .Q(n4565) );
  nnd2s1 U4818 ( .DIN1(\text_in[84] ), .DIN2(ld), .Q(n4564) );
  nnd2s1 U4819 ( .DIN1(n4566), .DIN2(n4567), .Q(n1302) );
  nnd2s1 U4820 ( .DIN1(text_in_r[83]), .DIN2(n1576), .Q(n4567) );
  nnd2s1 U4821 ( .DIN1(\text_in[83] ), .DIN2(ld), .Q(n4566) );
  nnd2s1 U4822 ( .DIN1(n4568), .DIN2(n4569), .Q(n1301) );
  nnd2s1 U4823 ( .DIN1(text_in_r[82]), .DIN2(n1576), .Q(n4569) );
  nnd2s1 U4824 ( .DIN1(\text_in[82] ), .DIN2(ld), .Q(n4568) );
  nnd2s1 U4825 ( .DIN1(n4570), .DIN2(n4571), .Q(n1300) );
  nnd2s1 U4826 ( .DIN1(text_in_r[81]), .DIN2(n1576), .Q(n4571) );
  nnd2s1 U4827 ( .DIN1(\text_in[81] ), .DIN2(ld), .Q(n4570) );
  nnd2s1 U4828 ( .DIN1(n4572), .DIN2(n4573), .Q(n1299) );
  nnd2s1 U4829 ( .DIN1(text_in_r[80]), .DIN2(n1576), .Q(n4573) );
  nnd2s1 U4830 ( .DIN1(\text_in[80] ), .DIN2(ld), .Q(n4572) );
  nnd2s1 U4831 ( .DIN1(n4574), .DIN2(n4575), .Q(n1298) );
  nnd2s1 U4832 ( .DIN1(text_in_r[79]), .DIN2(n1577), .Q(n4575) );
  nnd2s1 U4833 ( .DIN1(\text_in[79] ), .DIN2(ld), .Q(n4574) );
  nnd2s1 U4834 ( .DIN1(n4576), .DIN2(n4577), .Q(n1297) );
  nnd2s1 U4835 ( .DIN1(text_in_r[78]), .DIN2(n1577), .Q(n4577) );
  nnd2s1 U4836 ( .DIN1(\text_in[78] ), .DIN2(ld), .Q(n4576) );
  nnd2s1 U4837 ( .DIN1(n4578), .DIN2(n4579), .Q(n1296) );
  nnd2s1 U4838 ( .DIN1(text_in_r[77]), .DIN2(n1577), .Q(n4579) );
  nnd2s1 U4839 ( .DIN1(\text_in[77] ), .DIN2(ld), .Q(n4578) );
  nnd2s1 U4840 ( .DIN1(n4580), .DIN2(n4581), .Q(n1295) );
  nnd2s1 U4841 ( .DIN1(text_in_r[76]), .DIN2(n1577), .Q(n4581) );
  nnd2s1 U4842 ( .DIN1(\text_in[76] ), .DIN2(ld), .Q(n4580) );
  nnd2s1 U4843 ( .DIN1(n4582), .DIN2(n4583), .Q(n1294) );
  nnd2s1 U4844 ( .DIN1(text_in_r[75]), .DIN2(n1577), .Q(n4583) );
  nnd2s1 U4845 ( .DIN1(\text_in[75] ), .DIN2(ld), .Q(n4582) );
  nnd2s1 U4846 ( .DIN1(n4584), .DIN2(n4585), .Q(n1293) );
  nnd2s1 U4847 ( .DIN1(text_in_r[74]), .DIN2(n1577), .Q(n4585) );
  nnd2s1 U4848 ( .DIN1(\text_in[74] ), .DIN2(ld), .Q(n4584) );
  nnd2s1 U4849 ( .DIN1(n4586), .DIN2(n4587), .Q(n1292) );
  nnd2s1 U4850 ( .DIN1(text_in_r[73]), .DIN2(n1577), .Q(n4587) );
  nnd2s1 U4851 ( .DIN1(\text_in[73] ), .DIN2(ld), .Q(n4586) );
  nnd2s1 U4852 ( .DIN1(n4588), .DIN2(n4589), .Q(n1291) );
  nnd2s1 U4853 ( .DIN1(text_in_r[72]), .DIN2(n1578), .Q(n4589) );
  nnd2s1 U4854 ( .DIN1(\text_in[72] ), .DIN2(ld), .Q(n4588) );
  nnd2s1 U4855 ( .DIN1(n4590), .DIN2(n4591), .Q(n1290) );
  nnd2s1 U4856 ( .DIN1(text_in_r[71]), .DIN2(n1578), .Q(n4591) );
  nnd2s1 U4857 ( .DIN1(\text_in[71] ), .DIN2(ld), .Q(n4590) );
  nnd2s1 U4858 ( .DIN1(n4592), .DIN2(n4593), .Q(n1289) );
  nnd2s1 U4859 ( .DIN1(text_in_r[70]), .DIN2(n1578), .Q(n4593) );
  nnd2s1 U4860 ( .DIN1(\text_in[70] ), .DIN2(ld), .Q(n4592) );
  nnd2s1 U4861 ( .DIN1(n4594), .DIN2(n4595), .Q(n1288) );
  nnd2s1 U4862 ( .DIN1(text_in_r[69]), .DIN2(n1578), .Q(n4595) );
  nnd2s1 U4863 ( .DIN1(\text_in[69] ), .DIN2(ld), .Q(n4594) );
  nnd2s1 U4864 ( .DIN1(n4596), .DIN2(n4597), .Q(n1287) );
  nnd2s1 U4865 ( .DIN1(text_in_r[68]), .DIN2(n1578), .Q(n4597) );
  nnd2s1 U4866 ( .DIN1(\text_in[68] ), .DIN2(ld), .Q(n4596) );
  nnd2s1 U4867 ( .DIN1(n4598), .DIN2(n4599), .Q(n1286) );
  nnd2s1 U4868 ( .DIN1(text_in_r[67]), .DIN2(n1578), .Q(n4599) );
  nnd2s1 U4869 ( .DIN1(\text_in[67] ), .DIN2(ld), .Q(n4598) );
  nnd2s1 U4870 ( .DIN1(n4600), .DIN2(n4601), .Q(n1285) );
  nnd2s1 U4871 ( .DIN1(text_in_r[66]), .DIN2(n1578), .Q(n4601) );
  nnd2s1 U4872 ( .DIN1(\text_in[66] ), .DIN2(ld), .Q(n4600) );
  nnd2s1 U4873 ( .DIN1(n4602), .DIN2(n4603), .Q(n1284) );
  nnd2s1 U4874 ( .DIN1(text_in_r[65]), .DIN2(n1579), .Q(n4603) );
  nnd2s1 U4875 ( .DIN1(\text_in[65] ), .DIN2(ld), .Q(n4602) );
  nnd2s1 U4876 ( .DIN1(n4604), .DIN2(n4605), .Q(n1283) );
  nnd2s1 U4877 ( .DIN1(text_in_r[64]), .DIN2(n1579), .Q(n4605) );
  nnd2s1 U4878 ( .DIN1(\text_in[64] ), .DIN2(ld), .Q(n4604) );
  nnd2s1 U4879 ( .DIN1(n4606), .DIN2(n4607), .Q(n1282) );
  nnd2s1 U4880 ( .DIN1(text_in_r[63]), .DIN2(n1579), .Q(n4607) );
  nnd2s1 U4881 ( .DIN1(\text_in[63] ), .DIN2(ld), .Q(n4606) );
  nnd2s1 U4882 ( .DIN1(n4608), .DIN2(n4609), .Q(n1281) );
  nnd2s1 U4883 ( .DIN1(text_in_r[62]), .DIN2(n1579), .Q(n4609) );
  nnd2s1 U4884 ( .DIN1(\text_in[62] ), .DIN2(ld), .Q(n4608) );
  nnd2s1 U4885 ( .DIN1(n4610), .DIN2(n4611), .Q(n1280) );
  nnd2s1 U4886 ( .DIN1(text_in_r[61]), .DIN2(n1579), .Q(n4611) );
  nnd2s1 U4887 ( .DIN1(\text_in[61] ), .DIN2(ld), .Q(n4610) );
  nnd2s1 U4888 ( .DIN1(n4612), .DIN2(n4613), .Q(n1279) );
  nnd2s1 U4889 ( .DIN1(text_in_r[60]), .DIN2(n1579), .Q(n4613) );
  nnd2s1 U4890 ( .DIN1(\text_in[60] ), .DIN2(ld), .Q(n4612) );
  nnd2s1 U4891 ( .DIN1(n4614), .DIN2(n4615), .Q(n1278) );
  nnd2s1 U4892 ( .DIN1(text_in_r[59]), .DIN2(n1579), .Q(n4615) );
  nnd2s1 U4893 ( .DIN1(\text_in[59] ), .DIN2(ld), .Q(n4614) );
  nnd2s1 U4894 ( .DIN1(n4616), .DIN2(n4617), .Q(n1277) );
  nnd2s1 U4895 ( .DIN1(text_in_r[58]), .DIN2(n1580), .Q(n4617) );
  nnd2s1 U4896 ( .DIN1(\text_in[58] ), .DIN2(ld), .Q(n4616) );
  nnd2s1 U4897 ( .DIN1(n4618), .DIN2(n4619), .Q(n1276) );
  nnd2s1 U4898 ( .DIN1(text_in_r[57]), .DIN2(n1580), .Q(n4619) );
  nnd2s1 U4899 ( .DIN1(\text_in[57] ), .DIN2(ld), .Q(n4618) );
  nnd2s1 U4900 ( .DIN1(n4620), .DIN2(n4621), .Q(n1275) );
  nnd2s1 U4901 ( .DIN1(text_in_r[56]), .DIN2(n1580), .Q(n4621) );
  nnd2s1 U4902 ( .DIN1(\text_in[56] ), .DIN2(ld), .Q(n4620) );
  nnd2s1 U4903 ( .DIN1(n4622), .DIN2(n4623), .Q(n1274) );
  nnd2s1 U4904 ( .DIN1(text_in_r[55]), .DIN2(n1580), .Q(n4623) );
  nnd2s1 U4905 ( .DIN1(\text_in[55] ), .DIN2(ld), .Q(n4622) );
  nnd2s1 U4906 ( .DIN1(n4624), .DIN2(n4625), .Q(n1273) );
  nnd2s1 U4907 ( .DIN1(text_in_r[54]), .DIN2(n1580), .Q(n4625) );
  nnd2s1 U4908 ( .DIN1(\text_in[54] ), .DIN2(ld), .Q(n4624) );
  nnd2s1 U4909 ( .DIN1(n4626), .DIN2(n4627), .Q(n1272) );
  nnd2s1 U4910 ( .DIN1(text_in_r[53]), .DIN2(n1580), .Q(n4627) );
  nnd2s1 U4911 ( .DIN1(\text_in[53] ), .DIN2(ld), .Q(n4626) );
  nnd2s1 U4912 ( .DIN1(n4628), .DIN2(n4629), .Q(n1271) );
  nnd2s1 U4913 ( .DIN1(text_in_r[52]), .DIN2(n1580), .Q(n4629) );
  nnd2s1 U4914 ( .DIN1(\text_in[52] ), .DIN2(ld), .Q(n4628) );
  nnd2s1 U4915 ( .DIN1(n4630), .DIN2(n4631), .Q(n1270) );
  nnd2s1 U4916 ( .DIN1(text_in_r[51]), .DIN2(n1581), .Q(n4631) );
  nnd2s1 U4917 ( .DIN1(\text_in[51] ), .DIN2(ld), .Q(n4630) );
  nnd2s1 U4918 ( .DIN1(n4632), .DIN2(n4633), .Q(n1269) );
  nnd2s1 U4919 ( .DIN1(text_in_r[50]), .DIN2(n1581), .Q(n4633) );
  nnd2s1 U4920 ( .DIN1(\text_in[50] ), .DIN2(ld), .Q(n4632) );
  nnd2s1 U4921 ( .DIN1(n4634), .DIN2(n4635), .Q(n1268) );
  nnd2s1 U4922 ( .DIN1(text_in_r[49]), .DIN2(n1581), .Q(n4635) );
  nnd2s1 U4923 ( .DIN1(\text_in[49] ), .DIN2(ld), .Q(n4634) );
  nnd2s1 U4924 ( .DIN1(n4636), .DIN2(n4637), .Q(n1267) );
  nnd2s1 U4925 ( .DIN1(text_in_r[48]), .DIN2(n1581), .Q(n4637) );
  nnd2s1 U4926 ( .DIN1(\text_in[48] ), .DIN2(ld), .Q(n4636) );
  nnd2s1 U4927 ( .DIN1(n4638), .DIN2(n4639), .Q(n1266) );
  nnd2s1 U4928 ( .DIN1(text_in_r[47]), .DIN2(n1581), .Q(n4639) );
  nnd2s1 U4929 ( .DIN1(\text_in[47] ), .DIN2(ld), .Q(n4638) );
  nnd2s1 U4930 ( .DIN1(n4640), .DIN2(n4641), .Q(n1265) );
  nnd2s1 U4931 ( .DIN1(text_in_r[46]), .DIN2(n1581), .Q(n4641) );
  nnd2s1 U4932 ( .DIN1(\text_in[46] ), .DIN2(ld), .Q(n4640) );
  nnd2s1 U4933 ( .DIN1(n4642), .DIN2(n4643), .Q(n1264) );
  nnd2s1 U4934 ( .DIN1(text_in_r[45]), .DIN2(n1581), .Q(n4643) );
  nnd2s1 U4935 ( .DIN1(\text_in[45] ), .DIN2(ld), .Q(n4642) );
  nnd2s1 U4936 ( .DIN1(n4644), .DIN2(n4645), .Q(n1263) );
  nnd2s1 U4937 ( .DIN1(text_in_r[44]), .DIN2(n1582), .Q(n4645) );
  nnd2s1 U4938 ( .DIN1(\text_in[44] ), .DIN2(ld), .Q(n4644) );
  nnd2s1 U4939 ( .DIN1(n4646), .DIN2(n4647), .Q(n1262) );
  nnd2s1 U4940 ( .DIN1(text_in_r[43]), .DIN2(n1582), .Q(n4647) );
  nnd2s1 U4941 ( .DIN1(\text_in[43] ), .DIN2(ld), .Q(n4646) );
  nnd2s1 U4942 ( .DIN1(n4648), .DIN2(n4649), .Q(n1261) );
  nnd2s1 U4943 ( .DIN1(text_in_r[42]), .DIN2(n1582), .Q(n4649) );
  nnd2s1 U4944 ( .DIN1(\text_in[42] ), .DIN2(ld), .Q(n4648) );
  nnd2s1 U4945 ( .DIN1(n4650), .DIN2(n4651), .Q(n1260) );
  nnd2s1 U4946 ( .DIN1(text_in_r[41]), .DIN2(n1582), .Q(n4651) );
  nnd2s1 U4947 ( .DIN1(\text_in[41] ), .DIN2(ld), .Q(n4650) );
  nnd2s1 U4948 ( .DIN1(n4652), .DIN2(n4653), .Q(n1259) );
  nnd2s1 U4949 ( .DIN1(text_in_r[40]), .DIN2(n1582), .Q(n4653) );
  nnd2s1 U4950 ( .DIN1(\text_in[40] ), .DIN2(ld), .Q(n4652) );
  nnd2s1 U4951 ( .DIN1(n4654), .DIN2(n4655), .Q(n1258) );
  nnd2s1 U4952 ( .DIN1(text_in_r[39]), .DIN2(n1582), .Q(n4655) );
  nnd2s1 U4953 ( .DIN1(\text_in[39] ), .DIN2(ld), .Q(n4654) );
  nnd2s1 U4954 ( .DIN1(n4656), .DIN2(n4657), .Q(n1257) );
  nnd2s1 U4955 ( .DIN1(text_in_r[38]), .DIN2(n1582), .Q(n4657) );
  nnd2s1 U4956 ( .DIN1(\text_in[38] ), .DIN2(ld), .Q(n4656) );
  nnd2s1 U4957 ( .DIN1(n4658), .DIN2(n4659), .Q(n1256) );
  nnd2s1 U4958 ( .DIN1(text_in_r[37]), .DIN2(n1583), .Q(n4659) );
  nnd2s1 U4959 ( .DIN1(\text_in[37] ), .DIN2(ld), .Q(n4658) );
  nnd2s1 U4960 ( .DIN1(n4660), .DIN2(n4661), .Q(n1255) );
  nnd2s1 U4961 ( .DIN1(text_in_r[36]), .DIN2(n1583), .Q(n4661) );
  nnd2s1 U4962 ( .DIN1(\text_in[36] ), .DIN2(ld), .Q(n4660) );
  nnd2s1 U4963 ( .DIN1(n4662), .DIN2(n4663), .Q(n1254) );
  nnd2s1 U4964 ( .DIN1(text_in_r[35]), .DIN2(n1583), .Q(n4663) );
  nnd2s1 U4965 ( .DIN1(\text_in[35] ), .DIN2(ld), .Q(n4662) );
  nnd2s1 U4966 ( .DIN1(n4664), .DIN2(n4665), .Q(n1253) );
  nnd2s1 U4967 ( .DIN1(text_in_r[34]), .DIN2(n1583), .Q(n4665) );
  nnd2s1 U4968 ( .DIN1(\text_in[34] ), .DIN2(ld), .Q(n4664) );
  nnd2s1 U4969 ( .DIN1(n4666), .DIN2(n4667), .Q(n1252) );
  nnd2s1 U4970 ( .DIN1(text_in_r[33]), .DIN2(n1583), .Q(n4667) );
  nnd2s1 U4971 ( .DIN1(\text_in[33] ), .DIN2(ld), .Q(n4666) );
  nnd2s1 U4972 ( .DIN1(n4668), .DIN2(n4669), .Q(n1251) );
  nnd2s1 U4973 ( .DIN1(text_in_r[32]), .DIN2(n1583), .Q(n4669) );
  nnd2s1 U4974 ( .DIN1(\text_in[32] ), .DIN2(ld), .Q(n4668) );
  nnd2s1 U4975 ( .DIN1(n4670), .DIN2(n4671), .Q(n1250) );
  nnd2s1 U4976 ( .DIN1(text_in_r[31]), .DIN2(n1583), .Q(n4671) );
  nnd2s1 U4977 ( .DIN1(\text_in[31] ), .DIN2(ld), .Q(n4670) );
  nnd2s1 U4978 ( .DIN1(n4672), .DIN2(n4673), .Q(n1249) );
  nnd2s1 U4979 ( .DIN1(text_in_r[30]), .DIN2(n1584), .Q(n4673) );
  nnd2s1 U4980 ( .DIN1(\text_in[30] ), .DIN2(ld), .Q(n4672) );
  nnd2s1 U4981 ( .DIN1(n4674), .DIN2(n4675), .Q(n1248) );
  nnd2s1 U4982 ( .DIN1(text_in_r[29]), .DIN2(n1584), .Q(n4675) );
  nnd2s1 U4983 ( .DIN1(\text_in[29] ), .DIN2(ld), .Q(n4674) );
  nnd2s1 U4984 ( .DIN1(n4676), .DIN2(n4677), .Q(n1247) );
  nnd2s1 U4985 ( .DIN1(text_in_r[28]), .DIN2(n1584), .Q(n4677) );
  nnd2s1 U4986 ( .DIN1(\text_in[28] ), .DIN2(ld), .Q(n4676) );
  nnd2s1 U4987 ( .DIN1(n4678), .DIN2(n4679), .Q(n1246) );
  nnd2s1 U4988 ( .DIN1(text_in_r[27]), .DIN2(n1584), .Q(n4679) );
  nnd2s1 U4989 ( .DIN1(\text_in[27] ), .DIN2(ld), .Q(n4678) );
  nnd2s1 U4990 ( .DIN1(n4680), .DIN2(n4681), .Q(n1245) );
  nnd2s1 U4991 ( .DIN1(text_in_r[26]), .DIN2(n1584), .Q(n4681) );
  nnd2s1 U4992 ( .DIN1(\text_in[26] ), .DIN2(ld), .Q(n4680) );
  nnd2s1 U4993 ( .DIN1(n4682), .DIN2(n4683), .Q(n1244) );
  nnd2s1 U4994 ( .DIN1(text_in_r[25]), .DIN2(n1584), .Q(n4683) );
  nnd2s1 U4995 ( .DIN1(\text_in[25] ), .DIN2(ld), .Q(n4682) );
  nnd2s1 U4996 ( .DIN1(n4684), .DIN2(n4685), .Q(n1243) );
  nnd2s1 U4997 ( .DIN1(text_in_r[24]), .DIN2(n1584), .Q(n4685) );
  nnd2s1 U4998 ( .DIN1(\text_in[24] ), .DIN2(ld), .Q(n4684) );
  nnd2s1 U4999 ( .DIN1(n4686), .DIN2(n4687), .Q(n1242) );
  nnd2s1 U5000 ( .DIN1(text_in_r[23]), .DIN2(n1585), .Q(n4687) );
  nnd2s1 U5001 ( .DIN1(\text_in[23] ), .DIN2(ld), .Q(n4686) );
  nnd2s1 U5002 ( .DIN1(n4688), .DIN2(n4689), .Q(n1241) );
  nnd2s1 U5003 ( .DIN1(text_in_r[22]), .DIN2(n1585), .Q(n4689) );
  nnd2s1 U5004 ( .DIN1(\text_in[22] ), .DIN2(ld), .Q(n4688) );
  nnd2s1 U5005 ( .DIN1(n4690), .DIN2(n4691), .Q(n1240) );
  nnd2s1 U5006 ( .DIN1(text_in_r[21]), .DIN2(n1585), .Q(n4691) );
  nnd2s1 U5007 ( .DIN1(\text_in[21] ), .DIN2(ld), .Q(n4690) );
  nnd2s1 U5008 ( .DIN1(n4692), .DIN2(n4693), .Q(n1239) );
  nnd2s1 U5009 ( .DIN1(text_in_r[20]), .DIN2(n1585), .Q(n4693) );
  nnd2s1 U5010 ( .DIN1(\text_in[20] ), .DIN2(ld), .Q(n4692) );
  nnd2s1 U5011 ( .DIN1(n4694), .DIN2(n4695), .Q(n1238) );
  nnd2s1 U5012 ( .DIN1(text_in_r[19]), .DIN2(n1585), .Q(n4695) );
  nnd2s1 U5013 ( .DIN1(\text_in[19] ), .DIN2(ld), .Q(n4694) );
  nnd2s1 U5014 ( .DIN1(n4696), .DIN2(n4697), .Q(n1237) );
  nnd2s1 U5015 ( .DIN1(text_in_r[18]), .DIN2(n1585), .Q(n4697) );
  nnd2s1 U5016 ( .DIN1(\text_in[18] ), .DIN2(ld), .Q(n4696) );
  nnd2s1 U5017 ( .DIN1(n4698), .DIN2(n4699), .Q(n1236) );
  nnd2s1 U5018 ( .DIN1(text_in_r[17]), .DIN2(n1585), .Q(n4699) );
  nnd2s1 U5019 ( .DIN1(\text_in[17] ), .DIN2(ld), .Q(n4698) );
  nnd2s1 U5020 ( .DIN1(n4700), .DIN2(n4701), .Q(n1235) );
  nnd2s1 U5021 ( .DIN1(text_in_r[16]), .DIN2(n1586), .Q(n4701) );
  nnd2s1 U5022 ( .DIN1(\text_in[16] ), .DIN2(ld), .Q(n4700) );
  nnd2s1 U5023 ( .DIN1(n4702), .DIN2(n4703), .Q(n1234) );
  nnd2s1 U5024 ( .DIN1(text_in_r[15]), .DIN2(n1586), .Q(n4703) );
  nnd2s1 U5025 ( .DIN1(\text_in[15] ), .DIN2(ld), .Q(n4702) );
  nnd2s1 U5026 ( .DIN1(n4704), .DIN2(n4705), .Q(n1233) );
  nnd2s1 U5027 ( .DIN1(text_in_r[14]), .DIN2(n1586), .Q(n4705) );
  nnd2s1 U5028 ( .DIN1(\text_in[14] ), .DIN2(ld), .Q(n4704) );
  nnd2s1 U5029 ( .DIN1(n4706), .DIN2(n4707), .Q(n1232) );
  nnd2s1 U5030 ( .DIN1(text_in_r[13]), .DIN2(n1586), .Q(n4707) );
  nnd2s1 U5031 ( .DIN1(\text_in[13] ), .DIN2(ld), .Q(n4706) );
  nnd2s1 U5032 ( .DIN1(n4708), .DIN2(n4709), .Q(n1231) );
  nnd2s1 U5033 ( .DIN1(text_in_r[12]), .DIN2(n1586), .Q(n4709) );
  nnd2s1 U5034 ( .DIN1(\text_in[12] ), .DIN2(ld), .Q(n4708) );
  nnd2s1 U5035 ( .DIN1(n4710), .DIN2(n4711), .Q(n1230) );
  nnd2s1 U5036 ( .DIN1(text_in_r[11]), .DIN2(n1586), .Q(n4711) );
  nnd2s1 U5037 ( .DIN1(\text_in[11] ), .DIN2(ld), .Q(n4710) );
  nnd2s1 U5038 ( .DIN1(n4712), .DIN2(n4713), .Q(n1229) );
  nnd2s1 U5039 ( .DIN1(text_in_r[10]), .DIN2(n1586), .Q(n4713) );
  nnd2s1 U5040 ( .DIN1(\text_in[10] ), .DIN2(ld), .Q(n4712) );
  nnd2s1 U5041 ( .DIN1(n4714), .DIN2(n4715), .Q(n1228) );
  nnd2s1 U5042 ( .DIN1(text_in_r[9]), .DIN2(n1587), .Q(n4715) );
  nnd2s1 U5043 ( .DIN1(\text_in[9] ), .DIN2(ld), .Q(n4714) );
  nnd2s1 U5044 ( .DIN1(n4716), .DIN2(n4717), .Q(n1227) );
  nnd2s1 U5045 ( .DIN1(text_in_r[8]), .DIN2(n1587), .Q(n4717) );
  nnd2s1 U5046 ( .DIN1(\text_in[8] ), .DIN2(ld), .Q(n4716) );
  nnd2s1 U5047 ( .DIN1(n4718), .DIN2(n4719), .Q(n1226) );
  nnd2s1 U5048 ( .DIN1(text_in_r[7]), .DIN2(n1587), .Q(n4719) );
  nnd2s1 U5049 ( .DIN1(\text_in[7] ), .DIN2(ld), .Q(n4718) );
  nnd2s1 U5050 ( .DIN1(n4720), .DIN2(n4721), .Q(n1225) );
  nnd2s1 U5051 ( .DIN1(text_in_r[6]), .DIN2(n1587), .Q(n4721) );
  nnd2s1 U5052 ( .DIN1(\text_in[6] ), .DIN2(ld), .Q(n4720) );
  nnd2s1 U5053 ( .DIN1(n4722), .DIN2(n4723), .Q(n1224) );
  nnd2s1 U5054 ( .DIN1(text_in_r[5]), .DIN2(n1587), .Q(n4723) );
  nnd2s1 U5055 ( .DIN1(\text_in[5] ), .DIN2(ld), .Q(n4722) );
  nnd2s1 U5056 ( .DIN1(n4724), .DIN2(n4725), .Q(n1223) );
  nnd2s1 U5057 ( .DIN1(text_in_r[4]), .DIN2(n1587), .Q(n4725) );
  nnd2s1 U5058 ( .DIN1(\text_in[4] ), .DIN2(ld), .Q(n4724) );
  nnd2s1 U5059 ( .DIN1(n4726), .DIN2(n4727), .Q(n1222) );
  nnd2s1 U5060 ( .DIN1(text_in_r[3]), .DIN2(n1587), .Q(n4727) );
  nnd2s1 U5061 ( .DIN1(\text_in[3] ), .DIN2(ld), .Q(n4726) );
  nnd2s1 U5062 ( .DIN1(n4728), .DIN2(n4729), .Q(n1221) );
  nnd2s1 U5063 ( .DIN1(text_in_r[2]), .DIN2(n1592), .Q(n4729) );
  nnd2s1 U5064 ( .DIN1(\text_in[2] ), .DIN2(ld), .Q(n4728) );
  nnd2s1 U5065 ( .DIN1(n4730), .DIN2(n4731), .Q(n1220) );
  nnd2s1 U5066 ( .DIN1(text_in_r[1]), .DIN2(n1588), .Q(n4731) );
  nnd2s1 U5067 ( .DIN1(\text_in[1] ), .DIN2(ld), .Q(n4730) );
  nnd2s1 U5068 ( .DIN1(n4732), .DIN2(n4733), .Q(n1219) );
  nnd2s1 U5069 ( .DIN1(text_in_r[0]), .DIN2(n1560), .Q(n4733) );
  hi1s1 U5070 ( .DIN(ld), .Q(n1669) );
  nnd2s1 U5071 ( .DIN1(\text_in[0] ), .DIN2(ld), .Q(n4732) );
  nnd2s1 U5072 ( .DIN1(n4734), .DIN2(n4735), .Q(N99) );
  nnd2s1 U5073 ( .DIN1(n4736), .DIN2(n1630), .Q(n4735) );
  xor2s1 U5074 ( .DIN1(n4737), .DIN2(n4738), .Q(n4736) );
  xor2s1 U5075 ( .DIN1(n4739), .DIN2(n4740), .Q(n4738) );
  xnr2s1 U5076 ( .DIN1(n4742), .DIN2(n4741), .Q(n4740) );
  xor2s1 U5077 ( .DIN1(n4743), .DIN2(n4744), .Q(n4737) );
  xor2s1 U5078 ( .DIN1(n1479), .DIN2(n4745), .Q(n4743) );
  nnd2s1 U5079 ( .DIN1(n4746), .DIN2(n1599), .Q(n4734) );
  xor2s1 U5080 ( .DIN1(w2[1]), .DIN2(text_in_r[33]), .Q(n4746) );
  nnd2s1 U5081 ( .DIN1(n4747), .DIN2(n4748), .Q(N98) );
  nnd2s1 U5082 ( .DIN1(n4749), .DIN2(n1608), .Q(n4748) );
  xor2s1 U5083 ( .DIN1(n4750), .DIN2(n4751), .Q(n4749) );
  xor2s1 U5084 ( .DIN1(n4752), .DIN2(n4753), .Q(n4751) );
  xor2s1 U5085 ( .DIN1(n1450), .DIN2(n4754), .Q(n4750) );
  nnd2s1 U5086 ( .DIN1(n4755), .DIN2(n1607), .Q(n4747) );
  xor2s1 U5087 ( .DIN1(w2[0]), .DIN2(text_in_r[32]), .Q(n4755) );
  nnd2s1 U5088 ( .DIN1(n4756), .DIN2(n4757), .Q(N89) );
  nnd2s1 U5089 ( .DIN1(n4758), .DIN2(n1608), .Q(n4757) );
  xor2s1 U5090 ( .DIN1(n4759), .DIN2(n4760), .Q(n4758) );
  xor2s1 U5091 ( .DIN1(n4761), .DIN2(n4762), .Q(n4760) );
  xor2s1 U5092 ( .DIN1(n1416), .DIN2(n4763), .Q(n4759) );
  nnd2s1 U5093 ( .DIN1(n4764), .DIN2(n1607), .Q(n4756) );
  xor2s1 U5094 ( .DIN1(w3[31]), .DIN2(text_in_r[31]), .Q(n4764) );
  nnd2s1 U5095 ( .DIN1(n4765), .DIN2(n4766), .Q(N88) );
  nnd2s1 U5096 ( .DIN1(n4767), .DIN2(n1608), .Q(n4766) );
  xor2s1 U5097 ( .DIN1(n4768), .DIN2(n4769), .Q(n4767) );
  xor2s1 U5098 ( .DIN1(n4770), .DIN2(n4771), .Q(n4769) );
  xor2s1 U5099 ( .DIN1(n4772), .DIN2(w3[30]), .Q(n4768) );
  nnd2s1 U5100 ( .DIN1(n4773), .DIN2(n1607), .Q(n4765) );
  xor2s1 U5101 ( .DIN1(w3[30]), .DIN2(text_in_r[30]), .Q(n4773) );
  nnd2s1 U5102 ( .DIN1(n4774), .DIN2(n4775), .Q(N87) );
  nnd2s1 U5103 ( .DIN1(n4776), .DIN2(n1609), .Q(n4775) );
  xor2s1 U5104 ( .DIN1(n4777), .DIN2(n4778), .Q(n4776) );
  xor2s1 U5105 ( .DIN1(n4779), .DIN2(n4780), .Q(n4778) );
  xor2s1 U5106 ( .DIN1(n1374), .DIN2(n4781), .Q(n4777) );
  nnd2s1 U5107 ( .DIN1(n4782), .DIN2(n1607), .Q(n4774) );
  xor2s1 U5108 ( .DIN1(w3[29]), .DIN2(text_in_r[29]), .Q(n4782) );
  nnd3s1 U5109 ( .DIN1(n4783), .DIN2(n4784), .DIN3(n4785), .Q(N86) );
  nnd2s1 U5110 ( .DIN1(n1597), .DIN2(n4786), .Q(n4785) );
  xor2s1 U5111 ( .DIN1(w3[28]), .DIN2(text_in_r[28]), .Q(n4786) );
  nnd2s1 U5112 ( .DIN1(n4787), .DIN2(n4788), .Q(n4784) );
  nnd2s1 U5113 ( .DIN1(n4789), .DIN2(n4790), .Q(n4787) );
  nnd2s1 U5114 ( .DIN1(n4791), .DIN2(n4792), .Q(n4790) );
  nnd2s1 U5115 ( .DIN1(n4793), .DIN2(n4794), .Q(n4789) );
  nnd2s1 U5116 ( .DIN1(n4795), .DIN2(n4796), .Q(n4783) );
  nnd2s1 U5117 ( .DIN1(n4797), .DIN2(n4798), .Q(n4796) );
  nnd2s1 U5118 ( .DIN1(n4793), .DIN2(n4792), .Q(n4798) );
  nnd2s1 U5119 ( .DIN1(n4794), .DIN2(n4791), .Q(n4797) );
  hi1s1 U5120 ( .DIN(n4792), .Q(n4794) );
  xor2s1 U5121 ( .DIN1(n4799), .DIN2(n4800), .Q(n4792) );
  xor2s1 U5122 ( .DIN1(n1392), .DIN2(n4801), .Q(n4799) );
  nnd3s1 U5123 ( .DIN1(n4802), .DIN2(n4803), .DIN3(n4804), .Q(N85) );
  nnd2s1 U5124 ( .DIN1(n1596), .DIN2(n4805), .Q(n4804) );
  xor2s1 U5125 ( .DIN1(w3[27]), .DIN2(text_in_r[27]), .Q(n4805) );
  nnd2s1 U5126 ( .DIN1(n4806), .DIN2(n4807), .Q(n4803) );
  nnd2s1 U5127 ( .DIN1(n4808), .DIN2(n4809), .Q(n4806) );
  nnd2s1 U5128 ( .DIN1(n4810), .DIN2(n4811), .Q(n4809) );
  nnd2s1 U5129 ( .DIN1(n4812), .DIN2(n4813), .Q(n4808) );
  nnd2s1 U5130 ( .DIN1(n4814), .DIN2(n4815), .Q(n4802) );
  nnd2s1 U5131 ( .DIN1(n4816), .DIN2(n4817), .Q(n4815) );
  nnd2s1 U5132 ( .DIN1(n4812), .DIN2(n4811), .Q(n4817) );
  nnd2s1 U5133 ( .DIN1(n4813), .DIN2(n4810), .Q(n4816) );
  hi1s1 U5134 ( .DIN(n4811), .Q(n4813) );
  xor2s1 U5135 ( .DIN1(n4818), .DIN2(n4795), .Q(n4811) );
  xor2s1 U5136 ( .DIN1(n4819), .DIN2(w3[27]), .Q(n4818) );
  nnd2s1 U5137 ( .DIN1(n4820), .DIN2(n4821), .Q(N84) );
  nnd2s1 U5138 ( .DIN1(n4822), .DIN2(n1609), .Q(n4821) );
  xor2s1 U5139 ( .DIN1(n4823), .DIN2(n4824), .Q(n4822) );
  xor2s1 U5140 ( .DIN1(n4825), .DIN2(n1552), .Q(n4824) );
  xor2s1 U5141 ( .DIN1(n4827), .DIN2(w3[26]), .Q(n4823) );
  nnd2s1 U5142 ( .DIN1(n4828), .DIN2(n1606), .Q(n4820) );
  xor2s1 U5143 ( .DIN1(w3[26]), .DIN2(text_in_r[26]), .Q(n4828) );
  nnd2s1 U5144 ( .DIN1(n4829), .DIN2(n4830), .Q(N83) );
  nnd2s1 U5145 ( .DIN1(n4831), .DIN2(n1609), .Q(n4830) );
  xor2s1 U5146 ( .DIN1(n4832), .DIN2(n4833), .Q(n4831) );
  xor2s1 U5147 ( .DIN1(n1546), .DIN2(n4835), .Q(n4833) );
  xor2s1 U5148 ( .DIN1(n4836), .DIN2(n4795), .Q(n4832) );
  xor2s1 U5149 ( .DIN1(n1410), .DIN2(n4837), .Q(n4836) );
  nnd2s1 U5150 ( .DIN1(n4838), .DIN2(n1606), .Q(n4829) );
  xor2s1 U5151 ( .DIN1(w3[25]), .DIN2(text_in_r[25]), .Q(n4838) );
  nnd2s1 U5152 ( .DIN1(n4839), .DIN2(n4840), .Q(N82) );
  nnd2s1 U5153 ( .DIN1(n4841), .DIN2(n1610), .Q(n4840) );
  xor2s1 U5154 ( .DIN1(n4842), .DIN2(n4843), .Q(n4841) );
  xor2s1 U5155 ( .DIN1(n4795), .DIN2(n4844), .Q(n4843) );
  xor2s1 U5156 ( .DIN1(n1554), .DIN2(n4845), .Q(n4842) );
  nnd2s1 U5157 ( .DIN1(n4846), .DIN2(n1606), .Q(n4839) );
  xor2s1 U5158 ( .DIN1(n1555), .DIN2(text_in_r[24]), .Q(n4846) );
  nnd2s1 U5159 ( .DIN1(n4847), .DIN2(n4848), .Q(N73) );
  nnd2s1 U5160 ( .DIN1(n4849), .DIN2(n1610), .Q(n4848) );
  xor2s1 U5161 ( .DIN1(n4850), .DIN2(n4851), .Q(n4849) );
  xnr2s1 U5162 ( .DIN1(n4852), .DIN2(n4761), .Q(n4851) );
  xor2s1 U5163 ( .DIN1(n4853), .DIN2(n4854), .Q(n4850) );
  xor2s1 U5164 ( .DIN1(n1415), .DIN2(n4772), .Q(n4854) );
  nnd2s1 U5165 ( .DIN1(n4855), .DIN2(n1606), .Q(n4847) );
  xor2s1 U5166 ( .DIN1(w3[23]), .DIN2(text_in_r[23]), .Q(n4855) );
  nnd3s1 U5167 ( .DIN1(n4856), .DIN2(n4857), .DIN3(n4858), .Q(N72) );
  nnd2s1 U5168 ( .DIN1(n1597), .DIN2(n4859), .Q(n4858) );
  xor2s1 U5169 ( .DIN1(w3[22]), .DIN2(text_in_r[22]), .Q(n4859) );
  nnd2s1 U5170 ( .DIN1(n4860), .DIN2(n4861), .Q(n4857) );
  nnd2s1 U5171 ( .DIN1(n4862), .DIN2(n4863), .Q(n4860) );
  nnd2s1 U5172 ( .DIN1(n4864), .DIN2(n4865), .Q(n4863) );
  nnd2s1 U5173 ( .DIN1(n4866), .DIN2(n4867), .Q(n4862) );
  nnd2s1 U5174 ( .DIN1(n4770), .DIN2(n4868), .Q(n4856) );
  nnd2s1 U5175 ( .DIN1(n4869), .DIN2(n4870), .Q(n4868) );
  nnd2s1 U5176 ( .DIN1(n4866), .DIN2(n4865), .Q(n4870) );
  nnd2s1 U5177 ( .DIN1(n4867), .DIN2(n4864), .Q(n4869) );
  hi1s1 U5178 ( .DIN(n4865), .Q(n4867) );
  xor2s1 U5179 ( .DIN1(n4871), .DIN2(n4872), .Q(n4865) );
  xor2s1 U5180 ( .DIN1(n1438), .DIN2(n4873), .Q(n4872) );
  nnd3s1 U5181 ( .DIN1(n4874), .DIN2(n4875), .DIN3(n4876), .Q(N71) );
  nnd2s1 U5182 ( .DIN1(n1597), .DIN2(n4877), .Q(n4876) );
  xor2s1 U5183 ( .DIN1(w3[21]), .DIN2(text_in_r[21]), .Q(n4877) );
  nnd2s1 U5184 ( .DIN1(n4878), .DIN2(n4879), .Q(n4875) );
  hi1s1 U5185 ( .DIN(n4779), .Q(n4879) );
  nnd2s1 U5186 ( .DIN1(n4880), .DIN2(n4881), .Q(n4878) );
  nnd2s1 U5187 ( .DIN1(n4882), .DIN2(n4883), .Q(n4881) );
  nnd2s1 U5188 ( .DIN1(n4884), .DIN2(n4885), .Q(n4880) );
  nnd2s1 U5189 ( .DIN1(n4779), .DIN2(n4886), .Q(n4874) );
  nnd2s1 U5190 ( .DIN1(n4887), .DIN2(n4888), .Q(n4886) );
  nnd2s1 U5191 ( .DIN1(n4884), .DIN2(n4883), .Q(n4888) );
  nnd2s1 U5192 ( .DIN1(n4885), .DIN2(n4882), .Q(n4887) );
  hi1s1 U5193 ( .DIN(n4883), .Q(n4885) );
  xor2s1 U5194 ( .DIN1(n4889), .DIN2(n4890), .Q(n4883) );
  xor2s1 U5195 ( .DIN1(n1373), .DIN2(n4891), .Q(n4890) );
  nnd2s1 U5196 ( .DIN1(n4892), .DIN2(n4893), .Q(N70) );
  nnd2s1 U5197 ( .DIN1(n4894), .DIN2(n1610), .Q(n4893) );
  xor2s1 U5198 ( .DIN1(n4895), .DIN2(n4896), .Q(n4894) );
  xor2s1 U5199 ( .DIN1(n4897), .DIN2(n4898), .Q(n4896) );
  xnr2s1 U5200 ( .DIN1(n4899), .DIN2(n4800), .Q(n4898) );
  xor2s1 U5201 ( .DIN1(n4819), .DIN2(n4900), .Q(n4895) );
  xor2s1 U5202 ( .DIN1(n1376), .DIN2(n4901), .Q(n4900) );
  nnd2s1 U5203 ( .DIN1(n4902), .DIN2(n1606), .Q(n4892) );
  xor2s1 U5204 ( .DIN1(w3[20]), .DIN2(text_in_r[20]), .Q(n4902) );
  nnd2s1 U5205 ( .DIN1(n4903), .DIN2(n4904), .Q(N69) );
  nnd2s1 U5206 ( .DIN1(n4905), .DIN2(n1611), .Q(n4904) );
  xor2s1 U5207 ( .DIN1(n4906), .DIN2(n4907), .Q(n4905) );
  xor2s1 U5208 ( .DIN1(n4908), .DIN2(n4909), .Q(n4907) );
  xor2s1 U5209 ( .DIN1(n4910), .DIN2(n4814), .Q(n4909) );
  hi1s1 U5210 ( .DIN(n4807), .Q(n4814) );
  xor2s1 U5211 ( .DIN1(n4827), .DIN2(n4911), .Q(n4906) );
  xor2s1 U5212 ( .DIN1(n1439), .DIN2(n4912), .Q(n4911) );
  nnd2s1 U5213 ( .DIN1(n4913), .DIN2(n1606), .Q(n4903) );
  xor2s1 U5214 ( .DIN1(w3[19]), .DIN2(text_in_r[19]), .Q(n4913) );
  nnd2s1 U5215 ( .DIN1(n4914), .DIN2(n4915), .Q(N68) );
  nnd2s1 U5216 ( .DIN1(n4916), .DIN2(n1611), .Q(n4915) );
  xor2s1 U5217 ( .DIN1(n4917), .DIN2(n4918), .Q(n4916) );
  xor2s1 U5218 ( .DIN1(n4919), .DIN2(n4920), .Q(n4918) );
  xor2s1 U5219 ( .DIN1(n4921), .DIN2(n4922), .Q(n4917) );
  xor2s1 U5220 ( .DIN1(n1368), .DIN2(n4923), .Q(n4922) );
  nnd2s1 U5221 ( .DIN1(n4924), .DIN2(n1606), .Q(n4914) );
  xor2s1 U5222 ( .DIN1(w3[18]), .DIN2(text_in_r[18]), .Q(n4924) );
  nnd2s1 U5223 ( .DIN1(n4925), .DIN2(n4926), .Q(N67) );
  nnd2s1 U5224 ( .DIN1(n4927), .DIN2(n1611), .Q(n4926) );
  xor2s1 U5225 ( .DIN1(n4928), .DIN2(n4929), .Q(n4927) );
  xor2s1 U5226 ( .DIN1(n4908), .DIN2(n4930), .Q(n4929) );
  xnr2s1 U5227 ( .DIN1(n4931), .DIN2(n4835), .Q(n4930) );
  xnr2s1 U5228 ( .DIN1(n4845), .DIN2(n1551), .Q(n4928) );
  nnd2s1 U5229 ( .DIN1(n4934), .DIN2(n1606), .Q(n4925) );
  xor2s1 U5230 ( .DIN1(w3[17]), .DIN2(text_in_r[17]), .Q(n4934) );
  nnd2s1 U5231 ( .DIN1(n4935), .DIN2(n4936), .Q(N66) );
  nnd2s1 U5232 ( .DIN1(n4937), .DIN2(n1612), .Q(n4936) );
  xor2s1 U5233 ( .DIN1(n4938), .DIN2(n4939), .Q(n4937) );
  xor2s1 U5234 ( .DIN1(n4844), .DIN2(n4897), .Q(n4939) );
  hi1s1 U5235 ( .DIN(n4908), .Q(n4897) );
  xnr2s1 U5236 ( .DIN1(n4940), .DIN2(n4763), .Q(n4908) );
  xor2s1 U5237 ( .DIN1(n1558), .DIN2(n4941), .Q(n4938) );
  nnd2s1 U5238 ( .DIN1(n4942), .DIN2(n1606), .Q(n4935) );
  xor2s1 U5239 ( .DIN1(n1559), .DIN2(text_in_r[16]), .Q(n4942) );
  nnd2s1 U5240 ( .DIN1(n4943), .DIN2(n4944), .Q(N57) );
  nnd2s1 U5241 ( .DIN1(n4945), .DIN2(n1612), .Q(n4944) );
  xor2s1 U5242 ( .DIN1(n4946), .DIN2(n4947), .Q(n4945) );
  xor2s1 U5243 ( .DIN1(n4770), .DIN2(n4795), .Q(n4947) );
  hi1s1 U5244 ( .DIN(n4861), .Q(n4770) );
  xnr2s1 U5245 ( .DIN1(n4948), .DIN2(n4853), .Q(n4861) );
  xor2s1 U5246 ( .DIN1(n1414), .DIN2(n4949), .Q(n4946) );
  nnd2s1 U5247 ( .DIN1(n4950), .DIN2(n1606), .Q(n4943) );
  xor2s1 U5248 ( .DIN1(w3[15]), .DIN2(text_in_r[15]), .Q(n4950) );
  nnd2s1 U5249 ( .DIN1(n4951), .DIN2(n4952), .Q(N56) );
  nnd2s1 U5250 ( .DIN1(n4953), .DIN2(n1612), .Q(n4952) );
  xor2s1 U5251 ( .DIN1(n4954), .DIN2(n4955), .Q(n4953) );
  xor2s1 U5252 ( .DIN1(n4956), .DIN2(n4779), .Q(n4955) );
  xor2s1 U5253 ( .DIN1(n4957), .DIN2(n4958), .Q(n4779) );
  xor2s1 U5254 ( .DIN1(n4948), .DIN2(w3[14]), .Q(n4954) );
  nnd2s1 U5255 ( .DIN1(n4959), .DIN2(n1606), .Q(n4951) );
  xor2s1 U5256 ( .DIN1(w3[14]), .DIN2(text_in_r[14]), .Q(n4959) );
  nnd2s1 U5257 ( .DIN1(n4960), .DIN2(n4961), .Q(N55) );
  nnd2s1 U5258 ( .DIN1(n4962), .DIN2(n1613), .Q(n4961) );
  xor2s1 U5259 ( .DIN1(n4963), .DIN2(n4964), .Q(n4962) );
  xor2s1 U5260 ( .DIN1(n4771), .DIN2(n4800), .Q(n4964) );
  xor2s1 U5261 ( .DIN1(n4889), .DIN2(n4965), .Q(n4800) );
  xor2s1 U5262 ( .DIN1(n1372), .DIN2(n4957), .Q(n4963) );
  nnd2s1 U5263 ( .DIN1(n4966), .DIN2(n1606), .Q(n4960) );
  xor2s1 U5264 ( .DIN1(w3[13]), .DIN2(text_in_r[13]), .Q(n4966) );
  nnd2s1 U5265 ( .DIN1(n4967), .DIN2(n4968), .Q(N54) );
  nnd2s1 U5266 ( .DIN1(n4969), .DIN2(n1613), .Q(n4968) );
  xor2s1 U5267 ( .DIN1(n4970), .DIN2(n4971), .Q(n4969) );
  xnr2s1 U5268 ( .DIN1(n4761), .DIN2(n4972), .Q(n4971) );
  xor2s1 U5269 ( .DIN1(n1393), .DIN2(n4965), .Q(n4972) );
  xor2s1 U5270 ( .DIN1(n4780), .DIN2(n4807), .Q(n4970) );
  xnr2s1 U5271 ( .DIN1(n4973), .DIN2(n4899), .Q(n4807) );
  nnd2s1 U5272 ( .DIN1(n4974), .DIN2(n1605), .Q(n4967) );
  xor2s1 U5273 ( .DIN1(w3[12]), .DIN2(text_in_r[12]), .Q(n4974) );
  nnd3s1 U5274 ( .DIN1(n4975), .DIN2(n4976), .DIN3(n4977), .Q(N53) );
  nnd2s1 U5275 ( .DIN1(n1597), .DIN2(n4978), .Q(n4977) );
  xor2s1 U5276 ( .DIN1(w3[11]), .DIN2(text_in_r[11]), .Q(n4978) );
  nnd2s1 U5277 ( .DIN1(n4979), .DIN2(n4980), .Q(n4976) );
  nnd2s1 U5278 ( .DIN1(n4981), .DIN2(n4982), .Q(n4979) );
  nnd2s1 U5279 ( .DIN1(n4791), .DIN2(n4920), .Q(n4982) );
  nnd2s1 U5280 ( .DIN1(n4825), .DIN2(n4793), .Q(n4981) );
  nnd2s1 U5281 ( .DIN1(n4983), .DIN2(n4984), .Q(n4975) );
  nnd2s1 U5282 ( .DIN1(n4985), .DIN2(n4986), .Q(n4984) );
  nnd2s1 U5283 ( .DIN1(n4793), .DIN2(n4920), .Q(n4986) );
  nor2s1 U5284 ( .DIN1(n4987), .DIN2(n1594), .Q(n4793) );
  nnd2s1 U5285 ( .DIN1(n4825), .DIN2(n4791), .Q(n4985) );
  nor2s1 U5286 ( .DIN1(n4988), .DIN2(n1595), .Q(n4791) );
  hi1s1 U5287 ( .DIN(n4987), .Q(n4988) );
  hi1s1 U5288 ( .DIN(n4920), .Q(n4825) );
  xnr2s1 U5289 ( .DIN1(n4989), .DIN2(n4910), .Q(n4920) );
  hi1s1 U5290 ( .DIN(n4980), .Q(n4983) );
  xnr2s1 U5291 ( .DIN1(n4761), .DIN2(n4990), .Q(n4980) );
  xor2s1 U5292 ( .DIN1(n4973), .DIN2(w3[11]), .Q(n4990) );
  nnd2s1 U5293 ( .DIN1(n4991), .DIN2(n4992), .Q(N52) );
  nnd2s1 U5294 ( .DIN1(n4993), .DIN2(n1613), .Q(n4992) );
  xor2s1 U5295 ( .DIN1(n4994), .DIN2(n4995), .Q(n4993) );
  xor2s1 U5296 ( .DIN1(n4996), .DIN2(n4835), .Q(n4995) );
  xor2s1 U5297 ( .DIN1(n4919), .DIN2(n4997), .Q(n4835) );
  xor2s1 U5298 ( .DIN1(n4989), .DIN2(w3[10]), .Q(n4994) );
  nnd2s1 U5299 ( .DIN1(n4998), .DIN2(n1605), .Q(n4991) );
  xor2s1 U5300 ( .DIN1(w3[10]), .DIN2(text_in_r[10]), .Q(n4998) );
  nnd2s1 U5301 ( .DIN1(n4999), .DIN2(n5000), .Q(N51) );
  nnd2s1 U5302 ( .DIN1(n5001), .DIN2(n1614), .Q(n5000) );
  xor2s1 U5303 ( .DIN1(n5002), .DIN2(n5003), .Q(n5001) );
  xnr2s1 U5304 ( .DIN1(n4761), .DIN2(n5004), .Q(n5003) );
  xor2s1 U5305 ( .DIN1(n1547), .DIN2(n4997), .Q(n5004) );
  xnr2s1 U5306 ( .DIN1(n4844), .DIN2(n1552), .Q(n5002) );
  xor2s1 U5307 ( .DIN1(n4931), .DIN2(n5005), .Q(n4844) );
  nnd2s1 U5308 ( .DIN1(n5006), .DIN2(n1605), .Q(n4999) );
  xor2s1 U5309 ( .DIN1(w3[9]), .DIN2(text_in_r[9]), .Q(n5006) );
  xor2s1 U5310 ( .DIN1(n1556), .DIN2(n5005), .Q(N505) );
  hi1s1 U5311 ( .DIN(n4997), .Q(n5007) );
  xor2s1 U5312 ( .DIN1(n4989), .DIN2(w3[2]), .Q(N503) );
  xor2s1 U5313 ( .DIN1(n4973), .DIN2(w3[3]), .Q(N502) );
  xor2s1 U5314 ( .DIN1(w3[4]), .DIN2(n4965), .Q(N501) );
  xor2s1 U5315 ( .DIN1(n1375), .DIN2(n4957), .Q(N500) );
  nnd2s1 U5316 ( .DIN1(n5008), .DIN2(n5009), .Q(N50) );
  nnd2s1 U5317 ( .DIN1(n5010), .DIN2(n1614), .Q(n5009) );
  xor2s1 U5318 ( .DIN1(n5011), .DIN2(n5012), .Q(n5010) );
  xnr2s1 U5319 ( .DIN1(n4761), .DIN2(n1546), .Q(n5012) );
  xnr2s1 U5320 ( .DIN1(n4940), .DIN2(n4949), .Q(n4761) );
  xor2s1 U5321 ( .DIN1(n1361), .DIN2(n5005), .Q(n5011) );
  hi1s1 U5322 ( .DIN(n5013), .Q(n5005) );
  nnd2s1 U5323 ( .DIN1(n5014), .DIN2(n1605), .Q(n5008) );
  xor2s1 U5324 ( .DIN1(w3[8]), .DIN2(text_in_r[8]), .Q(n5014) );
  xor2s1 U5325 ( .DIN1(n4948), .DIN2(w3[6]), .Q(N499) );
  xor2s1 U5326 ( .DIN1(n1442), .DIN2(n4949), .Q(N498) );
  xor2s1 U5327 ( .DIN1(n1450), .DIN2(n4745), .Q(N497) );
  xor2s1 U5328 ( .DIN1(n5015), .DIN2(w2[1]), .Q(N496) );
  xor2s1 U5329 ( .DIN1(w2[2]), .DIN2(n5016), .Q(N495) );
  xor2s1 U5330 ( .DIN1(n5017), .DIN2(w2[3]), .Q(N494) );
  xor2s1 U5331 ( .DIN1(w2[4]), .DIN2(n5018), .Q(N493) );
  xor2s1 U5332 ( .DIN1(n1462), .DIN2(n5019), .Q(N492) );
  xnr2s1 U5333 ( .DIN1(n5020), .DIN2(w2[6]), .Q(N491) );
  xnr2s1 U5334 ( .DIN1(w2[7]), .DIN2(n5021), .Q(N490) );
  xor2s1 U5335 ( .DIN1(n1497), .DIN2(n5022), .Q(N489) );
  xor2s1 U5336 ( .DIN1(w1[1]), .DIN2(n5023), .Q(N488) );
  xor2s1 U5337 ( .DIN1(w1[2]), .DIN2(n5024), .Q(N487) );
  xor2s1 U5338 ( .DIN1(n5025), .DIN2(w1[3]), .Q(N486) );
  xor2s1 U5339 ( .DIN1(n1496), .DIN2(n5026), .Q(N485) );
  xor2s1 U5340 ( .DIN1(n1495), .DIN2(n5027), .Q(N484) );
  xor2s1 U5341 ( .DIN1(n5028), .DIN2(w1[6]), .Q(N483) );
  xnr2s1 U5342 ( .DIN1(w1[7]), .DIN2(n5029), .Q(N482) );
  xor2s1 U5343 ( .DIN1(n1473), .DIN2(n5030), .Q(N481) );
  xor2s1 U5344 ( .DIN1(w0[1]), .DIN2(n5031), .Q(N480) );
  xor2s1 U5345 ( .DIN1(w0[2]), .DIN2(n5032), .Q(N479) );
  xor2s1 U5346 ( .DIN1(n5033), .DIN2(w0[3]), .Q(N478) );
  xor2s1 U5347 ( .DIN1(n1472), .DIN2(n5034), .Q(N477) );
  xor2s1 U5348 ( .DIN1(n1471), .DIN2(n5035), .Q(N476) );
  xor2s1 U5349 ( .DIN1(n5036), .DIN2(w0[6]), .Q(N475) );
  xnr2s1 U5350 ( .DIN1(w0[7]), .DIN2(n5037), .Q(N474) );
  xor2s1 U5351 ( .DIN1(w3[9]), .DIN2(n4919), .Q(N472) );
  xor2s1 U5352 ( .DIN1(n4910), .DIN2(w3[10]), .Q(N471) );
  xor2s1 U5353 ( .DIN1(n4899), .DIN2(w3[11]), .Q(N470) );
  xor2s1 U5354 ( .DIN1(w3[12]), .DIN2(n4889), .Q(N469) );
  xor2s1 U5355 ( .DIN1(n1372), .DIN2(n4958), .Q(N468) );
  hi1s1 U5356 ( .DIN(n4871), .Q(n4958) );
  xor2s1 U5357 ( .DIN1(n4853), .DIN2(w3[14]), .Q(N467) );
  xor2s1 U5358 ( .DIN1(n1414), .DIN2(n4940), .Q(N466) );
  xor2s1 U5359 ( .DIN1(n1461), .DIN2(n4754), .Q(N465) );
  xor2s1 U5360 ( .DIN1(w2[9]), .DIN2(n5038), .Q(N464) );
  xor2s1 U5361 ( .DIN1(w2[10]), .DIN2(n5039), .Q(N463) );
  xor2s1 U5362 ( .DIN1(n5040), .DIN2(w2[11]), .Q(N462) );
  xor2s1 U5363 ( .DIN1(n1460), .DIN2(n5041), .Q(N461) );
  xor2s1 U5364 ( .DIN1(n1459), .DIN2(n5042), .Q(N460) );
  xor2s1 U5365 ( .DIN1(n5043), .DIN2(w2[14]), .Q(N459) );
  xor2s1 U5366 ( .DIN1(n1458), .DIN2(n5044), .Q(N458) );
  xor2s1 U5367 ( .DIN1(n1494), .DIN2(n5045), .Q(N457) );
  xor2s1 U5368 ( .DIN1(n5046), .DIN2(w1[9]), .Q(N456) );
  xor2s1 U5369 ( .DIN1(w1[10]), .DIN2(n5047), .Q(N455) );
  xor2s1 U5370 ( .DIN1(n5048), .DIN2(w1[11]), .Q(N454) );
  xor2s1 U5371 ( .DIN1(n1493), .DIN2(n5049), .Q(N453) );
  xor2s1 U5372 ( .DIN1(n1492), .DIN2(n5050), .Q(N452) );
  xor2s1 U5373 ( .DIN1(n5051), .DIN2(w1[14]), .Q(N451) );
  xor2s1 U5374 ( .DIN1(n1491), .DIN2(n5052), .Q(N450) );
  xor2s1 U5375 ( .DIN1(n1470), .DIN2(n5053), .Q(N449) );
  xor2s1 U5376 ( .DIN1(n5054), .DIN2(w0[9]), .Q(N448) );
  xor2s1 U5377 ( .DIN1(w0[10]), .DIN2(n5055), .Q(N447) );
  xor2s1 U5378 ( .DIN1(n5056), .DIN2(w0[11]), .Q(N446) );
  xor2s1 U5379 ( .DIN1(n1469), .DIN2(n5057), .Q(N445) );
  xor2s1 U5380 ( .DIN1(n1468), .DIN2(n5058), .Q(N444) );
  xor2s1 U5381 ( .DIN1(n5059), .DIN2(w0[14]), .Q(N443) );
  xor2s1 U5382 ( .DIN1(n1467), .DIN2(n5060), .Q(N442) );
  xor2s1 U5383 ( .DIN1(n1558), .DIN2(n4845), .Q(N441) );
  xor2s1 U5384 ( .DIN1(n4827), .DIN2(w3[18]), .Q(N439) );
  xor2s1 U5385 ( .DIN1(n4819), .DIN2(w3[19]), .Q(N438) );
  xor2s1 U5386 ( .DIN1(n1376), .DIN2(n4801), .Q(N437) );
  hi1s1 U5387 ( .DIN(n4891), .Q(n4801) );
  xor2s1 U5388 ( .DIN1(n1373), .DIN2(n4781), .Q(N436) );
  xor2s1 U5389 ( .DIN1(n4772), .DIN2(w3[22]), .Q(N435) );
  xor2s1 U5390 ( .DIN1(n1415), .DIN2(n4763), .Q(N434) );
  xor2s1 U5391 ( .DIN1(n1457), .DIN2(n5061), .Q(N433) );
  xor2s1 U5392 ( .DIN1(n1456), .DIN2(n5062), .Q(N432) );
  xor2s1 U5393 ( .DIN1(w2[18]), .DIN2(n5063), .Q(N431) );
  xor2s1 U5394 ( .DIN1(n5064), .DIN2(w2[19]), .Q(N430) );
  xor2s1 U5395 ( .DIN1(n1455), .DIN2(n5065), .Q(N429) );
  xnr2s1 U5396 ( .DIN1(w2[21]), .DIN2(n5066), .Q(N428) );
  xor2s1 U5397 ( .DIN1(n5067), .DIN2(w2[22]), .Q(N427) );
  xor2s1 U5398 ( .DIN1(w2[23]), .DIN2(n5068), .Q(N426) );
  xor2s1 U5399 ( .DIN1(n1490), .DIN2(n5069), .Q(N425) );
  xor2s1 U5400 ( .DIN1(n5070), .DIN2(w1[17]), .Q(N424) );
  xor2s1 U5401 ( .DIN1(n1489), .DIN2(n5071), .Q(N423) );
  xor2s1 U5402 ( .DIN1(n5072), .DIN2(w1[19]), .Q(N422) );
  xor2s1 U5403 ( .DIN1(n1488), .DIN2(n5073), .Q(N421) );
  xnr2s1 U5404 ( .DIN1(w1[21]), .DIN2(n5074), .Q(N420) );
  xor2s1 U5405 ( .DIN1(n5075), .DIN2(w1[22]), .Q(N419) );
  xor2s1 U5406 ( .DIN1(n1487), .DIN2(n5076), .Q(N418) );
  xor2s1 U5407 ( .DIN1(n1466), .DIN2(n5077), .Q(N417) );
  xor2s1 U5408 ( .DIN1(n5078), .DIN2(w0[17]), .Q(N416) );
  xor2s1 U5409 ( .DIN1(n1465), .DIN2(n5079), .Q(N415) );
  xor2s1 U5410 ( .DIN1(n5080), .DIN2(w0[19]), .Q(N414) );
  xor2s1 U5411 ( .DIN1(n1464), .DIN2(n5081), .Q(N413) );
  xnr2s1 U5412 ( .DIN1(w0[21]), .DIN2(n5082), .Q(N412) );
  xor2s1 U5413 ( .DIN1(n5083), .DIN2(w0[22]), .Q(N411) );
  xor2s1 U5414 ( .DIN1(n1463), .DIN2(n5084), .Q(N410) );
  nnd3s1 U5415 ( .DIN1(n5085), .DIN2(n5086), .DIN3(n5087), .Q(N41) );
  nnd2s1 U5416 ( .DIN1(n1597), .DIN2(n5088), .Q(n5087) );
  xor2s1 U5417 ( .DIN1(w3[7]), .DIN2(text_in_r[7]), .Q(n5088) );
  nnd2s1 U5418 ( .DIN1(n5089), .DIN2(n5090), .Q(n5086) );
  nnd2s1 U5419 ( .DIN1(n5091), .DIN2(n5092), .Q(n5089) );
  nnd2s1 U5420 ( .DIN1(n4864), .DIN2(n4788), .Q(n5092) );
  nnd2s1 U5421 ( .DIN1(n4866), .DIN2(n4795), .Q(n5091) );
  nnd2s1 U5422 ( .DIN1(n5093), .DIN2(n5094), .Q(n5085) );
  nnd2s1 U5423 ( .DIN1(n5095), .DIN2(n5096), .Q(n5094) );
  nnd2s1 U5424 ( .DIN1(n4866), .DIN2(n4788), .Q(n5096) );
  nor2s1 U5425 ( .DIN1(n5097), .DIN2(n1594), .Q(n4866) );
  nnd2s1 U5426 ( .DIN1(n4864), .DIN2(n4795), .Q(n5095) );
  hi1s1 U5427 ( .DIN(n4788), .Q(n4795) );
  xnr2s1 U5428 ( .DIN1(n4852), .DIN2(n4763), .Q(n4788) );
  nor4s1 U5429 ( .DIN1(n5098), .DIN2(n5099), .DIN3(n5100), .DIN4(n5101), 
        .Q(n4763) );
  nnd4s1 U5430 ( .DIN1(n5102), .DIN2(n5103), .DIN3(n5104), .DIN4(n5105), 
        .Q(n5101) );
  nnd2s1 U5431 ( .DIN1(n5106), .DIN2(n5107), .Q(n5105) );
  nnd2s1 U5432 ( .DIN1(n5108), .DIN2(n5109), .Q(n5104) );
  nnd2s1 U5433 ( .DIN1(n5110), .DIN2(n5111), .Q(n5103) );
  nnd4s1 U5434 ( .DIN1(n5112), .DIN2(n5113), .DIN3(n5114), .DIN4(n5115), 
        .Q(n5100) );
  nnd2s1 U5435 ( .DIN1(n5116), .DIN2(n5117), .Q(n5115) );
  nnd2s1 U5436 ( .DIN1(n5118), .DIN2(n5119), .Q(n5117) );
  nnd2s1 U5437 ( .DIN1(n5120), .DIN2(n5121), .Q(n5114) );
  nnd2s1 U5438 ( .DIN1(n5122), .DIN2(n5123), .Q(n5121) );
  nnd2s1 U5439 ( .DIN1(n5124), .DIN2(n5125), .Q(n5113) );
  nnd2s1 U5440 ( .DIN1(n5126), .DIN2(n5127), .Q(n5125) );
  nnd2s1 U5441 ( .DIN1(n5128), .DIN2(n5129), .Q(n5112) );
  nnd3s1 U5442 ( .DIN1(n5130), .DIN2(n5131), .DIN3(n5132), .Q(n5099) );
  nnd4s1 U5443 ( .DIN1(n5133), .DIN2(n5134), .DIN3(n5135), .DIN4(n5136), 
        .Q(n5098) );
  nnd2s1 U5444 ( .DIN1(n5137), .DIN2(n5138), .Q(n5135) );
  nnd2s1 U5445 ( .DIN1(n5139), .DIN2(n5140), .Q(n5134) );
  nor2s1 U5446 ( .DIN1(n5141), .DIN2(n1595), .Q(n4864) );
  hi1s1 U5447 ( .DIN(n5097), .Q(n5141) );
  hi1s1 U5448 ( .DIN(n5090), .Q(n5093) );
  xor2s1 U5449 ( .DIN1(n4948), .DIN2(n5142), .Q(n5090) );
  xor2s1 U5450 ( .DIN1(w3[7]), .DIN2(n4940), .Q(n5142) );
  nor4s1 U5451 ( .DIN1(n5143), .DIN2(n5144), .DIN3(n5145), .DIN4(n5146), 
        .Q(n4940) );
  nnd4s1 U5452 ( .DIN1(n5147), .DIN2(n5148), .DIN3(n5149), .DIN4(n5150), 
        .Q(n5146) );
  nnd2s1 U5453 ( .DIN1(n5151), .DIN2(n5152), .Q(n5150) );
  nnd2s1 U5454 ( .DIN1(n5153), .DIN2(n5154), .Q(n5149) );
  nnd2s1 U5455 ( .DIN1(n5155), .DIN2(n5156), .Q(n5148) );
  nnd4s1 U5456 ( .DIN1(n5157), .DIN2(n5158), .DIN3(n5159), .DIN4(n5160), 
        .Q(n5145) );
  nnd2s1 U5457 ( .DIN1(n5161), .DIN2(n5162), .Q(n5160) );
  nnd2s1 U5458 ( .DIN1(n5163), .DIN2(n5164), .Q(n5162) );
  nnd2s1 U5459 ( .DIN1(n5165), .DIN2(n5166), .Q(n5159) );
  nnd2s1 U5460 ( .DIN1(n5167), .DIN2(n5168), .Q(n5166) );
  nnd2s1 U5461 ( .DIN1(n5169), .DIN2(n5170), .Q(n5158) );
  nnd2s1 U5462 ( .DIN1(n5171), .DIN2(n5172), .Q(n5170) );
  nnd2s1 U5463 ( .DIN1(n5173), .DIN2(n5174), .Q(n5157) );
  nnd3s1 U5464 ( .DIN1(n5175), .DIN2(n5176), .DIN3(n5177), .Q(n5144) );
  nnd4s1 U5465 ( .DIN1(n5178), .DIN2(n5179), .DIN3(n5180), .DIN4(n5181), 
        .Q(n5143) );
  nnd2s1 U5466 ( .DIN1(n5182), .DIN2(n5183), .Q(n5180) );
  nnd2s1 U5467 ( .DIN1(n5184), .DIN2(n5185), .Q(n5179) );
  or3s1 U5468 ( .DIN1(n5186), .DIN2(n5187), .DIN3(n5188), .Q(n4948) );
  nnd4s1 U5469 ( .DIN1(n5189), .DIN2(n5190), .DIN3(n5191), .DIN4(n5192), 
        .Q(n5188) );
  and3s1 U5470 ( .DIN1(n5193), .DIN2(n5194), .DIN3(n5195), .Q(n5192) );
  nnd2s1 U5471 ( .DIN1(n5196), .DIN2(n5197), .Q(n5189) );
  nnd3s1 U5472 ( .DIN1(n5198), .DIN2(n5199), .DIN3(n5200), .Q(n5187) );
  or2s1 U5473 ( .DIN1(n5201), .DIN2(n5202), .Q(n5200) );
  or2s1 U5474 ( .DIN1(n5203), .DIN2(n5204), .Q(n5199) );
  nnd2s1 U5475 ( .DIN1(n5205), .DIN2(n5206), .Q(n5198) );
  nnd3s1 U5476 ( .DIN1(n5207), .DIN2(n5208), .DIN3(n5209), .Q(n5186) );
  nnd2s1 U5477 ( .DIN1(n5210), .DIN2(n5211), .Q(n5209) );
  nnd2s1 U5478 ( .DIN1(n5212), .DIN2(n5213), .Q(n5211) );
  nnd2s1 U5479 ( .DIN1(n5214), .DIN2(n5215), .Q(n5208) );
  nnd2s1 U5480 ( .DIN1(n5216), .DIN2(n5217), .Q(n5215) );
  hi1s1 U5481 ( .DIN(n5218), .Q(n5217) );
  nnd2s1 U5482 ( .DIN1(n5219), .DIN2(n5220), .Q(n5207) );
  nnd2s1 U5483 ( .DIN1(n5221), .DIN2(n5222), .Q(n5220) );
  xor2s1 U5484 ( .DIN1(n1554), .DIN2(n4941), .Q(N409) );
  xor2s1 U5485 ( .DIN1(n4923), .DIN2(w3[26]), .Q(N407) );
  xor2s1 U5486 ( .DIN1(n4912), .DIN2(w3[27]), .Q(N406) );
  xor2s1 U5487 ( .DIN1(w3[28]), .DIN2(n4901), .Q(N405) );
  xor2s1 U5488 ( .DIN1(n1374), .DIN2(n5224), .Q(N404) );
  xor2s1 U5489 ( .DIN1(n5097), .DIN2(w3[30]), .Q(N403) );
  xor2s1 U5490 ( .DIN1(n1416), .DIN2(n4852), .Q(N402) );
  xor2s1 U5491 ( .DIN1(n1454), .DIN2(n4741), .Q(N401) );
  xor2s1 U5492 ( .DIN1(w2[25]), .DIN2(n5225), .Q(N400) );
  nnd3s1 U5493 ( .DIN1(n5226), .DIN2(n5227), .DIN3(n5228), .Q(N40) );
  nnd2s1 U5494 ( .DIN1(n1597), .DIN2(n5229), .Q(n5228) );
  xor2s1 U5495 ( .DIN1(w3[6]), .DIN2(text_in_r[6]), .Q(n5229) );
  nnd2s1 U5496 ( .DIN1(n5230), .DIN2(n5231), .Q(n5227) );
  nnd2s1 U5497 ( .DIN1(n5232), .DIN2(n5233), .Q(n5230) );
  nnd2s1 U5498 ( .DIN1(n4882), .DIN2(n4762), .Q(n5233) );
  nnd2s1 U5499 ( .DIN1(n4956), .DIN2(n4884), .Q(n5232) );
  nnd2s1 U5500 ( .DIN1(n5234), .DIN2(n5235), .Q(n5226) );
  nnd2s1 U5501 ( .DIN1(n5236), .DIN2(n5237), .Q(n5235) );
  nnd2s1 U5502 ( .DIN1(n4884), .DIN2(n4762), .Q(n5237) );
  hi1s1 U5503 ( .DIN(n4956), .Q(n4762) );
  nor2s1 U5504 ( .DIN1(n5238), .DIN2(n1594), .Q(n4884) );
  nnd2s1 U5505 ( .DIN1(n4956), .DIN2(n4882), .Q(n5236) );
  nor2s1 U5506 ( .DIN1(n5224), .DIN2(n1595), .Q(n4882) );
  hi1s1 U5507 ( .DIN(n5238), .Q(n5224) );
  xor2s1 U5508 ( .DIN1(n5097), .DIN2(n4772), .Q(n4956) );
  or3s1 U5509 ( .DIN1(n5239), .DIN2(n5240), .DIN3(n5241), .Q(n4772) );
  nnd4s1 U5510 ( .DIN1(n5242), .DIN2(n5243), .DIN3(n5244), .DIN4(n5245), 
        .Q(n5241) );
  and3s1 U5511 ( .DIN1(n5246), .DIN2(n5247), .DIN3(n5248), .Q(n5245) );
  nnd2s1 U5512 ( .DIN1(n5249), .DIN2(n5108), .Q(n5243) );
  nnd2s1 U5513 ( .DIN1(n5138), .DIN2(n5250), .Q(n5242) );
  nnd3s1 U5514 ( .DIN1(n5251), .DIN2(n5252), .DIN3(n5253), .Q(n5240) );
  or2s1 U5515 ( .DIN1(n5254), .DIN2(n5255), .Q(n5253) );
  or2s1 U5516 ( .DIN1(n5123), .DIN2(n5256), .Q(n5252) );
  nnd2s1 U5517 ( .DIN1(n5124), .DIN2(n5257), .Q(n5251) );
  nnd3s1 U5518 ( .DIN1(n5258), .DIN2(n5259), .DIN3(n5260), .Q(n5239) );
  nnd2s1 U5519 ( .DIN1(n5261), .DIN2(n5262), .Q(n5260) );
  nnd2s1 U5520 ( .DIN1(n5263), .DIN2(n5264), .Q(n5262) );
  nnd2s1 U5521 ( .DIN1(n5265), .DIN2(n5266), .Q(n5259) );
  nnd2s1 U5522 ( .DIN1(n5267), .DIN2(n5268), .Q(n5266) );
  nnd2s1 U5523 ( .DIN1(n5139), .DIN2(n5269), .Q(n5258) );
  nnd2s1 U5524 ( .DIN1(n5270), .DIN2(n5271), .Q(n5269) );
  hi1s1 U5525 ( .DIN(n5272), .Q(n5271) );
  or3s1 U5526 ( .DIN1(n5273), .DIN2(n5274), .DIN3(n5275), .Q(n5097) );
  nnd4s1 U5527 ( .DIN1(n5276), .DIN2(n5277), .DIN3(n5278), .DIN4(n5279), 
        .Q(n5275) );
  and3s1 U5528 ( .DIN1(n5280), .DIN2(n5281), .DIN3(n5282), .Q(n5279) );
  nnd2s1 U5529 ( .DIN1(n5283), .DIN2(n5284), .Q(n5277) );
  nnd2s1 U5530 ( .DIN1(n5285), .DIN2(n5286), .Q(n5276) );
  nnd3s1 U5531 ( .DIN1(n5287), .DIN2(n5288), .DIN3(n5289), .Q(n5274) );
  or2s1 U5532 ( .DIN1(n5290), .DIN2(n5291), .Q(n5289) );
  or2s1 U5533 ( .DIN1(n5292), .DIN2(n5293), .Q(n5288) );
  nnd2s1 U5534 ( .DIN1(n5294), .DIN2(n5295), .Q(n5287) );
  nnd3s1 U5535 ( .DIN1(n5296), .DIN2(n5297), .DIN3(n5298), .Q(n5273) );
  nnd2s1 U5536 ( .DIN1(n5299), .DIN2(n5300), .Q(n5298) );
  nnd2s1 U5537 ( .DIN1(n5301), .DIN2(n5302), .Q(n5300) );
  nnd2s1 U5538 ( .DIN1(n5303), .DIN2(n5304), .Q(n5297) );
  nnd2s1 U5539 ( .DIN1(n5305), .DIN2(n5306), .Q(n5304) );
  nnd2s1 U5540 ( .DIN1(n5307), .DIN2(n5308), .Q(n5296) );
  nnd2s1 U5541 ( .DIN1(n5309), .DIN2(n5310), .Q(n5308) );
  hi1s1 U5542 ( .DIN(n5311), .Q(n5310) );
  hi1s1 U5543 ( .DIN(n5231), .Q(n5234) );
  xnr2s1 U5544 ( .DIN1(n4957), .DIN2(n5312), .Q(n5231) );
  xor2s1 U5545 ( .DIN1(n1391), .DIN2(n4853), .Q(n5312) );
  or3s1 U5546 ( .DIN1(n5313), .DIN2(n5314), .DIN3(n5315), .Q(n4853) );
  nnd4s1 U5547 ( .DIN1(n5316), .DIN2(n5317), .DIN3(n5318), .DIN4(n5319), 
        .Q(n5315) );
  and3s1 U5548 ( .DIN1(n5320), .DIN2(n5321), .DIN3(n5322), .Q(n5319) );
  nnd2s1 U5549 ( .DIN1(n5323), .DIN2(n5153), .Q(n5317) );
  nnd2s1 U5550 ( .DIN1(n5183), .DIN2(n5324), .Q(n5316) );
  nnd3s1 U5551 ( .DIN1(n5325), .DIN2(n5326), .DIN3(n5327), .Q(n5314) );
  or2s1 U5552 ( .DIN1(n5328), .DIN2(n5329), .Q(n5327) );
  or2s1 U5553 ( .DIN1(n5168), .DIN2(n5330), .Q(n5326) );
  nnd2s1 U5554 ( .DIN1(n5169), .DIN2(n5331), .Q(n5325) );
  nnd3s1 U5555 ( .DIN1(n5332), .DIN2(n5333), .DIN3(n5334), .Q(n5313) );
  nnd2s1 U5556 ( .DIN1(n5335), .DIN2(n5336), .Q(n5334) );
  nnd2s1 U5557 ( .DIN1(n5337), .DIN2(n5338), .Q(n5336) );
  nnd2s1 U5558 ( .DIN1(n5339), .DIN2(n5340), .Q(n5333) );
  nnd2s1 U5559 ( .DIN1(n5341), .DIN2(n5342), .Q(n5340) );
  nnd2s1 U5560 ( .DIN1(n5184), .DIN2(n5343), .Q(n5332) );
  nnd2s1 U5561 ( .DIN1(n5344), .DIN2(n5345), .Q(n5343) );
  hi1s1 U5562 ( .DIN(n5346), .Q(n5345) );
  nor3s1 U5563 ( .DIN1(n5347), .DIN2(n5348), .DIN3(n5349), .Q(n4957) );
  nnd4s1 U5564 ( .DIN1(n5350), .DIN2(n5194), .DIN3(n5351), .DIN4(n5352), 
        .Q(n5349) );
  and4s1 U5565 ( .DIN1(n5353), .DIN2(n5354), .DIN3(n5355), .DIN4(n5356), 
        .Q(n5352) );
  nnd2s1 U5566 ( .DIN1(n5196), .DIN2(n5357), .Q(n5356) );
  nnd2s1 U5567 ( .DIN1(n5210), .DIN2(n5358), .Q(n5355) );
  nnd2s1 U5568 ( .DIN1(n5359), .DIN2(n5219), .Q(n5354) );
  nor2s1 U5569 ( .DIN1(n5360), .DIN2(n5361), .Q(n5194) );
  nnd4s1 U5570 ( .DIN1(n5362), .DIN2(n5363), .DIN3(n5364), .DIN4(n5365), 
        .Q(n5361) );
  nnd2s1 U5571 ( .DIN1(n5366), .DIN2(n5367), .Q(n5365) );
  nnd3s1 U5572 ( .DIN1(n5222), .DIN2(n5368), .DIN3(n5369), .Q(n5367) );
  nnd2s1 U5573 ( .DIN1(n5370), .DIN2(n5371), .Q(n5364) );
  nnd2s1 U5574 ( .DIN1(n5359), .DIN2(n5372), .Q(n5363) );
  nnd2s1 U5575 ( .DIN1(n5373), .DIN2(n5357), .Q(n5362) );
  nnd4s1 U5576 ( .DIN1(n5374), .DIN2(n5375), .DIN3(n5376), .DIN4(n5377), 
        .Q(n5360) );
  nnd2s1 U5577 ( .DIN1(n5378), .DIN2(n5379), .Q(n5377) );
  nnd2s1 U5578 ( .DIN1(n5380), .DIN2(n5381), .Q(n5379) );
  nnd2s1 U5579 ( .DIN1(n5358), .DIN2(n5382), .Q(n5376) );
  nnd2s1 U5580 ( .DIN1(n5383), .DIN2(n5384), .Q(n5382) );
  nnd2s1 U5581 ( .DIN1(n5385), .DIN2(n5386), .Q(n5375) );
  nnd2s1 U5582 ( .DIN1(n5387), .DIN2(n5213), .Q(n5386) );
  nnd2s1 U5583 ( .DIN1(n5388), .DIN2(n5389), .Q(n5374) );
  nnd2s1 U5584 ( .DIN1(n5222), .DIN2(n5390), .Q(n5389) );
  nnd4s1 U5585 ( .DIN1(n5391), .DIN2(n5392), .DIN3(n5393), .DIN4(n5394), 
        .Q(n5348) );
  or2s1 U5586 ( .DIN1(n5395), .DIN2(n5396), .Q(n5394) );
  nnd2s1 U5587 ( .DIN1(n5373), .DIN2(n5397), .Q(n5393) );
  nnd2s1 U5588 ( .DIN1(n5398), .DIN2(n5399), .Q(n5392) );
  nnd2s1 U5589 ( .DIN1(n5370), .DIN2(n5400), .Q(n5391) );
  nnd4s1 U5590 ( .DIN1(n5401), .DIN2(n5402), .DIN3(n5403), .DIN4(n5404), 
        .Q(n5347) );
  nnd2s1 U5591 ( .DIN1(n5405), .DIN2(n5406), .Q(n5404) );
  nnd2s1 U5592 ( .DIN1(n5368), .DIN2(n5407), .Q(n5406) );
  nnd2s1 U5593 ( .DIN1(n5408), .DIN2(n5409), .Q(n5403) );
  nnd2s1 U5594 ( .DIN1(n5212), .DIN2(n5410), .Q(n5409) );
  nnd2s1 U5595 ( .DIN1(n5205), .DIN2(n5411), .Q(n5402) );
  nnd2s1 U5596 ( .DIN1(n5412), .DIN2(n5413), .Q(n5411) );
  nnd2s1 U5597 ( .DIN1(n5414), .DIN2(n5415), .Q(n5401) );
  xor2s1 U5598 ( .DIN1(n1453), .DIN2(n5416), .Q(N399) );
  xor2s1 U5599 ( .DIN1(w2[27]), .DIN2(n5417), .Q(N398) );
  xor2s1 U5600 ( .DIN1(w2[28]), .DIN2(n5418), .Q(N397) );
  xor2s1 U5601 ( .DIN1(n1452), .DIN2(n5419), .Q(N396) );
  xor2s1 U5602 ( .DIN1(n5420), .DIN2(w2[30]), .Q(N395) );
  xor2s1 U5603 ( .DIN1(n1451), .DIN2(n5421), .Q(N394) );
  xor2s1 U5604 ( .DIN1(n1486), .DIN2(n5422), .Q(N393) );
  xor2s1 U5605 ( .DIN1(n5423), .DIN2(w1[25]), .Q(N392) );
  xor2s1 U5606 ( .DIN1(w1[26]), .DIN2(n5424), .Q(N391) );
  xor2s1 U5607 ( .DIN1(n5425), .DIN2(w1[27]), .Q(N390) );
  nnd2s1 U5608 ( .DIN1(n5426), .DIN2(n5427), .Q(N39) );
  nnd2s1 U5609 ( .DIN1(n5428), .DIN2(n1614), .Q(n5427) );
  xor2s1 U5610 ( .DIN1(n5429), .DIN2(n5430), .Q(n5428) );
  xnr2s1 U5611 ( .DIN1(n4965), .DIN2(n4771), .Q(n5430) );
  xnr2s1 U5612 ( .DIN1(n5238), .DIN2(n4781), .Q(n4771) );
  hi1s1 U5613 ( .DIN(n4873), .Q(n4781) );
  or3s1 U5614 ( .DIN1(n5431), .DIN2(n5432), .DIN3(n5433), .Q(n4873) );
  nnd4s1 U5615 ( .DIN1(n5434), .DIN2(n5247), .DIN3(n5435), .DIN4(n5436), 
        .Q(n5433) );
  and4s1 U5616 ( .DIN1(n5437), .DIN2(n5438), .DIN3(n5439), .DIN4(n5136), 
        .Q(n5436) );
  nnd2s1 U5617 ( .DIN1(n5440), .DIN2(n5265), .Q(n5136) );
  nnd2s1 U5618 ( .DIN1(n5261), .DIN2(n5441), .Q(n5439) );
  nnd2s1 U5619 ( .DIN1(n5442), .DIN2(n5140), .Q(n5438) );
  nor2s1 U5620 ( .DIN1(n5443), .DIN2(n5444), .Q(n5247) );
  nnd4s1 U5621 ( .DIN1(n5445), .DIN2(n5446), .DIN3(n5447), .DIN4(n5448), 
        .Q(n5444) );
  or2s1 U5622 ( .DIN1(n5449), .DIN2(n5450), .Q(n5448) );
  nnd2s1 U5623 ( .DIN1(n5442), .DIN2(n5451), .Q(n5447) );
  nnd2s1 U5624 ( .DIN1(n5440), .DIN2(n5138), .Q(n5446) );
  nnd2s1 U5625 ( .DIN1(n5111), .DIN2(n5452), .Q(n5445) );
  nnd4s1 U5626 ( .DIN1(n5453), .DIN2(n5454), .DIN3(n5455), .DIN4(n5456), 
        .Q(n5443) );
  nnd2s1 U5627 ( .DIN1(n5110), .DIN2(n5457), .Q(n5456) );
  nnd2s1 U5628 ( .DIN1(n5267), .DIN2(n5458), .Q(n5457) );
  nnd2s1 U5629 ( .DIN1(n5459), .DIN2(n5460), .Q(n5455) );
  nnd2s1 U5630 ( .DIN1(n5263), .DIN2(n5461), .Q(n5460) );
  nnd2s1 U5631 ( .DIN1(n5441), .DIN2(n5462), .Q(n5454) );
  nnd2s1 U5632 ( .DIN1(n5463), .DIN2(n5464), .Q(n5462) );
  nnd2s1 U5633 ( .DIN1(n5120), .DIN2(n5465), .Q(n5453) );
  nnd3s1 U5634 ( .DIN1(n5267), .DIN2(n5466), .DIN3(n5467), .Q(n5465) );
  nnd4s1 U5635 ( .DIN1(n5468), .DIN2(n5469), .DIN3(n5470), .DIN4(n5471), 
        .Q(n5432) );
  nnd2s1 U5636 ( .DIN1(n5472), .DIN2(n5473), .Q(n5471) );
  nnd2s1 U5637 ( .DIN1(n5111), .DIN2(n5474), .Q(n5470) );
  nnd2s1 U5638 ( .DIN1(n5137), .DIN2(n5475), .Q(n5469) );
  nnd2s1 U5639 ( .DIN1(n5249), .DIN2(n5452), .Q(n5468) );
  nnd4s1 U5640 ( .DIN1(n5476), .DIN2(n5477), .DIN3(n5478), .DIN4(n5479), 
        .Q(n5431) );
  nnd2s1 U5641 ( .DIN1(n5128), .DIN2(n5480), .Q(n5479) );
  nnd2s1 U5642 ( .DIN1(n5264), .DIN2(n5481), .Q(n5480) );
  nnd2s1 U5643 ( .DIN1(n5482), .DIN2(n5483), .Q(n5478) );
  nnd2s1 U5644 ( .DIN1(n5124), .DIN2(n5484), .Q(n5477) );
  nnd2s1 U5645 ( .DIN1(n5485), .DIN2(n5119), .Q(n5484) );
  nnd2s1 U5646 ( .DIN1(n5108), .DIN2(n5486), .Q(n5476) );
  or3s1 U5647 ( .DIN1(n5487), .DIN2(n5488), .DIN3(n5489), .Q(n5238) );
  nnd4s1 U5648 ( .DIN1(n5490), .DIN2(n5281), .DIN3(n5491), .DIN4(n5492), 
        .Q(n5489) );
  and4s1 U5649 ( .DIN1(n5493), .DIN2(n5494), .DIN3(n5495), .DIN4(n5496), 
        .Q(n5492) );
  nnd2s1 U5650 ( .DIN1(n5497), .DIN2(n5299), .Q(n5495) );
  nnd2s1 U5651 ( .DIN1(n5498), .DIN2(n5499), .Q(n5494) );
  nor2s1 U5652 ( .DIN1(n5500), .DIN2(n5501), .Q(n5281) );
  nnd4s1 U5653 ( .DIN1(n5502), .DIN2(n5503), .DIN3(n5504), .DIN4(n5505), 
        .Q(n5501) );
  or2s1 U5654 ( .DIN1(n5506), .DIN2(n5507), .Q(n5505) );
  nnd2s1 U5655 ( .DIN1(n5508), .DIN2(n5499), .Q(n5504) );
  nnd2s1 U5656 ( .DIN1(n5286), .DIN2(n5509), .Q(n5503) );
  nnd2s1 U5657 ( .DIN1(n5510), .DIN2(n5511), .Q(n5502) );
  nnd4s1 U5658 ( .DIN1(n5512), .DIN2(n5513), .DIN3(n5514), .DIN4(n5515), 
        .Q(n5500) );
  nnd2s1 U5659 ( .DIN1(n5516), .DIN2(n5517), .Q(n5515) );
  nnd2s1 U5660 ( .DIN1(n5305), .DIN2(n5518), .Q(n5517) );
  nnd2s1 U5661 ( .DIN1(n5519), .DIN2(n5520), .Q(n5514) );
  nnd2s1 U5662 ( .DIN1(n5301), .DIN2(n5521), .Q(n5520) );
  nnd2s1 U5663 ( .DIN1(n5497), .DIN2(n5522), .Q(n5513) );
  nnd2s1 U5664 ( .DIN1(n5523), .DIN2(n5524), .Q(n5522) );
  nnd2s1 U5665 ( .DIN1(n5525), .DIN2(n5526), .Q(n5512) );
  nnd3s1 U5666 ( .DIN1(n5527), .DIN2(n5305), .DIN3(n5528), .Q(n5526) );
  nnd4s1 U5667 ( .DIN1(n5529), .DIN2(n5530), .DIN3(n5531), .DIN4(n5532), 
        .Q(n5488) );
  nnd2s1 U5668 ( .DIN1(n5533), .DIN2(n5534), .Q(n5532) );
  nnd2s1 U5669 ( .DIN1(n5510), .DIN2(n5535), .Q(n5531) );
  nnd2s1 U5670 ( .DIN1(n5536), .DIN2(n5537), .Q(n5530) );
  nnd2s1 U5671 ( .DIN1(n5511), .DIN2(n5284), .Q(n5529) );
  nnd4s1 U5672 ( .DIN1(n5538), .DIN2(n5539), .DIN3(n5540), .DIN4(n5541), 
        .Q(n5487) );
  nnd2s1 U5673 ( .DIN1(n5542), .DIN2(n5543), .Q(n5541) );
  nnd2s1 U5674 ( .DIN1(n5302), .DIN2(n5544), .Q(n5543) );
  nnd2s1 U5675 ( .DIN1(n5545), .DIN2(n5546), .Q(n5540) );
  nnd2s1 U5676 ( .DIN1(n5294), .DIN2(n5547), .Q(n5539) );
  nnd2s1 U5677 ( .DIN1(n5548), .DIN2(n5549), .Q(n5547) );
  nnd2s1 U5678 ( .DIN1(n5283), .DIN2(n5550), .Q(n5538) );
  or3s1 U5679 ( .DIN1(n5551), .DIN2(n5552), .DIN3(n5553), .Q(n4965) );
  nnd4s1 U5680 ( .DIN1(n5554), .DIN2(n5555), .DIN3(n5556), .DIN4(n5557), 
        .Q(n5553) );
  and4s1 U5681 ( .DIN1(n5558), .DIN2(n5559), .DIN3(n5560), .DIN4(n5561), 
        .Q(n5557) );
  nnd2s1 U5682 ( .DIN1(n5196), .DIN2(n5562), .Q(n5561) );
  nnd2s1 U5683 ( .DIN1(n5563), .DIN2(n5564), .Q(n5562) );
  nnd2s1 U5684 ( .DIN1(n5565), .DIN2(n5566), .Q(n5560) );
  nnd2s1 U5685 ( .DIN1(n5212), .DIN2(n5390), .Q(n5566) );
  nnd2s1 U5686 ( .DIN1(n5219), .DIN2(n5567), .Q(n5559) );
  nnd2s1 U5687 ( .DIN1(n5568), .DIN2(n5569), .Q(n5558) );
  nnd2s1 U5688 ( .DIN1(n5570), .DIN2(n5571), .Q(n5569) );
  nnd2s1 U5689 ( .DIN1(n5370), .DIN2(n5572), .Q(n5556) );
  nnd2s1 U5690 ( .DIN1(n5197), .DIN2(n5415), .Q(n5555) );
  nnd2s1 U5691 ( .DIN1(n5358), .DIN2(n5397), .Q(n5554) );
  nnd3s1 U5692 ( .DIN1(n5350), .DIN2(n5195), .DIN3(n5573), .Q(n5552) );
  nor4s1 U5693 ( .DIN1(n5574), .DIN2(n5575), .DIN3(n5576), .DIN4(n5577), 
        .Q(n5195) );
  nnd4s1 U5694 ( .DIN1(n5578), .DIN2(n5579), .DIN3(n5580), .DIN4(n5581), 
        .Q(n5577) );
  nnd2s1 U5695 ( .DIN1(n5408), .DIN2(n5582), .Q(n5581) );
  nnd2s1 U5696 ( .DIN1(n5565), .DIN2(n5196), .Q(n5580) );
  nnd2s1 U5697 ( .DIN1(n5214), .DIN2(n5359), .Q(n5579) );
  nnd2s1 U5698 ( .DIN1(n5385), .DIN2(n5583), .Q(n5578) );
  nnd3s1 U5699 ( .DIN1(n5584), .DIN2(n5585), .DIN3(n5586), .Q(n5576) );
  nnd2s1 U5700 ( .DIN1(n5388), .DIN2(n5587), .Q(n5586) );
  nnd2s1 U5701 ( .DIN1(n5588), .DIN2(n5589), .Q(n5587) );
  nnd2s1 U5702 ( .DIN1(n5414), .DIN2(n5590), .Q(n5585) );
  nnd2s1 U5703 ( .DIN1(n5591), .DIN2(n5592), .Q(n5590) );
  nnd2s1 U5704 ( .DIN1(n5366), .DIN2(n5593), .Q(n5584) );
  nnd2s1 U5705 ( .DIN1(n5594), .DIN2(n5410), .Q(n5593) );
  nor2s1 U5706 ( .DIN1(n5387), .DIN2(n5595), .Q(n5575) );
  and2s1 U5707 ( .DIN1(n5372), .DIN2(n5596), .Q(n5574) );
  nnd3s1 U5708 ( .DIN1(n5212), .DIN2(n5597), .DIN3(n5222), .Q(n5596) );
  nor3s1 U5709 ( .DIN1(n5598), .DIN2(n5599), .DIN3(n5600), .Q(n5350) );
  nnd4s1 U5710 ( .DIN1(n5193), .DIN2(n5601), .DIN3(n5602), .DIN4(n5603), 
        .Q(n5600) );
  and3s1 U5711 ( .DIN1(n5604), .DIN2(n5605), .DIN3(n5606), .Q(n5603) );
  nnd2s1 U5712 ( .DIN1(n5359), .DIN2(n5357), .Q(n5605) );
  nnd2s1 U5713 ( .DIN1(n5408), .DIN2(n5358), .Q(n5604) );
  nor2s1 U5714 ( .DIN1(n5607), .DIN2(n5608), .Q(n5193) );
  nnd4s1 U5715 ( .DIN1(n5609), .DIN2(n5610), .DIN3(n5611), .DIN4(n5612), 
        .Q(n5608) );
  nnd2s1 U5716 ( .DIN1(n5210), .DIN2(n5613), .Q(n5612) );
  nnd2s1 U5717 ( .DIN1(n5205), .DIN2(n5614), .Q(n5611) );
  nnd2s1 U5718 ( .DIN1(n5565), .DIN2(n5572), .Q(n5610) );
  nnd2s1 U5719 ( .DIN1(n5366), .DIN2(n5378), .Q(n5609) );
  nnd4s1 U5720 ( .DIN1(n5615), .DIN2(n5616), .DIN3(n5617), .DIN4(n5618), 
        .Q(n5607) );
  nnd2s1 U5721 ( .DIN1(n5398), .DIN2(n5619), .Q(n5618) );
  nnd2s1 U5722 ( .DIN1(n5563), .DIN2(n5571), .Q(n5619) );
  nnd2s1 U5723 ( .DIN1(n5196), .DIN2(n5614), .Q(n5617) );
  nnd2s1 U5724 ( .DIN1(n5388), .DIN2(n5620), .Q(n5616) );
  nnd2s1 U5725 ( .DIN1(n5221), .DIN2(n5387), .Q(n5620) );
  nnd2s1 U5726 ( .DIN1(n5621), .DIN2(n5622), .Q(n5615) );
  nnd3s1 U5727 ( .DIN1(n5623), .DIN2(n5395), .DIN3(n5564), .Q(n5622) );
  nnd3s1 U5728 ( .DIN1(n5624), .DIN2(n5625), .DIN3(n5626), .Q(n5599) );
  nnd2s1 U5729 ( .DIN1(n5627), .DIN2(n5373), .Q(n5626) );
  nnd2s1 U5730 ( .DIN1(n5398), .DIN2(n5628), .Q(n5625) );
  nnd3s1 U5731 ( .DIN1(n5384), .DIN2(n5629), .DIN3(n5204), .Q(n5628) );
  nor2s1 U5732 ( .DIN1(n5214), .DIN2(n5405), .Q(n5204) );
  nnd2s1 U5733 ( .DIN1(n5621), .DIN2(n5214), .Q(n5624) );
  nnd3s1 U5734 ( .DIN1(n5630), .DIN2(n5631), .DIN3(n5632), .Q(n5598) );
  nnd2s1 U5735 ( .DIN1(n5210), .DIN2(n5633), .Q(n5632) );
  nnd2s1 U5736 ( .DIN1(n5634), .DIN2(n5203), .Q(n5633) );
  nnd2s1 U5737 ( .DIN1(n5414), .DIN2(n5635), .Q(n5631) );
  nnd2s1 U5738 ( .DIN1(n5410), .DIN2(n5589), .Q(n5635) );
  nnd2s1 U5739 ( .DIN1(n5197), .DIN2(n5636), .Q(n5630) );
  nnd2s1 U5740 ( .DIN1(n5387), .DIN2(n5589), .Q(n5636) );
  nnd3s1 U5741 ( .DIN1(n5637), .DIN2(n5638), .DIN3(n5639), .Q(n5551) );
  xor2s1 U5742 ( .DIN1(n4871), .DIN2(n5640), .Q(n5429) );
  xor2s1 U5743 ( .DIN1(n1375), .DIN2(n4901), .Q(n5640) );
  or3s1 U5744 ( .DIN1(n5641), .DIN2(n5642), .DIN3(n5643), .Q(n4871) );
  nnd4s1 U5745 ( .DIN1(n5644), .DIN2(n5321), .DIN3(n5645), .DIN4(n5646), 
        .Q(n5643) );
  and4s1 U5746 ( .DIN1(n5647), .DIN2(n5648), .DIN3(n5649), .DIN4(n5181), 
        .Q(n5646) );
  nnd2s1 U5747 ( .DIN1(n5650), .DIN2(n5339), .Q(n5181) );
  nnd2s1 U5748 ( .DIN1(n5335), .DIN2(n5651), .Q(n5649) );
  nnd2s1 U5749 ( .DIN1(n5652), .DIN2(n5185), .Q(n5648) );
  nor2s1 U5750 ( .DIN1(n5653), .DIN2(n5654), .Q(n5321) );
  nnd4s1 U5751 ( .DIN1(n5655), .DIN2(n5656), .DIN3(n5657), .DIN4(n5658), 
        .Q(n5654) );
  or2s1 U5752 ( .DIN1(n5659), .DIN2(n5660), .Q(n5658) );
  nnd2s1 U5753 ( .DIN1(n5652), .DIN2(n5661), .Q(n5657) );
  nnd2s1 U5754 ( .DIN1(n5650), .DIN2(n5183), .Q(n5656) );
  nnd2s1 U5755 ( .DIN1(n5156), .DIN2(n5662), .Q(n5655) );
  nnd4s1 U5756 ( .DIN1(n5663), .DIN2(n5664), .DIN3(n5665), .DIN4(n5666), 
        .Q(n5653) );
  nnd2s1 U5757 ( .DIN1(n5155), .DIN2(n5667), .Q(n5666) );
  nnd2s1 U5758 ( .DIN1(n5341), .DIN2(n5668), .Q(n5667) );
  nnd2s1 U5759 ( .DIN1(n5669), .DIN2(n5670), .Q(n5665) );
  nnd2s1 U5760 ( .DIN1(n5337), .DIN2(n5671), .Q(n5670) );
  nnd2s1 U5761 ( .DIN1(n5651), .DIN2(n5672), .Q(n5664) );
  nnd2s1 U5762 ( .DIN1(n5673), .DIN2(n5674), .Q(n5672) );
  nnd2s1 U5763 ( .DIN1(n5165), .DIN2(n5675), .Q(n5663) );
  nnd3s1 U5764 ( .DIN1(n5341), .DIN2(n5676), .DIN3(n5677), .Q(n5675) );
  nnd4s1 U5765 ( .DIN1(n5678), .DIN2(n5679), .DIN3(n5680), .DIN4(n5681), 
        .Q(n5642) );
  nnd2s1 U5766 ( .DIN1(n5682), .DIN2(n5683), .Q(n5681) );
  nnd2s1 U5767 ( .DIN1(n5156), .DIN2(n5684), .Q(n5680) );
  nnd2s1 U5768 ( .DIN1(n5182), .DIN2(n5685), .Q(n5679) );
  nnd2s1 U5769 ( .DIN1(n5323), .DIN2(n5662), .Q(n5678) );
  nnd4s1 U5770 ( .DIN1(n5686), .DIN2(n5687), .DIN3(n5688), .DIN4(n5689), 
        .Q(n5641) );
  nnd2s1 U5771 ( .DIN1(n5173), .DIN2(n5690), .Q(n5689) );
  nnd2s1 U5772 ( .DIN1(n5338), .DIN2(n5691), .Q(n5690) );
  nnd2s1 U5773 ( .DIN1(n5692), .DIN2(n5693), .Q(n5688) );
  nnd2s1 U5774 ( .DIN1(n5169), .DIN2(n5694), .Q(n5687) );
  nnd2s1 U5775 ( .DIN1(n5695), .DIN2(n5164), .Q(n5694) );
  nnd2s1 U5776 ( .DIN1(n5153), .DIN2(n5696), .Q(n5686) );
  nnd2s1 U5777 ( .DIN1(n5697), .DIN2(n1605), .Q(n5426) );
  xor2s1 U5778 ( .DIN1(w3[5]), .DIN2(text_in_r[5]), .Q(n5697) );
  xor2s1 U5779 ( .DIN1(w1[28]), .DIN2(n5698), .Q(N389) );
  xor2s1 U5780 ( .DIN1(n1485), .DIN2(n5699), .Q(N388) );
  xor2s1 U5781 ( .DIN1(n5700), .DIN2(w1[30]), .Q(N387) );
  xor2s1 U5782 ( .DIN1(w1[31]), .DIN2(n5701), .Q(N386) );
  xor2s1 U5783 ( .DIN1(n1481), .DIN2(n5702), .Q(N385) );
  xor2s1 U5784 ( .DIN1(n5703), .DIN2(w0[25]), .Q(N384) );
  xor2s1 U5785 ( .DIN1(w0[26]), .DIN2(n5704), .Q(N383) );
  xor2s1 U5786 ( .DIN1(n5705), .DIN2(w0[27]), .Q(N382) );
  xor2s1 U5787 ( .DIN1(w0[28]), .DIN2(n5706), .Q(N381) );
  xor2s1 U5788 ( .DIN1(n1480), .DIN2(n5707), .Q(N380) );
  nnd2s1 U5789 ( .DIN1(n5708), .DIN2(n5709), .Q(N38) );
  nnd2s1 U5790 ( .DIN1(n5710), .DIN2(n1615), .Q(n5709) );
  xor2s1 U5791 ( .DIN1(n5711), .DIN2(n5712), .Q(n5710) );
  xor2s1 U5792 ( .DIN1(n5713), .DIN2(n5714), .Q(n5712) );
  xnr2s1 U5793 ( .DIN1(n4973), .DIN2(n4780), .Q(n5714) );
  xor2s1 U5794 ( .DIN1(n4901), .DIN2(n4891), .Q(n4780) );
  or3s1 U5795 ( .DIN1(n5715), .DIN2(n5716), .DIN3(n5717), .Q(n4891) );
  nnd4s1 U5796 ( .DIN1(n5434), .DIN2(n5248), .DIN3(n5718), .DIN4(n5719), 
        .Q(n5717) );
  and3s1 U5797 ( .DIN1(n5720), .DIN2(n5721), .DIN3(n5722), .Q(n5719) );
  nor4s1 U5798 ( .DIN1(n5723), .DIN2(n5724), .DIN3(n5725), .DIN4(n5726), 
        .Q(n5248) );
  nnd4s1 U5799 ( .DIN1(n5727), .DIN2(n5728), .DIN3(n5729), .DIN4(n5730), 
        .Q(n5726) );
  nnd2s1 U5800 ( .DIN1(n5106), .DIN2(n5249), .Q(n5730) );
  nnd2s1 U5801 ( .DIN1(n5442), .DIN2(n5731), .Q(n5728) );
  nnd2s1 U5802 ( .DIN1(n5459), .DIN2(n5107), .Q(n5727) );
  nnd3s1 U5803 ( .DIN1(n5732), .DIN2(n5733), .DIN3(n5734), .Q(n5725) );
  nnd2s1 U5804 ( .DIN1(n5472), .DIN2(n5735), .Q(n5734) );
  nnd2s1 U5805 ( .DIN1(n5736), .DIN2(n5122), .Q(n5735) );
  nnd2s1 U5806 ( .DIN1(n5120), .DIN2(n5737), .Q(n5733) );
  nnd2s1 U5807 ( .DIN1(n5738), .DIN2(n5481), .Q(n5737) );
  nnd2s1 U5808 ( .DIN1(n5440), .DIN2(n5739), .Q(n5732) );
  nnd2s1 U5809 ( .DIN1(n5740), .DIN2(n5119), .Q(n5739) );
  nor2s1 U5810 ( .DIN1(n5741), .DIN2(n5742), .Q(n5724) );
  and2s1 U5811 ( .DIN1(n5138), .DIN2(n5743), .Q(n5723) );
  nnd3s1 U5812 ( .DIN1(n5744), .DIN2(n5264), .DIN3(n5267), .Q(n5743) );
  nor3s1 U5813 ( .DIN1(n5745), .DIN2(n5746), .DIN3(n5747), .Q(n5434) );
  nnd4s1 U5814 ( .DIN1(n5246), .DIN2(n5748), .DIN3(n5749), .DIN4(n5750), 
        .Q(n5747) );
  and3s1 U5815 ( .DIN1(n5751), .DIN2(n5752), .DIN3(n5753), .Q(n5750) );
  nnd2s1 U5816 ( .DIN1(n5440), .DIN2(n5452), .Q(n5753) );
  nnd2s1 U5817 ( .DIN1(n5754), .DIN2(n5139), .Q(n5752) );
  nnd2s1 U5818 ( .DIN1(n5755), .DIN2(n5111), .Q(n5751) );
  nor2s1 U5819 ( .DIN1(n5756), .DIN2(n5757), .Q(n5246) );
  nnd4s1 U5820 ( .DIN1(n5758), .DIN2(n5759), .DIN3(n5760), .DIN4(n5761), 
        .Q(n5757) );
  nnd2s1 U5821 ( .DIN1(n5261), .DIN2(n5762), .Q(n5761) );
  nnd2s1 U5822 ( .DIN1(n5124), .DIN2(n5763), .Q(n5760) );
  nnd2s1 U5823 ( .DIN1(n5106), .DIN2(n5764), .Q(n5759) );
  nnd2s1 U5824 ( .DIN1(n5120), .DIN2(n5250), .Q(n5758) );
  nnd4s1 U5825 ( .DIN1(n5765), .DIN2(n5766), .DIN3(n5767), .DIN4(n5768), 
        .Q(n5756) );
  nnd2s1 U5826 ( .DIN1(n5249), .DIN2(n5763), .Q(n5768) );
  nnd2s1 U5827 ( .DIN1(n5110), .DIN2(n5769), .Q(n5767) );
  nnd2s1 U5828 ( .DIN1(n5268), .DIN2(n5461), .Q(n5769) );
  nnd2s1 U5829 ( .DIN1(n5137), .DIN2(n5770), .Q(n5766) );
  nnd2s1 U5830 ( .DIN1(n5771), .DIN2(n5772), .Q(n5770) );
  nnd2s1 U5831 ( .DIN1(n5754), .DIN2(n5773), .Q(n5765) );
  nnd3s1 U5832 ( .DIN1(n5127), .DIN2(n5774), .DIN3(n5775), .Q(n5773) );
  nnd3s1 U5833 ( .DIN1(n5776), .DIN2(n5777), .DIN3(n5102), .Q(n5746) );
  nnd2s1 U5834 ( .DIN1(n5459), .DIN2(n5451), .Q(n5102) );
  nnd2s1 U5835 ( .DIN1(n5137), .DIN2(n5778), .Q(n5777) );
  nnd3s1 U5836 ( .DIN1(n5464), .DIN2(n5779), .DIN3(n5256), .Q(n5778) );
  nor2s1 U5837 ( .DIN1(n5482), .DIN2(n5139), .Q(n5256) );
  nnd2s1 U5838 ( .DIN1(n5441), .DIN2(n5128), .Q(n5776) );
  nnd3s1 U5839 ( .DIN1(n5780), .DIN2(n5781), .DIN3(n5782), .Q(n5745) );
  nnd2s1 U5840 ( .DIN1(n5472), .DIN2(n5783), .Q(n5782) );
  nnd2s1 U5841 ( .DIN1(n5449), .DIN2(n5481), .Q(n5783) );
  nnd2s1 U5842 ( .DIN1(n5108), .DIN2(n5784), .Q(n5781) );
  nnd2s1 U5843 ( .DIN1(n5461), .DIN2(n5449), .Q(n5784) );
  nnd2s1 U5844 ( .DIN1(n5261), .DIN2(n5785), .Q(n5780) );
  nnd2s1 U5845 ( .DIN1(n5738), .DIN2(n5268), .Q(n5785) );
  nnd3s1 U5846 ( .DIN1(n5786), .DIN2(n5787), .DIN3(n5788), .Q(n5716) );
  nnd2s1 U5847 ( .DIN1(n5442), .DIN2(n5764), .Q(n5788) );
  nnd2s1 U5848 ( .DIN1(n5108), .DIN2(n5473), .Q(n5787) );
  nnd2s1 U5849 ( .DIN1(n5441), .DIN2(n5474), .Q(n5786) );
  nnd4s1 U5850 ( .DIN1(n5789), .DIN2(n5790), .DIN3(n5791), .DIN4(n5792), 
        .Q(n5715) );
  nnd2s1 U5851 ( .DIN1(n5106), .DIN2(n5793), .Q(n5792) );
  nnd2s1 U5852 ( .DIN1(n5458), .DIN2(n5264), .Q(n5793) );
  nnd2s1 U5853 ( .DIN1(n5249), .DIN2(n5794), .Q(n5791) );
  nnd2s1 U5854 ( .DIN1(n5775), .DIN2(n5771), .Q(n5794) );
  nnd2s1 U5855 ( .DIN1(n5265), .DIN2(n5795), .Q(n5790) );
  nnd2s1 U5856 ( .DIN1(n5116), .DIN2(n5796), .Q(n5789) );
  nnd2s1 U5857 ( .DIN1(n5797), .DIN2(n5772), .Q(n5796) );
  or3s1 U5858 ( .DIN1(n5798), .DIN2(n5799), .DIN3(n5800), .Q(n4901) );
  nnd4s1 U5859 ( .DIN1(n5490), .DIN2(n5282), .DIN3(n5801), .DIN4(n5802), 
        .Q(n5800) );
  and3s1 U5860 ( .DIN1(n5803), .DIN2(n5804), .DIN3(n5805), .Q(n5802) );
  nor4s1 U5861 ( .DIN1(n5806), .DIN2(n5807), .DIN3(n5808), .DIN4(n5809), 
        .Q(n5282) );
  nnd4s1 U5862 ( .DIN1(n5810), .DIN2(n5811), .DIN3(n5812), .DIN4(n5813), 
        .Q(n5809) );
  nnd2s1 U5863 ( .DIN1(n5284), .DIN2(n5814), .Q(n5813) );
  nnd2s1 U5864 ( .DIN1(n5499), .DIN2(n5815), .Q(n5811) );
  nnd2s1 U5865 ( .DIN1(n5816), .DIN2(n5519), .Q(n5810) );
  nnd3s1 U5866 ( .DIN1(n5817), .DIN2(n5818), .DIN3(n5819), .Q(n5808) );
  nnd2s1 U5867 ( .DIN1(n5533), .DIN2(n5820), .Q(n5819) );
  nnd2s1 U5868 ( .DIN1(n5821), .DIN2(n5822), .Q(n5820) );
  nnd2s1 U5869 ( .DIN1(n5525), .DIN2(n5823), .Q(n5818) );
  nnd2s1 U5870 ( .DIN1(n5824), .DIN2(n5544), .Q(n5823) );
  nnd2s1 U5871 ( .DIN1(n5509), .DIN2(n5825), .Q(n5817) );
  nnd2s1 U5872 ( .DIN1(n5826), .DIN2(n5549), .Q(n5825) );
  nor2s1 U5873 ( .DIN1(n5827), .DIN2(n5828), .Q(n5807) );
  and2s1 U5874 ( .DIN1(n5286), .DIN2(n5829), .Q(n5806) );
  nnd3s1 U5875 ( .DIN1(n5302), .DIN2(n5305), .DIN3(n5830), .Q(n5829) );
  nor3s1 U5876 ( .DIN1(n5831), .DIN2(n5832), .DIN3(n5833), .Q(n5490) );
  nnd4s1 U5877 ( .DIN1(n5280), .DIN2(n5834), .DIN3(n5835), .DIN4(n5836), 
        .Q(n5833) );
  and3s1 U5878 ( .DIN1(n5837), .DIN2(n5838), .DIN3(n5839), .Q(n5836) );
  nnd2s1 U5879 ( .DIN1(n5511), .DIN2(n5509), .Q(n5839) );
  nnd2s1 U5880 ( .DIN1(n5307), .DIN2(n5840), .Q(n5838) );
  nnd2s1 U5881 ( .DIN1(n5841), .DIN2(n5510), .Q(n5837) );
  nor2s1 U5882 ( .DIN1(n5842), .DIN2(n5843), .Q(n5280) );
  nnd4s1 U5883 ( .DIN1(n5844), .DIN2(n5845), .DIN3(n5846), .DIN4(n5847), 
        .Q(n5843) );
  nnd2s1 U5884 ( .DIN1(n5299), .DIN2(n5848), .Q(n5847) );
  nnd2s1 U5885 ( .DIN1(n5294), .DIN2(n5849), .Q(n5846) );
  nnd2s1 U5886 ( .DIN1(n5814), .DIN2(n5850), .Q(n5845) );
  nnd2s1 U5887 ( .DIN1(n5285), .DIN2(n5525), .Q(n5844) );
  nnd4s1 U5888 ( .DIN1(n5851), .DIN2(n5852), .DIN3(n5853), .DIN4(n5854), 
        .Q(n5842) );
  nnd2s1 U5889 ( .DIN1(n5284), .DIN2(n5849), .Q(n5854) );
  nnd2s1 U5890 ( .DIN1(n5516), .DIN2(n5855), .Q(n5853) );
  nnd2s1 U5891 ( .DIN1(n5306), .DIN2(n5521), .Q(n5855) );
  nnd2s1 U5892 ( .DIN1(n5537), .DIN2(n5856), .Q(n5852) );
  nnd2s1 U5893 ( .DIN1(n5857), .DIN2(n5858), .Q(n5856) );
  nnd2s1 U5894 ( .DIN1(n5840), .DIN2(n5859), .Q(n5851) );
  nnd3s1 U5895 ( .DIN1(n5860), .DIN2(n5861), .DIN3(n5862), .Q(n5859) );
  nnd3s1 U5896 ( .DIN1(n5863), .DIN2(n5864), .DIN3(n5865), .Q(n5832) );
  nnd2s1 U5897 ( .DIN1(n5537), .DIN2(n5866), .Q(n5864) );
  nnd3s1 U5898 ( .DIN1(n5524), .DIN2(n5867), .DIN3(n5293), .Q(n5866) );
  nor2s1 U5899 ( .DIN1(n5545), .DIN2(n5307), .Q(n5293) );
  nnd2s1 U5900 ( .DIN1(n5497), .DIN2(n5542), .Q(n5863) );
  nnd3s1 U5901 ( .DIN1(n5868), .DIN2(n5869), .DIN3(n5870), .Q(n5831) );
  nnd2s1 U5902 ( .DIN1(n5533), .DIN2(n5871), .Q(n5870) );
  nnd2s1 U5903 ( .DIN1(n5506), .DIN2(n5544), .Q(n5871) );
  nnd2s1 U5904 ( .DIN1(n5283), .DIN2(n5872), .Q(n5869) );
  nnd2s1 U5905 ( .DIN1(n5521), .DIN2(n5506), .Q(n5872) );
  nnd2s1 U5906 ( .DIN1(n5299), .DIN2(n5873), .Q(n5868) );
  nnd2s1 U5907 ( .DIN1(n5824), .DIN2(n5306), .Q(n5873) );
  nnd3s1 U5908 ( .DIN1(n5874), .DIN2(n5875), .DIN3(n5876), .Q(n5799) );
  nnd2s1 U5909 ( .DIN1(n5499), .DIN2(n5850), .Q(n5876) );
  nnd2s1 U5910 ( .DIN1(n5283), .DIN2(n5534), .Q(n5875) );
  nnd2s1 U5911 ( .DIN1(n5497), .DIN2(n5535), .Q(n5874) );
  nnd4s1 U5912 ( .DIN1(n5877), .DIN2(n5878), .DIN3(n5879), .DIN4(n5880), 
        .Q(n5798) );
  nnd2s1 U5913 ( .DIN1(n5814), .DIN2(n5881), .Q(n5880) );
  nnd2s1 U5914 ( .DIN1(n5518), .DIN2(n5302), .Q(n5881) );
  nnd2s1 U5915 ( .DIN1(n5284), .DIN2(n5882), .Q(n5879) );
  nnd2s1 U5916 ( .DIN1(n5862), .DIN2(n5857), .Q(n5882) );
  nnd2s1 U5917 ( .DIN1(n5303), .DIN2(n5883), .Q(n5878) );
  nnd2s1 U5918 ( .DIN1(n5884), .DIN2(n5885), .Q(n5877) );
  nnd2s1 U5919 ( .DIN1(n5886), .DIN2(n5858), .Q(n5885) );
  or3s1 U5920 ( .DIN1(n5887), .DIN2(n5888), .DIN3(n5889), .Q(n4973) );
  nnd4s1 U5921 ( .DIN1(n5890), .DIN2(n5891), .DIN3(n5191), .DIN4(n5892), 
        .Q(n5889) );
  and3s1 U5922 ( .DIN1(n5351), .DIN2(n5602), .DIN3(n5573), .Q(n5892) );
  nor4s1 U5923 ( .DIN1(n5893), .DIN2(n5894), .DIN3(n5895), .DIN4(n5896), 
        .Q(n5573) );
  nnd4s1 U5924 ( .DIN1(n5897), .DIN2(n5898), .DIN3(n5899), .DIN4(n5900), 
        .Q(n5896) );
  nor2s1 U5925 ( .DIN1(n5901), .DIN2(n5902), .Q(n5900) );
  nor2s1 U5926 ( .DIN1(n5903), .DIN2(n5201), .Q(n5902) );
  nor2s1 U5927 ( .DIN1(n5563), .DIN2(n5904), .Q(n5901) );
  nnd2s1 U5928 ( .DIN1(n5400), .DIN2(n5357), .Q(n5899) );
  nnd2s1 U5929 ( .DIN1(n5414), .DIN2(n5371), .Q(n5898) );
  nnd2s1 U5930 ( .DIN1(n5565), .DIN2(n5378), .Q(n5897) );
  nnd3s1 U5931 ( .DIN1(n5905), .DIN2(n5906), .DIN3(n5907), .Q(n5895) );
  or2s1 U5932 ( .DIN1(n5588), .DIN2(n5908), .Q(n5907) );
  nnd2s1 U5933 ( .DIN1(n5627), .DIN2(n5909), .Q(n5906) );
  nnd3s1 U5934 ( .DIN1(n5589), .DIN2(n5203), .DIN3(n5213), .Q(n5909) );
  nnd2s1 U5935 ( .DIN1(n5910), .DIN2(n5911), .Q(n5905) );
  nnd3s1 U5936 ( .DIN1(n5380), .DIN2(n5395), .DIN3(n5912), .Q(n5911) );
  nor2s1 U5937 ( .DIN1(n5410), .DIN2(n5595), .Q(n5894) );
  nor2s1 U5938 ( .DIN1(n5396), .DIN2(n5564), .Q(n5893) );
  nor4s1 U5939 ( .DIN1(n5913), .DIN2(n5914), .DIN3(n5915), .DIN4(n5916), 
        .Q(n5602) );
  nnd4s1 U5940 ( .DIN1(n5917), .DIN2(n5918), .DIN3(n5919), .DIN4(n5920), 
        .Q(n5916) );
  nnd2s1 U5941 ( .DIN1(n5372), .DIN2(n5583), .Q(n5920) );
  nor2s1 U5942 ( .DIN1(n5921), .DIN2(n5922), .Q(n5919) );
  nor2s1 U5943 ( .DIN1(n5912), .DIN2(n5588), .Q(n5922) );
  nor2s1 U5944 ( .DIN1(n5390), .DIN2(n5595), .Q(n5921) );
  nnd2s1 U5945 ( .DIN1(n5408), .DIN2(n5378), .Q(n5918) );
  nnd2s1 U5946 ( .DIN1(n5197), .DIN2(n5358), .Q(n5917) );
  nnd3s1 U5947 ( .DIN1(n5923), .DIN2(n5924), .DIN3(n5925), .Q(n5915) );
  nnd2s1 U5948 ( .DIN1(n5196), .DIN2(n5926), .Q(n5925) );
  nnd2s1 U5949 ( .DIN1(n5570), .DIN2(n5380), .Q(n5926) );
  nnd2s1 U5950 ( .DIN1(n5357), .DIN2(n5927), .Q(n5924) );
  nnd2s1 U5951 ( .DIN1(n5928), .DIN2(n5589), .Q(n5927) );
  nnd2s1 U5952 ( .DIN1(n5400), .DIN2(n5929), .Q(n5923) );
  nnd2s1 U5953 ( .DIN1(n5629), .DIN2(n5413), .Q(n5929) );
  nor2s1 U5954 ( .DIN1(n5930), .DIN2(n5412), .Q(n5914) );
  nor2s1 U5955 ( .DIN1(n5582), .DIN2(n5568), .Q(n5930) );
  nor2s1 U5956 ( .DIN1(n5931), .DIN2(n5212), .Q(n5913) );
  nor2s1 U5957 ( .DIN1(n5627), .DIN2(n5405), .Q(n5931) );
  nor4s1 U5958 ( .DIN1(n5932), .DIN2(n5933), .DIN3(n5934), .DIN4(n5935), 
        .Q(n5351) );
  nnd4s1 U5959 ( .DIN1(n5936), .DIN2(n5937), .DIN3(n5938), .DIN4(n5939), 
        .Q(n5935) );
  nor2s1 U5960 ( .DIN1(n5940), .DIN2(n5941), .Q(n5938) );
  nor2s1 U5961 ( .DIN1(n5571), .DIN2(n5222), .Q(n5941) );
  nor2s1 U5962 ( .DIN1(n5368), .DIN2(n5595), .Q(n5940) );
  nnd2s1 U5963 ( .DIN1(n5565), .DIN2(n5583), .Q(n5937) );
  nnd2s1 U5964 ( .DIN1(n5359), .DIN2(n5385), .Q(n5936) );
  nnd3s1 U5965 ( .DIN1(n5942), .DIN2(n5943), .DIN3(n5944), .Q(n5934) );
  nnd2s1 U5966 ( .DIN1(n5197), .DIN2(n5945), .Q(n5944) );
  nnd2s1 U5967 ( .DIN1(n5205), .DIN2(n5946), .Q(n5943) );
  nnd2s1 U5968 ( .DIN1(n5380), .DIN2(n5571), .Q(n5946) );
  nnd2s1 U5969 ( .DIN1(n5627), .DIN2(n5947), .Q(n5942) );
  nnd3s1 U5970 ( .DIN1(n5588), .DIN2(n5597), .DIN3(n5948), .Q(n5947) );
  nor2s1 U5971 ( .DIN1(n5381), .DIN2(n5221), .Q(n5933) );
  nor2s1 U5972 ( .DIN1(n5216), .DIN2(n5412), .Q(n5932) );
  nor3s1 U5973 ( .DIN1(n5949), .DIN2(n5950), .DIN3(n5951), .Q(n5191) );
  nnd4s1 U5974 ( .DIN1(n5601), .DIN2(n5353), .DIN3(n5639), .DIN4(n5952), 
        .Q(n5951) );
  and3s1 U5975 ( .DIN1(n5953), .DIN2(n5954), .DIN3(n5955), .Q(n5952) );
  nnd2s1 U5976 ( .DIN1(n5197), .DIN2(n5568), .Q(n5955) );
  nnd2s1 U5977 ( .DIN1(n5370), .DIN2(n5583), .Q(n5954) );
  nnd2s1 U5978 ( .DIN1(n5398), .DIN2(n5219), .Q(n5953) );
  nor4s1 U5979 ( .DIN1(n5956), .DIN2(n5957), .DIN3(n5958), .DIN4(n5959), 
        .Q(n5639) );
  nnd4s1 U5980 ( .DIN1(n5960), .DIN2(n5961), .DIN3(n5962), .DIN4(n5963), 
        .Q(n5959) );
  nnd2s1 U5981 ( .DIN1(n5219), .DIN2(n5964), .Q(n5963) );
  nor2s1 U5982 ( .DIN1(n5965), .DIN2(n5966), .Q(n5962) );
  nor2s1 U5983 ( .DIN1(n5967), .DIN2(n5597), .Q(n5966) );
  nor2s1 U5984 ( .DIN1(n5370), .DIN2(n5565), .Q(n5967) );
  nor2s1 U5985 ( .DIN1(n5968), .DIN2(n5413), .Q(n5965) );
  nor2s1 U5986 ( .DIN1(n5398), .DIN2(n5218), .Q(n5968) );
  nnd2s1 U5987 ( .DIN1(n5568), .DIN2(n5969), .Q(n5961) );
  nnd3s1 U5988 ( .DIN1(n5623), .DIN2(n5563), .DIN3(n5381), .Q(n5969) );
  nnd2s1 U5989 ( .DIN1(n5970), .DIN2(n5405), .Q(n5960) );
  nnd3s1 U5990 ( .DIN1(n5971), .DIN2(n5972), .DIN3(n5973), .Q(n5958) );
  nnd2s1 U5991 ( .DIN1(n5627), .DIN2(n5582), .Q(n5973) );
  nnd2s1 U5992 ( .DIN1(n5400), .DIN2(n5414), .Q(n5971) );
  nor2s1 U5993 ( .DIN1(n5588), .DIN2(n5570), .Q(n5957) );
  nor2s1 U5994 ( .DIN1(n5410), .DIN2(n5412), .Q(n5956) );
  nor4s1 U5995 ( .DIN1(n5974), .DIN2(n5975), .DIN3(n5976), .DIN4(n5977), 
        .Q(n5353) );
  nnd4s1 U5996 ( .DIN1(n5978), .DIN2(n5979), .DIN3(n5980), .DIN4(n5981), 
        .Q(n5977) );
  nnd2s1 U5997 ( .DIN1(n5568), .DIN2(n5414), .Q(n5981) );
  nnd2s1 U5998 ( .DIN1(n5405), .DIN2(n5910), .Q(n5980) );
  nnd2s1 U5999 ( .DIN1(n5408), .DIN2(n5583), .Q(n5979) );
  nnd2s1 U6000 ( .DIN1(n5219), .DIN2(n5371), .Q(n5978) );
  nnd3s1 U6001 ( .DIN1(n5982), .DIN2(n5983), .DIN3(n5984), .Q(n5976) );
  nnd2s1 U6002 ( .DIN1(n5214), .DIN2(n5985), .Q(n5984) );
  nnd2s1 U6003 ( .DIN1(n5634), .DIN2(n5387), .Q(n5985) );
  nor2s1 U6004 ( .DIN1(n5400), .DIN2(n5582), .Q(n5634) );
  nnd2s1 U6005 ( .DIN1(n5399), .DIN2(n5986), .Q(n5983) );
  nnd2s1 U6006 ( .DIN1(n5928), .DIN2(n5387), .Q(n5986) );
  nor2s1 U6007 ( .DIN1(n5582), .DIN2(n5970), .Q(n5928) );
  nnd2s1 U6008 ( .DIN1(n5621), .DIN2(n5987), .Q(n5982) );
  nnd2s1 U6009 ( .DIN1(n5570), .DIN2(n5595), .Q(n5987) );
  nor2s1 U6010 ( .DIN1(n5588), .DIN2(n5595), .Q(n5975) );
  nor2s1 U6011 ( .DIN1(n5369), .DIN2(n5571), .Q(n5974) );
  hi1s1 U6012 ( .DIN(n5988), .Q(n5369) );
  nor2s1 U6013 ( .DIN1(n5989), .DIN2(n5990), .Q(n5601) );
  nnd4s1 U6014 ( .DIN1(n5991), .DIN2(n5992), .DIN3(n5993), .DIN4(n5994), 
        .Q(n5990) );
  nnd2s1 U6015 ( .DIN1(n5583), .DIN2(n5995), .Q(n5994) );
  nnd3s1 U6016 ( .DIN1(n5912), .DIN2(n5571), .DIN3(n5381), .Q(n5995) );
  nnd2s1 U6017 ( .DIN1(n5565), .DIN2(n5358), .Q(n5991) );
  nnd4s1 U6018 ( .DIN1(n5996), .DIN2(n5997), .DIN3(n5998), .DIN4(n5999), 
        .Q(n5989) );
  nnd2s1 U6019 ( .DIN1(n5372), .DIN2(n6000), .Q(n5999) );
  nnd2s1 U6020 ( .DIN1(n5621), .DIN2(n6001), .Q(n5998) );
  nnd2s1 U6021 ( .DIN1(n5202), .DIN2(n5563), .Q(n6001) );
  nnd2s1 U6022 ( .DIN1(n5408), .DIN2(n6002), .Q(n5997) );
  nnd2s1 U6023 ( .DIN1(n6003), .DIN2(n5221), .Q(n6002) );
  nnd2s1 U6024 ( .DIN1(n5205), .DIN2(n6004), .Q(n5996) );
  nnd2s1 U6025 ( .DIN1(n5564), .DIN2(n5381), .Q(n6004) );
  nnd3s1 U6026 ( .DIN1(n6005), .DIN2(n6006), .DIN3(n6007), .Q(n5950) );
  nnd2s1 U6027 ( .DIN1(n5366), .DIN2(n5970), .Q(n6007) );
  nnd2s1 U6028 ( .DIN1(n5582), .DIN2(n6008), .Q(n6006) );
  nnd3s1 U6029 ( .DIN1(n5912), .DIN2(n5623), .DIN3(n6009), .Q(n6008) );
  or2s1 U6030 ( .DIN1(n5387), .DIN2(n6010), .Q(n6005) );
  nnd3s1 U6031 ( .DIN1(n6011), .DIN2(n6012), .DIN3(n6013), .Q(n5949) );
  nnd2s1 U6032 ( .DIN1(n5205), .DIN2(n6014), .Q(n6013) );
  nnd2s1 U6033 ( .DIN1(n5395), .DIN2(n5629), .Q(n6014) );
  nnd2s1 U6034 ( .DIN1(n5405), .DIN2(n6015), .Q(n6012) );
  nnd2s1 U6035 ( .DIN1(n5592), .DIN2(n5589), .Q(n6015) );
  nnd2s1 U6036 ( .DIN1(n5385), .DIN2(n6016), .Q(n6011) );
  nnd2s1 U6037 ( .DIN1(n5396), .DIN2(n5597), .Q(n6016) );
  nor2s1 U6038 ( .DIN1(n5373), .DIN2(n5400), .Q(n5396) );
  nnd2s1 U6039 ( .DIN1(n5366), .DIN2(n5359), .Q(n5891) );
  nnd3s1 U6040 ( .DIN1(n6017), .DIN2(n6018), .DIN3(n6019), .Q(n5888) );
  nnd2s1 U6041 ( .DIN1(n5219), .DIN2(n5378), .Q(n6019) );
  nnd2s1 U6042 ( .DIN1(n6020), .DIN2(n6021), .Q(n6018) );
  nnd2s1 U6043 ( .DIN1(n5970), .DIN2(n5408), .Q(n6017) );
  nnd4s1 U6044 ( .DIN1(n6022), .DIN2(n6023), .DIN3(n6024), .DIN4(n6025), 
        .Q(n5887) );
  nnd2s1 U6045 ( .DIN1(n5399), .DIN2(n6026), .Q(n6025) );
  nnd2s1 U6046 ( .DIN1(n5216), .DIN2(n5410), .Q(n6026) );
  nor2s1 U6047 ( .DIN1(n5371), .DIN2(n5358), .Q(n5216) );
  nnd2s1 U6048 ( .DIN1(n5400), .DIN2(n6027), .Q(n6024) );
  nnd2s1 U6049 ( .DIN1(n5623), .DIN2(n5384), .Q(n6027) );
  nnd2s1 U6050 ( .DIN1(n5371), .DIN2(n6028), .Q(n6023) );
  nnd2s1 U6051 ( .DIN1(n5383), .DIN2(n5395), .Q(n6028) );
  nnd2s1 U6052 ( .DIN1(n5568), .DIN2(n5614), .Q(n6022) );
  xor2s1 U6053 ( .DIN1(n4912), .DIN2(n6029), .Q(n5711) );
  xor2s1 U6054 ( .DIN1(n1441), .DIN2(n4889), .Q(n6029) );
  or3s1 U6055 ( .DIN1(n6030), .DIN2(n6031), .DIN3(n6032), .Q(n4889) );
  nnd4s1 U6056 ( .DIN1(n5644), .DIN2(n5322), .DIN3(n6033), .DIN4(n6034), 
        .Q(n6032) );
  and3s1 U6057 ( .DIN1(n6035), .DIN2(n6036), .DIN3(n6037), .Q(n6034) );
  nor4s1 U6058 ( .DIN1(n6038), .DIN2(n6039), .DIN3(n6040), .DIN4(n6041), 
        .Q(n5322) );
  nnd4s1 U6059 ( .DIN1(n6042), .DIN2(n6043), .DIN3(n6044), .DIN4(n6045), 
        .Q(n6041) );
  nnd2s1 U6060 ( .DIN1(n5151), .DIN2(n5323), .Q(n6045) );
  nnd2s1 U6061 ( .DIN1(n5652), .DIN2(n6046), .Q(n6043) );
  nnd2s1 U6062 ( .DIN1(n5669), .DIN2(n5152), .Q(n6042) );
  nnd3s1 U6063 ( .DIN1(n6047), .DIN2(n6048), .DIN3(n6049), .Q(n6040) );
  nnd2s1 U6064 ( .DIN1(n5682), .DIN2(n6050), .Q(n6049) );
  nnd2s1 U6065 ( .DIN1(n6051), .DIN2(n5167), .Q(n6050) );
  nnd2s1 U6066 ( .DIN1(n5165), .DIN2(n6052), .Q(n6048) );
  nnd2s1 U6067 ( .DIN1(n6053), .DIN2(n5691), .Q(n6052) );
  nnd2s1 U6068 ( .DIN1(n5650), .DIN2(n6054), .Q(n6047) );
  nnd2s1 U6069 ( .DIN1(n6055), .DIN2(n5164), .Q(n6054) );
  nor2s1 U6070 ( .DIN1(n6056), .DIN2(n6057), .Q(n6039) );
  and2s1 U6071 ( .DIN1(n5183), .DIN2(n6058), .Q(n6038) );
  nnd3s1 U6072 ( .DIN1(n6059), .DIN2(n5338), .DIN3(n5341), .Q(n6058) );
  nor3s1 U6073 ( .DIN1(n6060), .DIN2(n6061), .DIN3(n6062), .Q(n5644) );
  nnd4s1 U6074 ( .DIN1(n5320), .DIN2(n6063), .DIN3(n6064), .DIN4(n6065), 
        .Q(n6062) );
  and3s1 U6075 ( .DIN1(n6066), .DIN2(n6067), .DIN3(n6068), .Q(n6065) );
  nnd2s1 U6076 ( .DIN1(n5650), .DIN2(n5662), .Q(n6068) );
  nnd2s1 U6077 ( .DIN1(n6069), .DIN2(n5184), .Q(n6067) );
  nnd2s1 U6078 ( .DIN1(n6070), .DIN2(n5156), .Q(n6066) );
  nor2s1 U6079 ( .DIN1(n6071), .DIN2(n6072), .Q(n5320) );
  nnd4s1 U6080 ( .DIN1(n6073), .DIN2(n6074), .DIN3(n6075), .DIN4(n6076), 
        .Q(n6072) );
  nnd2s1 U6081 ( .DIN1(n5335), .DIN2(n6077), .Q(n6076) );
  nnd2s1 U6082 ( .DIN1(n5169), .DIN2(n6078), .Q(n6075) );
  nnd2s1 U6083 ( .DIN1(n5151), .DIN2(n6079), .Q(n6074) );
  nnd2s1 U6084 ( .DIN1(n5165), .DIN2(n5324), .Q(n6073) );
  nnd4s1 U6085 ( .DIN1(n6080), .DIN2(n6081), .DIN3(n6082), .DIN4(n6083), 
        .Q(n6071) );
  nnd2s1 U6086 ( .DIN1(n5323), .DIN2(n6078), .Q(n6083) );
  nnd2s1 U6087 ( .DIN1(n5155), .DIN2(n6084), .Q(n6082) );
  nnd2s1 U6088 ( .DIN1(n5342), .DIN2(n5671), .Q(n6084) );
  nnd2s1 U6089 ( .DIN1(n5182), .DIN2(n6085), .Q(n6081) );
  nnd2s1 U6090 ( .DIN1(n6086), .DIN2(n6087), .Q(n6085) );
  nnd2s1 U6091 ( .DIN1(n6069), .DIN2(n6088), .Q(n6080) );
  nnd3s1 U6092 ( .DIN1(n5172), .DIN2(n6089), .DIN3(n6090), .Q(n6088) );
  nnd3s1 U6093 ( .DIN1(n6091), .DIN2(n6092), .DIN3(n5147), .Q(n6061) );
  nnd2s1 U6094 ( .DIN1(n5669), .DIN2(n5661), .Q(n5147) );
  nnd2s1 U6095 ( .DIN1(n5182), .DIN2(n6093), .Q(n6092) );
  nnd3s1 U6096 ( .DIN1(n5674), .DIN2(n6094), .DIN3(n5330), .Q(n6093) );
  nor2s1 U6097 ( .DIN1(n5692), .DIN2(n5184), .Q(n5330) );
  nnd2s1 U6098 ( .DIN1(n5651), .DIN2(n5173), .Q(n6091) );
  nnd3s1 U6099 ( .DIN1(n6095), .DIN2(n6096), .DIN3(n6097), .Q(n6060) );
  nnd2s1 U6100 ( .DIN1(n5682), .DIN2(n6098), .Q(n6097) );
  nnd2s1 U6101 ( .DIN1(n5659), .DIN2(n5691), .Q(n6098) );
  nnd2s1 U6102 ( .DIN1(n5153), .DIN2(n6099), .Q(n6096) );
  nnd2s1 U6103 ( .DIN1(n5671), .DIN2(n5659), .Q(n6099) );
  nnd2s1 U6104 ( .DIN1(n5335), .DIN2(n6100), .Q(n6095) );
  nnd2s1 U6105 ( .DIN1(n6053), .DIN2(n5342), .Q(n6100) );
  nnd3s1 U6106 ( .DIN1(n6101), .DIN2(n6102), .DIN3(n6103), .Q(n6031) );
  nnd2s1 U6107 ( .DIN1(n5652), .DIN2(n6079), .Q(n6103) );
  nnd2s1 U6108 ( .DIN1(n5153), .DIN2(n5683), .Q(n6102) );
  nnd2s1 U6109 ( .DIN1(n5651), .DIN2(n5684), .Q(n6101) );
  nnd4s1 U6110 ( .DIN1(n6104), .DIN2(n6105), .DIN3(n6106), .DIN4(n6107), 
        .Q(n6030) );
  nnd2s1 U6111 ( .DIN1(n5151), .DIN2(n6108), .Q(n6107) );
  nnd2s1 U6112 ( .DIN1(n5668), .DIN2(n5338), .Q(n6108) );
  nnd2s1 U6113 ( .DIN1(n5323), .DIN2(n6109), .Q(n6106) );
  nnd2s1 U6114 ( .DIN1(n6090), .DIN2(n6086), .Q(n6109) );
  nnd2s1 U6115 ( .DIN1(n5339), .DIN2(n6110), .Q(n6105) );
  nnd2s1 U6116 ( .DIN1(n5161), .DIN2(n6111), .Q(n6104) );
  nnd2s1 U6117 ( .DIN1(n6112), .DIN2(n6087), .Q(n6111) );
  nnd2s1 U6118 ( .DIN1(n6113), .DIN2(n1605), .Q(n5708) );
  xor2s1 U6119 ( .DIN1(w3[4]), .DIN2(text_in_r[4]), .Q(n6113) );
  xor2s1 U6120 ( .DIN1(n6114), .DIN2(w0[30]), .Q(N379) );
  xor2s1 U6121 ( .DIN1(w0[31]), .DIN2(n6115), .Q(N378) );
  nnd2s1 U6122 ( .DIN1(n6116), .DIN2(n6117), .Q(N37) );
  nnd2s1 U6123 ( .DIN1(n6118), .DIN2(n1615), .Q(n6117) );
  xor2s1 U6124 ( .DIN1(n6119), .DIN2(n6120), .Q(n6118) );
  xor2s1 U6125 ( .DIN1(n5713), .DIN2(n6121), .Q(n6120) );
  xor2s1 U6126 ( .DIN1(n4989), .DIN2(n4987), .Q(n6121) );
  xnr2s1 U6127 ( .DIN1(n4912), .DIN2(n4819), .Q(n4987) );
  or3s1 U6128 ( .DIN1(n6122), .DIN2(n6123), .DIN3(n6124), .Q(n4819) );
  nnd4s1 U6129 ( .DIN1(n6125), .DIN2(n6126), .DIN3(n5244), .DIN4(n6127), 
        .Q(n6124) );
  and3s1 U6130 ( .DIN1(n5435), .DIN2(n5749), .DIN3(n5718), .Q(n6127) );
  nor4s1 U6131 ( .DIN1(n6128), .DIN2(n6129), .DIN3(n6130), .DIN4(n6131), 
        .Q(n5718) );
  nnd4s1 U6132 ( .DIN1(n6132), .DIN2(n6133), .DIN3(n6134), .DIN4(n6135), 
        .Q(n6131) );
  nnd2s1 U6133 ( .DIN1(n5111), .DIN2(n5265), .Q(n6135) );
  nor2s1 U6134 ( .DIN1(n6136), .DIN2(n6137), .Q(n6134) );
  nor2s1 U6135 ( .DIN1(n5264), .DIN2(n6138), .Q(n6137) );
  nor2s1 U6136 ( .DIN1(n5481), .DIN2(n6139), .Q(n6136) );
  nnd2s1 U6137 ( .DIN1(n5140), .DIN2(n5452), .Q(n6133) );
  nnd2s1 U6138 ( .DIN1(n5459), .DIN2(n5124), .Q(n6132) );
  nnd3s1 U6139 ( .DIN1(n6140), .DIN2(n6141), .DIN3(n6142), .Q(n6130) );
  nnd2s1 U6140 ( .DIN1(n5482), .DIN2(n5486), .Q(n6142) );
  nnd2s1 U6141 ( .DIN1(n5109), .DIN2(n6143), .Q(n6141) );
  nnd3s1 U6142 ( .DIN1(n5774), .DIN2(n5740), .DIN3(n6138), .Q(n6143) );
  nnd2s1 U6143 ( .DIN1(n5755), .DIN2(n6144), .Q(n6140) );
  nnd3s1 U6144 ( .DIN1(n5449), .DIN2(n5123), .DIN3(n5263), .Q(n6144) );
  nor2s1 U6145 ( .DIN1(n5449), .DIN2(n5127), .Q(n6129) );
  nor2s1 U6146 ( .DIN1(n6145), .DIN2(n6146), .Q(n6128) );
  nor4s1 U6147 ( .DIN1(n6147), .DIN2(n6148), .DIN3(n6149), .DIN4(n6150), 
        .Q(n5749) );
  nnd4s1 U6148 ( .DIN1(n6151), .DIN2(n6152), .DIN3(n6153), .DIN4(n6154), 
        .Q(n6150) );
  nor2s1 U6149 ( .DIN1(n6155), .DIN2(n6156), .Q(n6154) );
  nor2s1 U6150 ( .DIN1(n6138), .DIN2(n6146), .Q(n6156) );
  nor2s1 U6151 ( .DIN1(n5485), .DIN2(n5123), .Q(n6155) );
  nnd2s1 U6152 ( .DIN1(n5250), .DIN2(n5128), .Q(n6152) );
  nnd2s1 U6153 ( .DIN1(n5441), .DIN2(n5108), .Q(n6151) );
  nnd3s1 U6154 ( .DIN1(n6157), .DIN2(n6158), .DIN3(n6159), .Q(n6149) );
  nnd2s1 U6155 ( .DIN1(n5451), .DIN2(n6160), .Q(n6159) );
  nnd2s1 U6156 ( .DIN1(n5775), .DIN2(n5464), .Q(n6160) );
  nnd2s1 U6157 ( .DIN1(n5249), .DIN2(n6161), .Q(n6158) );
  nnd2s1 U6158 ( .DIN1(n5797), .DIN2(n5740), .Q(n6161) );
  nnd2s1 U6159 ( .DIN1(n5110), .DIN2(n5483), .Q(n6157) );
  nnd2s1 U6160 ( .DIN1(n5466), .DIN2(n5741), .Q(n5483) );
  nor2s1 U6161 ( .DIN1(n6162), .DIN2(n5268), .Q(n6148) );
  nor2s1 U6162 ( .DIN1(n5138), .DIN2(n5120), .Q(n6162) );
  nor2s1 U6163 ( .DIN1(n6163), .DIN2(n5772), .Q(n6147) );
  and2s1 U6164 ( .DIN1(n5449), .DIN2(n6164), .Q(n6163) );
  nor4s1 U6165 ( .DIN1(n6165), .DIN2(n6166), .DIN3(n6167), .DIN4(n6168), 
        .Q(n5435) );
  nnd4s1 U6166 ( .DIN1(n6169), .DIN2(n6170), .DIN3(n6171), .DIN4(n6172), 
        .Q(n6168) );
  nnd2s1 U6167 ( .DIN1(n5754), .DIN2(n5452), .Q(n6172) );
  nor2s1 U6168 ( .DIN1(n6173), .DIN2(n6174), .Q(n6171) );
  nor2s1 U6169 ( .DIN1(n5268), .DIN2(n6175), .Q(n6173) );
  nnd2s1 U6170 ( .DIN1(n5440), .DIN2(n5459), .Q(n6170) );
  nnd2s1 U6171 ( .DIN1(n5442), .DIN2(n5116), .Q(n6169) );
  nnd3s1 U6172 ( .DIN1(n6176), .DIN2(n6177), .DIN3(n6178), .Q(n6167) );
  nnd2s1 U6173 ( .DIN1(n5108), .DIN2(n6179), .Q(n6178) );
  nnd2s1 U6174 ( .DIN1(n5124), .DIN2(n6180), .Q(n6177) );
  nnd2s1 U6175 ( .DIN1(n5772), .DIN2(n5740), .Q(n6180) );
  nnd2s1 U6176 ( .DIN1(n5755), .DIN2(n6181), .Q(n6176) );
  nnd3s1 U6177 ( .DIN1(n5744), .DIN2(n6146), .DIN3(n6182), .Q(n6181) );
  nor2s1 U6178 ( .DIN1(n5123), .DIN2(n5127), .Q(n6166) );
  nor2s1 U6179 ( .DIN1(n5270), .DIN2(n5119), .Q(n6165) );
  nor3s1 U6180 ( .DIN1(n6183), .DIN2(n6184), .DIN3(n6185), .Q(n5244) );
  nnd4s1 U6181 ( .DIN1(n5748), .DIN2(n5437), .DIN3(n5722), .DIN4(n6186), 
        .Q(n6185) );
  and3s1 U6182 ( .DIN1(n6187), .DIN2(n6188), .DIN3(n6189), .Q(n6186) );
  nnd2s1 U6183 ( .DIN1(n5442), .DIN2(n5107), .Q(n6189) );
  nnd2s1 U6184 ( .DIN1(n5137), .DIN2(n5265), .Q(n6187) );
  nor4s1 U6185 ( .DIN1(n6190), .DIN2(n6191), .DIN3(n6192), .DIN4(n6193), 
        .Q(n5722) );
  nnd4s1 U6186 ( .DIN1(n6194), .DIN2(n6195), .DIN3(n6196), .DIN4(n6197), 
        .Q(n6193) );
  nnd2s1 U6187 ( .DIN1(n5442), .DIN2(n6198), .Q(n6197) );
  nnd2s1 U6188 ( .DIN1(n6199), .DIN2(n5744), .Q(n6198) );
  nor2s1 U6189 ( .DIN1(n6200), .DIN2(n6201), .Q(n6196) );
  nor2s1 U6190 ( .DIN1(n6202), .DIN2(n5485), .Q(n6201) );
  nor2s1 U6191 ( .DIN1(n5137), .DIN2(n5272), .Q(n6202) );
  nor2s1 U6192 ( .DIN1(n6203), .DIN2(n5126), .Q(n6200) );
  nor2s1 U6193 ( .DIN1(n6204), .DIN2(n5441), .Q(n6203) );
  nnd2s1 U6194 ( .DIN1(n5116), .DIN2(n6205), .Q(n6195) );
  nnd3s1 U6195 ( .DIN1(n5127), .DIN2(n5771), .DIN3(n6175), .Q(n6205) );
  nnd2s1 U6196 ( .DIN1(n5755), .DIN2(n6204), .Q(n6194) );
  nnd3s1 U6197 ( .DIN1(n6206), .DIN2(n6207), .DIN3(n6208), .Q(n6192) );
  nnd2s1 U6198 ( .DIN1(n6209), .DIN2(n5482), .Q(n6208) );
  nnd2s1 U6199 ( .DIN1(n5106), .DIN2(n5109), .Q(n6207) );
  nnd2s1 U6200 ( .DIN1(n5110), .DIN2(n5249), .Q(n6206) );
  nor2s1 U6201 ( .DIN1(n6138), .DIN2(n5268), .Q(n6191) );
  nor2s1 U6202 ( .DIN1(n6146), .DIN2(n5797), .Q(n6190) );
  nor4s1 U6203 ( .DIN1(n6210), .DIN2(n6211), .DIN3(n6212), .DIN4(n6213), 
        .Q(n5437) );
  nnd4s1 U6204 ( .DIN1(n6214), .DIN2(n6215), .DIN3(n6216), .DIN4(n6217), 
        .Q(n6213) );
  nnd2s1 U6205 ( .DIN1(n5107), .DIN2(n5128), .Q(n6217) );
  nnd2s1 U6206 ( .DIN1(n5265), .DIN2(n5451), .Q(n6216) );
  nnd2s1 U6207 ( .DIN1(n5472), .DIN2(n5116), .Q(n6215) );
  nnd2s1 U6208 ( .DIN1(n5442), .DIN2(n5440), .Q(n6214) );
  nnd3s1 U6209 ( .DIN1(n6218), .DIN2(n6219), .DIN3(n6220), .Q(n6212) );
  nnd2s1 U6210 ( .DIN1(n5139), .DIN2(n6221), .Q(n6220) );
  nnd3s1 U6211 ( .DIN1(n5461), .DIN2(n5268), .DIN3(n5741), .Q(n6221) );
  nnd2s1 U6212 ( .DIN1(n5475), .DIN2(n6222), .Q(n6219) );
  nnd2s1 U6213 ( .DIN1(n6164), .DIN2(n5461), .Q(n6222) );
  nor2s1 U6214 ( .DIN1(n6209), .DIN2(n6204), .Q(n6164) );
  nnd2s1 U6215 ( .DIN1(n5754), .DIN2(n6223), .Q(n6218) );
  nnd2s1 U6216 ( .DIN1(n6139), .DIN2(n5797), .Q(n6223) );
  nor2s1 U6217 ( .DIN1(n5744), .DIN2(n5775), .Q(n6211) );
  nor2s1 U6218 ( .DIN1(n5467), .DIN2(n5772), .Q(n6210) );
  hi1s1 U6219 ( .DIN(n5129), .Q(n5467) );
  nor2s1 U6220 ( .DIN1(n6224), .DIN2(n6225), .Q(n5748) );
  nnd4s1 U6221 ( .DIN1(n6226), .DIN2(n6227), .DIN3(n6228), .DIN4(n6229), 
        .Q(n6225) );
  nnd2s1 U6222 ( .DIN1(n5107), .DIN2(n6230), .Q(n6229) );
  nnd3s1 U6223 ( .DIN1(n5772), .DIN2(n6138), .DIN3(n6175), .Q(n6230) );
  nnd2s1 U6224 ( .DIN1(n5106), .DIN2(n5441), .Q(n6227) );
  nnd4s1 U6225 ( .DIN1(n6231), .DIN2(n6232), .DIN3(n6233), .DIN4(n6234), 
        .Q(n6224) );
  nnd2s1 U6226 ( .DIN1(n5128), .DIN2(n6235), .Q(n6234) );
  nnd2s1 U6227 ( .DIN1(n6236), .DIN2(n5268), .Q(n6235) );
  nnd2s1 U6228 ( .DIN1(n5138), .DIN2(n6237), .Q(n6233) );
  nnd2s1 U6229 ( .DIN1(n5124), .DIN2(n6238), .Q(n6232) );
  nnd2s1 U6230 ( .DIN1(n5775), .DIN2(n6175), .Q(n6238) );
  nnd2s1 U6231 ( .DIN1(n5754), .DIN2(n6239), .Q(n6231) );
  nnd2s1 U6232 ( .DIN1(n5255), .DIN2(n5771), .Q(n6239) );
  nnd3s1 U6233 ( .DIN1(n6240), .DIN2(n6241), .DIN3(n6242), .Q(n6184) );
  nnd2s1 U6234 ( .DIN1(n5108), .DIN2(n5116), .Q(n6242) );
  nnd2s1 U6235 ( .DIN1(n6204), .DIN2(n6243), .Q(n6241) );
  nnd3s1 U6236 ( .DIN1(n6138), .DIN2(n5127), .DIN3(n6244), .Q(n6243) );
  or2s1 U6237 ( .DIN1(n5461), .DIN2(n6245), .Q(n6240) );
  nnd3s1 U6238 ( .DIN1(n6246), .DIN2(n6247), .DIN3(n6248), .Q(n6183) );
  nnd2s1 U6239 ( .DIN1(n5124), .DIN2(n6249), .Q(n6248) );
  nnd2s1 U6240 ( .DIN1(n5779), .DIN2(n5774), .Q(n6249) );
  nnd2s1 U6241 ( .DIN1(n5459), .DIN2(n6250), .Q(n6247) );
  or2s1 U6242 ( .DIN1(n5486), .DIN2(n5109), .Q(n6250) );
  nnd2s1 U6243 ( .DIN1(n5268), .DIN2(n5254), .Q(n5486) );
  nnd2s1 U6244 ( .DIN1(n5482), .DIN2(n6251), .Q(n6246) );
  nnd2s1 U6245 ( .DIN1(n5122), .DIN2(n5449), .Q(n6251) );
  nnd2s1 U6246 ( .DIN1(n5265), .DIN2(n5250), .Q(n6126) );
  nnd2s1 U6247 ( .DIN1(n5120), .DIN2(n5440), .Q(n6125) );
  nnd3s1 U6248 ( .DIN1(n6252), .DIN2(n6253), .DIN3(n6254), .Q(n6123) );
  nnd2s1 U6249 ( .DIN1(n6209), .DIN2(n5128), .Q(n6254) );
  nnd2s1 U6250 ( .DIN1(n5731), .DIN2(n6255), .Q(n6253) );
  nnd4s1 U6251 ( .DIN1(n6256), .DIN2(n6257), .DIN3(n6258), .DIN4(n6259), 
        .Q(n6122) );
  nnd2s1 U6252 ( .DIN1(n5475), .DIN2(n6260), .Q(n6259) );
  nnd2s1 U6253 ( .DIN1(n5270), .DIN2(n5481), .Q(n6260) );
  nor2s1 U6254 ( .DIN1(n5441), .DIN2(n5451), .Q(n5270) );
  nnd2s1 U6255 ( .DIN1(n5451), .DIN2(n6261), .Q(n6258) );
  nnd2s1 U6256 ( .DIN1(n5463), .DIN2(n5774), .Q(n6261) );
  nnd2s1 U6257 ( .DIN1(n5140), .DIN2(n6262), .Q(n6257) );
  nnd2s1 U6258 ( .DIN1(n5464), .DIN2(n5127), .Q(n6262) );
  nnd2s1 U6259 ( .DIN1(n5116), .DIN2(n5763), .Q(n6256) );
  or3s1 U6260 ( .DIN1(n6263), .DIN2(n6264), .DIN3(n6265), .Q(n4912) );
  nnd4s1 U6261 ( .DIN1(n6266), .DIN2(n6267), .DIN3(n5278), .DIN4(n6268), 
        .Q(n6265) );
  and3s1 U6262 ( .DIN1(n5491), .DIN2(n5835), .DIN3(n5801), .Q(n6268) );
  nor4s1 U6263 ( .DIN1(n6269), .DIN2(n6270), .DIN3(n6271), .DIN4(n6272), 
        .Q(n5801) );
  nnd4s1 U6264 ( .DIN1(n6273), .DIN2(n6274), .DIN3(n6275), .DIN4(n6276), 
        .Q(n6272) );
  nnd2s1 U6265 ( .DIN1(n5303), .DIN2(n5510), .Q(n6276) );
  nor2s1 U6266 ( .DIN1(n6277), .DIN2(n6278), .Q(n6275) );
  nor2s1 U6267 ( .DIN1(n6279), .DIN2(n5302), .Q(n6278) );
  nor2s1 U6268 ( .DIN1(n5544), .DIN2(n6280), .Q(n6277) );
  nnd2s1 U6269 ( .DIN1(n5498), .DIN2(n5511), .Q(n6274) );
  nnd2s1 U6270 ( .DIN1(n5294), .DIN2(n5519), .Q(n6273) );
  nnd3s1 U6271 ( .DIN1(n6281), .DIN2(n6282), .DIN3(n6283), .Q(n6271) );
  nnd2s1 U6272 ( .DIN1(n5545), .DIN2(n5550), .Q(n6283) );
  nnd2s1 U6273 ( .DIN1(n6284), .DIN2(n6285), .Q(n6282) );
  nnd3s1 U6274 ( .DIN1(n5861), .DIN2(n5826), .DIN3(n6279), .Q(n6285) );
  nnd2s1 U6275 ( .DIN1(n5841), .DIN2(n6286), .Q(n6281) );
  nnd3s1 U6276 ( .DIN1(n5506), .DIN2(n5292), .DIN3(n5301), .Q(n6286) );
  nor2s1 U6277 ( .DIN1(n5860), .DIN2(n5506), .Q(n6270) );
  nor2s1 U6278 ( .DIN1(n6287), .DIN2(n6288), .Q(n6269) );
  nor4s1 U6279 ( .DIN1(n6289), .DIN2(n6290), .DIN3(n6291), .DIN4(n6292), 
        .Q(n5835) );
  nnd4s1 U6280 ( .DIN1(n6293), .DIN2(n6294), .DIN3(n6295), .DIN4(n6296), 
        .Q(n6292) );
  nor2s1 U6281 ( .DIN1(n6297), .DIN2(n6298), .Q(n6296) );
  nor2s1 U6282 ( .DIN1(n6288), .DIN2(n6279), .Q(n6298) );
  nor2s1 U6283 ( .DIN1(n5548), .DIN2(n5292), .Q(n6297) );
  nnd2s1 U6284 ( .DIN1(n5285), .DIN2(n5542), .Q(n6294) );
  nnd2s1 U6285 ( .DIN1(n5283), .DIN2(n5497), .Q(n6293) );
  nnd3s1 U6286 ( .DIN1(n6299), .DIN2(n6300), .DIN3(n6301), .Q(n6291) );
  nnd2s1 U6287 ( .DIN1(n5508), .DIN2(n6302), .Q(n6301) );
  nnd2s1 U6288 ( .DIN1(n5862), .DIN2(n5524), .Q(n6302) );
  nnd2s1 U6289 ( .DIN1(n5284), .DIN2(n6303), .Q(n6300) );
  nnd2s1 U6290 ( .DIN1(n5886), .DIN2(n5826), .Q(n6303) );
  nnd2s1 U6291 ( .DIN1(n5516), .DIN2(n5546), .Q(n6299) );
  nnd2s1 U6292 ( .DIN1(n5527), .DIN2(n5827), .Q(n5546) );
  nor2s1 U6293 ( .DIN1(n6304), .DIN2(n5306), .Q(n6290) );
  nor2s1 U6294 ( .DIN1(n5286), .DIN2(n5525), .Q(n6304) );
  nor2s1 U6295 ( .DIN1(n6305), .DIN2(n5858), .Q(n6289) );
  and2s1 U6296 ( .DIN1(n5506), .DIN2(n6306), .Q(n6305) );
  nor4s1 U6297 ( .DIN1(n6307), .DIN2(n6308), .DIN3(n6309), .DIN4(n6310), 
        .Q(n5491) );
  nnd4s1 U6298 ( .DIN1(n6311), .DIN2(n6312), .DIN3(n6313), .DIN4(n6314), 
        .Q(n6310) );
  nnd2s1 U6299 ( .DIN1(n5511), .DIN2(n5840), .Q(n6314) );
  nor2s1 U6300 ( .DIN1(n6315), .DIN2(n6316), .Q(n6313) );
  nor2s1 U6301 ( .DIN1(n5306), .DIN2(n6317), .Q(n6315) );
  nnd2s1 U6302 ( .DIN1(n5519), .DIN2(n5509), .Q(n6312) );
  nnd2s1 U6303 ( .DIN1(n5884), .DIN2(n5499), .Q(n6311) );
  nnd3s1 U6304 ( .DIN1(n6318), .DIN2(n6319), .DIN3(n6320), .Q(n6309) );
  nnd2s1 U6305 ( .DIN1(n5283), .DIN2(n6321), .Q(n6320) );
  nnd2s1 U6306 ( .DIN1(n5294), .DIN2(n6322), .Q(n6319) );
  nnd2s1 U6307 ( .DIN1(n5858), .DIN2(n5826), .Q(n6322) );
  nnd2s1 U6308 ( .DIN1(n5841), .DIN2(n6323), .Q(n6318) );
  nnd3s1 U6309 ( .DIN1(n5830), .DIN2(n6288), .DIN3(n6324), .Q(n6323) );
  nor2s1 U6310 ( .DIN1(n5860), .DIN2(n5292), .Q(n6308) );
  nor2s1 U6311 ( .DIN1(n5309), .DIN2(n5549), .Q(n6307) );
  nor3s1 U6312 ( .DIN1(n6325), .DIN2(n6326), .DIN3(n6327), .Q(n5278) );
  nnd4s1 U6313 ( .DIN1(n5834), .DIN2(n5493), .DIN3(n5805), .DIN4(n6328), 
        .Q(n6327) );
  and3s1 U6314 ( .DIN1(n6329), .DIN2(n6330), .DIN3(n6331), .Q(n6328) );
  nnd2s1 U6315 ( .DIN1(n5816), .DIN2(n5499), .Q(n6331) );
  nnd2s1 U6316 ( .DIN1(n5303), .DIN2(n5537), .Q(n6329) );
  nor4s1 U6317 ( .DIN1(n6332), .DIN2(n6333), .DIN3(n6334), .DIN4(n6335), 
        .Q(n5805) );
  nnd4s1 U6318 ( .DIN1(n6336), .DIN2(n6337), .DIN3(n6338), .DIN4(n6339), 
        .Q(n6335) );
  nnd2s1 U6319 ( .DIN1(n5499), .DIN2(n6340), .Q(n6339) );
  nnd2s1 U6320 ( .DIN1(n6341), .DIN2(n5830), .Q(n6340) );
  nor2s1 U6321 ( .DIN1(n6342), .DIN2(n6343), .Q(n6338) );
  nor2s1 U6322 ( .DIN1(n6344), .DIN2(n5548), .Q(n6343) );
  nor2s1 U6323 ( .DIN1(n5537), .DIN2(n5311), .Q(n6344) );
  nor2s1 U6324 ( .DIN1(n6345), .DIN2(n6346), .Q(n6342) );
  nor2s1 U6325 ( .DIN1(n6347), .DIN2(n5497), .Q(n6345) );
  nnd2s1 U6326 ( .DIN1(n5884), .DIN2(n6348), .Q(n6337) );
  nnd3s1 U6327 ( .DIN1(n5860), .DIN2(n5857), .DIN3(n6317), .Q(n6348) );
  nnd2s1 U6328 ( .DIN1(n5841), .DIN2(n6347), .Q(n6336) );
  nnd3s1 U6329 ( .DIN1(n6349), .DIN2(n6350), .DIN3(n6351), .Q(n6334) );
  nnd2s1 U6330 ( .DIN1(n6352), .DIN2(n5545), .Q(n6351) );
  nnd2s1 U6331 ( .DIN1(n6284), .DIN2(n5814), .Q(n6350) );
  nnd2s1 U6332 ( .DIN1(n5516), .DIN2(n5284), .Q(n6349) );
  nor2s1 U6333 ( .DIN1(n6279), .DIN2(n5306), .Q(n6333) );
  nor2s1 U6334 ( .DIN1(n6288), .DIN2(n5886), .Q(n6332) );
  nor4s1 U6335 ( .DIN1(n6353), .DIN2(n6354), .DIN3(n6355), .DIN4(n6356), 
        .Q(n5493) );
  nnd4s1 U6336 ( .DIN1(n6357), .DIN2(n6358), .DIN3(n6359), .DIN4(n6360), 
        .Q(n6356) );
  nnd2s1 U6337 ( .DIN1(n5816), .DIN2(n5542), .Q(n6360) );
  nnd2s1 U6338 ( .DIN1(n5303), .DIN2(n5508), .Q(n6359) );
  nnd2s1 U6339 ( .DIN1(n5884), .DIN2(n5533), .Q(n6358) );
  nnd2s1 U6340 ( .DIN1(n5499), .DIN2(n5509), .Q(n6357) );
  nnd3s1 U6341 ( .DIN1(n6361), .DIN2(n6362), .DIN3(n6363), .Q(n6355) );
  nnd2s1 U6342 ( .DIN1(n5307), .DIN2(n6364), .Q(n6363) );
  nnd3s1 U6343 ( .DIN1(n5827), .DIN2(n5521), .DIN3(n5306), .Q(n6364) );
  nnd2s1 U6344 ( .DIN1(n5536), .DIN2(n6365), .Q(n6362) );
  nnd2s1 U6345 ( .DIN1(n6306), .DIN2(n5521), .Q(n6365) );
  nor2s1 U6346 ( .DIN1(n6352), .DIN2(n6347), .Q(n6306) );
  nnd2s1 U6347 ( .DIN1(n5840), .DIN2(n6366), .Q(n6361) );
  nnd2s1 U6348 ( .DIN1(n6280), .DIN2(n5886), .Q(n6366) );
  nor2s1 U6349 ( .DIN1(n5830), .DIN2(n5862), .Q(n6354) );
  nor2s1 U6350 ( .DIN1(n5528), .DIN2(n5858), .Q(n6353) );
  hi1s1 U6351 ( .DIN(n6367), .Q(n5528) );
  nor2s1 U6352 ( .DIN1(n6368), .DIN2(n6369), .Q(n5834) );
  nnd4s1 U6353 ( .DIN1(n6370), .DIN2(n6371), .DIN3(n6372), .DIN4(n6373), 
        .Q(n6369) );
  nnd2s1 U6354 ( .DIN1(n5816), .DIN2(n6374), .Q(n6373) );
  nnd3s1 U6355 ( .DIN1(n5858), .DIN2(n6279), .DIN3(n6317), .Q(n6374) );
  nnd2s1 U6356 ( .DIN1(n5497), .DIN2(n5814), .Q(n6371) );
  nnd4s1 U6357 ( .DIN1(n6375), .DIN2(n6376), .DIN3(n6377), .DIN4(n6378), 
        .Q(n6368) );
  nnd2s1 U6358 ( .DIN1(n5542), .DIN2(n6379), .Q(n6378) );
  nnd2s1 U6359 ( .DIN1(n6380), .DIN2(n5306), .Q(n6379) );
  nnd2s1 U6360 ( .DIN1(n5286), .DIN2(n6381), .Q(n6377) );
  nnd2s1 U6361 ( .DIN1(n5294), .DIN2(n6382), .Q(n6376) );
  nnd2s1 U6362 ( .DIN1(n5862), .DIN2(n6317), .Q(n6382) );
  nnd2s1 U6363 ( .DIN1(n5840), .DIN2(n6383), .Q(n6375) );
  nnd2s1 U6364 ( .DIN1(n5291), .DIN2(n5857), .Q(n6383) );
  nnd3s1 U6365 ( .DIN1(n6384), .DIN2(n6385), .DIN3(n6386), .Q(n6326) );
  nnd2s1 U6366 ( .DIN1(n5283), .DIN2(n5884), .Q(n6386) );
  nnd2s1 U6367 ( .DIN1(n6347), .DIN2(n6387), .Q(n6385) );
  nnd3s1 U6368 ( .DIN1(n5860), .DIN2(n6279), .DIN3(n6388), .Q(n6387) );
  or2s1 U6369 ( .DIN1(n5521), .DIN2(n6389), .Q(n6384) );
  nnd3s1 U6370 ( .DIN1(n6390), .DIN2(n6391), .DIN3(n6392), .Q(n6325) );
  nnd2s1 U6371 ( .DIN1(n5294), .DIN2(n6393), .Q(n6392) );
  nnd2s1 U6372 ( .DIN1(n5867), .DIN2(n5861), .Q(n6393) );
  nnd2s1 U6373 ( .DIN1(n5519), .DIN2(n6394), .Q(n6391) );
  or2s1 U6374 ( .DIN1(n5550), .DIN2(n6284), .Q(n6394) );
  nnd2s1 U6375 ( .DIN1(n5306), .DIN2(n5290), .Q(n5550) );
  nnd2s1 U6376 ( .DIN1(n5545), .DIN2(n6395), .Q(n6390) );
  nnd2s1 U6377 ( .DIN1(n5822), .DIN2(n5506), .Q(n6395) );
  nnd2s1 U6378 ( .DIN1(n5303), .DIN2(n5285), .Q(n6267) );
  nnd2s1 U6379 ( .DIN1(n5509), .DIN2(n5525), .Q(n6266) );
  nnd3s1 U6380 ( .DIN1(n6396), .DIN2(n6397), .DIN3(n6398), .Q(n6264) );
  nnd2s1 U6381 ( .DIN1(n6352), .DIN2(n5542), .Q(n6398) );
  nnd2s1 U6382 ( .DIN1(n5815), .DIN2(n6399), .Q(n6397) );
  nnd4s1 U6383 ( .DIN1(n6400), .DIN2(n6401), .DIN3(n6402), .DIN4(n6403), 
        .Q(n6263) );
  nnd2s1 U6384 ( .DIN1(n5536), .DIN2(n6404), .Q(n6403) );
  nnd2s1 U6385 ( .DIN1(n5309), .DIN2(n5544), .Q(n6404) );
  nor2s1 U6386 ( .DIN1(n5497), .DIN2(n5508), .Q(n5309) );
  nnd2s1 U6387 ( .DIN1(n5508), .DIN2(n6405), .Q(n6402) );
  nnd2s1 U6388 ( .DIN1(n5523), .DIN2(n5861), .Q(n6405) );
  nnd2s1 U6389 ( .DIN1(n5498), .DIN2(n6406), .Q(n6401) );
  nnd2s1 U6390 ( .DIN1(n5524), .DIN2(n5860), .Q(n6406) );
  nnd2s1 U6391 ( .DIN1(n5884), .DIN2(n5849), .Q(n6400) );
  or3s1 U6392 ( .DIN1(n6407), .DIN2(n6408), .DIN3(n6409), .Q(n4989) );
  nnd4s1 U6393 ( .DIN1(n6410), .DIN2(n6411), .DIN3(n6412), .DIN4(n6413), 
        .Q(n6409) );
  and3s1 U6394 ( .DIN1(n6414), .DIN2(n6415), .DIN3(n6416), .Q(n6413) );
  nnd2s1 U6395 ( .DIN1(n5366), .DIN2(n5373), .Q(n6411) );
  nnd2s1 U6396 ( .DIN1(n5359), .DIN2(n5197), .Q(n6410) );
  nnd3s1 U6397 ( .DIN1(n6417), .DIN2(n6418), .DIN3(n6419), .Q(n6408) );
  nnd2s1 U6398 ( .DIN1(n5568), .DIN2(n5357), .Q(n6419) );
  or2s1 U6399 ( .DIN1(n5592), .DIN2(n6420), .Q(n6418) );
  nnd2s1 U6400 ( .DIN1(n5621), .DIN2(n5408), .Q(n6417) );
  nnd4s1 U6401 ( .DIN1(n6421), .DIN2(n6422), .DIN3(n6423), .DIN4(n6424), 
        .Q(n6407) );
  nnd2s1 U6402 ( .DIN1(n5970), .DIN2(n6425), .Q(n6424) );
  nnd2s1 U6403 ( .DIN1(n6010), .DIN2(n5563), .Q(n6425) );
  nnd2s1 U6404 ( .DIN1(n5372), .DIN2(n6426), .Q(n6423) );
  nnd2s1 U6405 ( .DIN1(n5594), .DIN2(n5212), .Q(n6426) );
  nor2s1 U6406 ( .DIN1(n5583), .DIN2(n5582), .Q(n5594) );
  nnd2s1 U6407 ( .DIN1(n5400), .DIN2(n6427), .Q(n6422) );
  nnd2s1 U6408 ( .DIN1(n5412), .DIN2(n5564), .Q(n6427) );
  nnd2s1 U6409 ( .DIN1(n5214), .DIN2(n6428), .Q(n6421) );
  xor2s1 U6410 ( .DIN1(n4923), .DIN2(n6429), .Q(n6119) );
  xor2s1 U6411 ( .DIN1(n1440), .DIN2(n4899), .Q(n6429) );
  or3s1 U6412 ( .DIN1(n6430), .DIN2(n6431), .DIN3(n6432), .Q(n4899) );
  nnd4s1 U6413 ( .DIN1(n6433), .DIN2(n6434), .DIN3(n5318), .DIN4(n6435), 
        .Q(n6432) );
  and3s1 U6414 ( .DIN1(n5645), .DIN2(n6064), .DIN3(n6033), .Q(n6435) );
  nor4s1 U6415 ( .DIN1(n6436), .DIN2(n6437), .DIN3(n6438), .DIN4(n6439), 
        .Q(n6033) );
  nnd4s1 U6416 ( .DIN1(n6440), .DIN2(n6441), .DIN3(n6442), .DIN4(n6443), 
        .Q(n6439) );
  nnd2s1 U6417 ( .DIN1(n5156), .DIN2(n5339), .Q(n6443) );
  nor2s1 U6418 ( .DIN1(n6444), .DIN2(n6445), .Q(n6442) );
  nor2s1 U6419 ( .DIN1(n5338), .DIN2(n6446), .Q(n6445) );
  nor2s1 U6420 ( .DIN1(n5691), .DIN2(n6447), .Q(n6444) );
  nnd2s1 U6421 ( .DIN1(n5185), .DIN2(n5662), .Q(n6441) );
  nnd2s1 U6422 ( .DIN1(n5669), .DIN2(n5169), .Q(n6440) );
  nnd3s1 U6423 ( .DIN1(n6448), .DIN2(n6449), .DIN3(n6450), .Q(n6438) );
  nnd2s1 U6424 ( .DIN1(n5692), .DIN2(n5696), .Q(n6450) );
  nnd2s1 U6425 ( .DIN1(n5154), .DIN2(n6451), .Q(n6449) );
  nnd3s1 U6426 ( .DIN1(n6089), .DIN2(n6055), .DIN3(n6446), .Q(n6451) );
  nnd2s1 U6427 ( .DIN1(n6070), .DIN2(n6452), .Q(n6448) );
  nnd3s1 U6428 ( .DIN1(n5659), .DIN2(n5168), .DIN3(n5337), .Q(n6452) );
  nor2s1 U6429 ( .DIN1(n5659), .DIN2(n5172), .Q(n6437) );
  nor2s1 U6430 ( .DIN1(n6453), .DIN2(n6454), .Q(n6436) );
  nor4s1 U6431 ( .DIN1(n6455), .DIN2(n6456), .DIN3(n6457), .DIN4(n6458), 
        .Q(n6064) );
  nnd4s1 U6432 ( .DIN1(n6459), .DIN2(n6460), .DIN3(n6461), .DIN4(n6462), 
        .Q(n6458) );
  nor2s1 U6433 ( .DIN1(n6463), .DIN2(n6464), .Q(n6462) );
  nor2s1 U6434 ( .DIN1(n6446), .DIN2(n6454), .Q(n6464) );
  nor2s1 U6435 ( .DIN1(n5695), .DIN2(n5168), .Q(n6463) );
  nnd2s1 U6436 ( .DIN1(n5324), .DIN2(n5173), .Q(n6460) );
  nnd2s1 U6437 ( .DIN1(n5651), .DIN2(n5153), .Q(n6459) );
  nnd3s1 U6438 ( .DIN1(n6465), .DIN2(n6466), .DIN3(n6467), .Q(n6457) );
  nnd2s1 U6439 ( .DIN1(n5661), .DIN2(n6468), .Q(n6467) );
  nnd2s1 U6440 ( .DIN1(n6090), .DIN2(n5674), .Q(n6468) );
  nnd2s1 U6441 ( .DIN1(n5323), .DIN2(n6469), .Q(n6466) );
  nnd2s1 U6442 ( .DIN1(n6112), .DIN2(n6055), .Q(n6469) );
  nnd2s1 U6443 ( .DIN1(n5155), .DIN2(n5693), .Q(n6465) );
  nnd2s1 U6444 ( .DIN1(n5676), .DIN2(n6056), .Q(n5693) );
  nor2s1 U6445 ( .DIN1(n6470), .DIN2(n5342), .Q(n6456) );
  nor2s1 U6446 ( .DIN1(n5183), .DIN2(n5165), .Q(n6470) );
  nor2s1 U6447 ( .DIN1(n6471), .DIN2(n6087), .Q(n6455) );
  and2s1 U6448 ( .DIN1(n5659), .DIN2(n6472), .Q(n6471) );
  nor4s1 U6449 ( .DIN1(n6473), .DIN2(n6474), .DIN3(n6475), .DIN4(n6476), 
        .Q(n5645) );
  nnd4s1 U6450 ( .DIN1(n6477), .DIN2(n6478), .DIN3(n6479), .DIN4(n6480), 
        .Q(n6476) );
  nnd2s1 U6451 ( .DIN1(n6069), .DIN2(n5662), .Q(n6480) );
  nor2s1 U6452 ( .DIN1(n6481), .DIN2(n6482), .Q(n6479) );
  nor2s1 U6453 ( .DIN1(n5342), .DIN2(n6483), .Q(n6481) );
  nnd2s1 U6454 ( .DIN1(n5650), .DIN2(n5669), .Q(n6478) );
  nnd2s1 U6455 ( .DIN1(n5652), .DIN2(n5161), .Q(n6477) );
  nnd3s1 U6456 ( .DIN1(n6484), .DIN2(n6485), .DIN3(n6486), .Q(n6475) );
  nnd2s1 U6457 ( .DIN1(n5153), .DIN2(n6487), .Q(n6486) );
  nnd2s1 U6458 ( .DIN1(n5169), .DIN2(n6488), .Q(n6485) );
  nnd2s1 U6459 ( .DIN1(n6087), .DIN2(n6055), .Q(n6488) );
  nnd2s1 U6460 ( .DIN1(n6070), .DIN2(n6489), .Q(n6484) );
  nnd3s1 U6461 ( .DIN1(n6059), .DIN2(n6454), .DIN3(n6490), .Q(n6489) );
  nor2s1 U6462 ( .DIN1(n5168), .DIN2(n5172), .Q(n6474) );
  nor2s1 U6463 ( .DIN1(n5344), .DIN2(n5164), .Q(n6473) );
  nor3s1 U6464 ( .DIN1(n6491), .DIN2(n6492), .DIN3(n6493), .Q(n5318) );
  nnd4s1 U6465 ( .DIN1(n6063), .DIN2(n5647), .DIN3(n6037), .DIN4(n6494), 
        .Q(n6493) );
  and3s1 U6466 ( .DIN1(n6495), .DIN2(n6496), .DIN3(n6497), .Q(n6494) );
  nnd2s1 U6467 ( .DIN1(n5652), .DIN2(n5152), .Q(n6497) );
  nnd2s1 U6468 ( .DIN1(n5182), .DIN2(n5339), .Q(n6495) );
  nor4s1 U6469 ( .DIN1(n6498), .DIN2(n6499), .DIN3(n6500), .DIN4(n6501), 
        .Q(n6037) );
  nnd4s1 U6470 ( .DIN1(n6502), .DIN2(n6503), .DIN3(n6504), .DIN4(n6505), 
        .Q(n6501) );
  nnd2s1 U6471 ( .DIN1(n5652), .DIN2(n6506), .Q(n6505) );
  nnd2s1 U6472 ( .DIN1(n6507), .DIN2(n6059), .Q(n6506) );
  nor2s1 U6473 ( .DIN1(n6508), .DIN2(n6509), .Q(n6504) );
  nor2s1 U6474 ( .DIN1(n6510), .DIN2(n5695), .Q(n6509) );
  nor2s1 U6475 ( .DIN1(n5182), .DIN2(n5346), .Q(n6510) );
  nor2s1 U6476 ( .DIN1(n6511), .DIN2(n5171), .Q(n6508) );
  nor2s1 U6477 ( .DIN1(n6512), .DIN2(n5651), .Q(n6511) );
  nnd2s1 U6478 ( .DIN1(n5161), .DIN2(n6513), .Q(n6503) );
  nnd3s1 U6479 ( .DIN1(n5172), .DIN2(n6086), .DIN3(n6483), .Q(n6513) );
  nnd2s1 U6480 ( .DIN1(n6070), .DIN2(n6512), .Q(n6502) );
  nnd3s1 U6481 ( .DIN1(n6514), .DIN2(n6515), .DIN3(n6516), .Q(n6500) );
  nnd2s1 U6482 ( .DIN1(n6517), .DIN2(n5692), .Q(n6516) );
  nnd2s1 U6483 ( .DIN1(n5151), .DIN2(n5154), .Q(n6515) );
  nnd2s1 U6484 ( .DIN1(n5155), .DIN2(n5323), .Q(n6514) );
  nor2s1 U6485 ( .DIN1(n6446), .DIN2(n5342), .Q(n6499) );
  nor2s1 U6486 ( .DIN1(n6454), .DIN2(n6112), .Q(n6498) );
  nor4s1 U6487 ( .DIN1(n6518), .DIN2(n6519), .DIN3(n6520), .DIN4(n6521), 
        .Q(n5647) );
  nnd4s1 U6488 ( .DIN1(n6522), .DIN2(n6523), .DIN3(n6524), .DIN4(n6525), 
        .Q(n6521) );
  nnd2s1 U6489 ( .DIN1(n5152), .DIN2(n5173), .Q(n6525) );
  nnd2s1 U6490 ( .DIN1(n5339), .DIN2(n5661), .Q(n6524) );
  nnd2s1 U6491 ( .DIN1(n5682), .DIN2(n5161), .Q(n6523) );
  nnd2s1 U6492 ( .DIN1(n5652), .DIN2(n5650), .Q(n6522) );
  nnd3s1 U6493 ( .DIN1(n6526), .DIN2(n6527), .DIN3(n6528), .Q(n6520) );
  nnd2s1 U6494 ( .DIN1(n5184), .DIN2(n6529), .Q(n6528) );
  nnd3s1 U6495 ( .DIN1(n5671), .DIN2(n5342), .DIN3(n6056), .Q(n6529) );
  nnd2s1 U6496 ( .DIN1(n5685), .DIN2(n6530), .Q(n6527) );
  nnd2s1 U6497 ( .DIN1(n6472), .DIN2(n5671), .Q(n6530) );
  nor2s1 U6498 ( .DIN1(n6517), .DIN2(n6512), .Q(n6472) );
  nnd2s1 U6499 ( .DIN1(n6069), .DIN2(n6531), .Q(n6526) );
  nnd2s1 U6500 ( .DIN1(n6447), .DIN2(n6112), .Q(n6531) );
  nor2s1 U6501 ( .DIN1(n6059), .DIN2(n6090), .Q(n6519) );
  nor2s1 U6502 ( .DIN1(n5677), .DIN2(n6087), .Q(n6518) );
  hi1s1 U6503 ( .DIN(n5174), .Q(n5677) );
  nor2s1 U6504 ( .DIN1(n6532), .DIN2(n6533), .Q(n6063) );
  nnd4s1 U6505 ( .DIN1(n6534), .DIN2(n6535), .DIN3(n6536), .DIN4(n6537), 
        .Q(n6533) );
  nnd2s1 U6506 ( .DIN1(n5152), .DIN2(n6538), .Q(n6537) );
  nnd3s1 U6507 ( .DIN1(n6087), .DIN2(n6446), .DIN3(n6483), .Q(n6538) );
  nnd2s1 U6508 ( .DIN1(n5151), .DIN2(n5651), .Q(n6535) );
  nnd4s1 U6509 ( .DIN1(n6539), .DIN2(n6540), .DIN3(n6541), .DIN4(n6542), 
        .Q(n6532) );
  nnd2s1 U6510 ( .DIN1(n5173), .DIN2(n6543), .Q(n6542) );
  nnd2s1 U6511 ( .DIN1(n6544), .DIN2(n5342), .Q(n6543) );
  nnd2s1 U6512 ( .DIN1(n5183), .DIN2(n6545), .Q(n6541) );
  nnd2s1 U6513 ( .DIN1(n5169), .DIN2(n6546), .Q(n6540) );
  nnd2s1 U6514 ( .DIN1(n6090), .DIN2(n6483), .Q(n6546) );
  nnd2s1 U6515 ( .DIN1(n6069), .DIN2(n6547), .Q(n6539) );
  nnd2s1 U6516 ( .DIN1(n5329), .DIN2(n6086), .Q(n6547) );
  nnd3s1 U6517 ( .DIN1(n6548), .DIN2(n6549), .DIN3(n6550), .Q(n6492) );
  nnd2s1 U6518 ( .DIN1(n5153), .DIN2(n5161), .Q(n6550) );
  nnd2s1 U6519 ( .DIN1(n6512), .DIN2(n6551), .Q(n6549) );
  nnd3s1 U6520 ( .DIN1(n6446), .DIN2(n5172), .DIN3(n6552), .Q(n6551) );
  or2s1 U6521 ( .DIN1(n5671), .DIN2(n6553), .Q(n6548) );
  nnd3s1 U6522 ( .DIN1(n6554), .DIN2(n6555), .DIN3(n6556), .Q(n6491) );
  nnd2s1 U6523 ( .DIN1(n5169), .DIN2(n6557), .Q(n6556) );
  nnd2s1 U6524 ( .DIN1(n6094), .DIN2(n6089), .Q(n6557) );
  nnd2s1 U6525 ( .DIN1(n5669), .DIN2(n6558), .Q(n6555) );
  or2s1 U6526 ( .DIN1(n5696), .DIN2(n5154), .Q(n6558) );
  nnd2s1 U6527 ( .DIN1(n5342), .DIN2(n5328), .Q(n5696) );
  nnd2s1 U6528 ( .DIN1(n5692), .DIN2(n6559), .Q(n6554) );
  nnd2s1 U6529 ( .DIN1(n5167), .DIN2(n5659), .Q(n6559) );
  nnd2s1 U6530 ( .DIN1(n5339), .DIN2(n5324), .Q(n6434) );
  nnd2s1 U6531 ( .DIN1(n5165), .DIN2(n5650), .Q(n6433) );
  nnd3s1 U6532 ( .DIN1(n6560), .DIN2(n6561), .DIN3(n6562), .Q(n6431) );
  nnd2s1 U6533 ( .DIN1(n6517), .DIN2(n5173), .Q(n6562) );
  nnd2s1 U6534 ( .DIN1(n6046), .DIN2(n6563), .Q(n6561) );
  nnd4s1 U6535 ( .DIN1(n6564), .DIN2(n6565), .DIN3(n6566), .DIN4(n6567), 
        .Q(n6430) );
  nnd2s1 U6536 ( .DIN1(n5685), .DIN2(n6568), .Q(n6567) );
  nnd2s1 U6537 ( .DIN1(n5344), .DIN2(n5691), .Q(n6568) );
  nor2s1 U6538 ( .DIN1(n5651), .DIN2(n5661), .Q(n5344) );
  nnd2s1 U6539 ( .DIN1(n5661), .DIN2(n6569), .Q(n6566) );
  nnd2s1 U6540 ( .DIN1(n5673), .DIN2(n6089), .Q(n6569) );
  nnd2s1 U6541 ( .DIN1(n5185), .DIN2(n6570), .Q(n6565) );
  nnd2s1 U6542 ( .DIN1(n5674), .DIN2(n5172), .Q(n6570) );
  nnd2s1 U6543 ( .DIN1(n5161), .DIN2(n6078), .Q(n6564) );
  nnd2s1 U6544 ( .DIN1(n6571), .DIN2(n1605), .Q(n6116) );
  xor2s1 U6545 ( .DIN1(w3[3]), .DIN2(text_in_r[3]), .Q(n6571) );
  nnd3s1 U6546 ( .DIN1(n6572), .DIN2(n6573), .DIN3(n6574), .Q(N36) );
  nnd2s1 U6547 ( .DIN1(n1597), .DIN2(n6575), .Q(n6574) );
  xor2s1 U6548 ( .DIN1(w3[2]), .DIN2(text_in_r[2]), .Q(n6575) );
  nnd2s1 U6549 ( .DIN1(n6576), .DIN2(n4933), .Q(n6573) );
  nnd2s1 U6550 ( .DIN1(n6577), .DIN2(n6578), .Q(n6576) );
  nnd2s1 U6551 ( .DIN1(n4810), .DIN2(n6579), .Q(n6578) );
  nnd2s1 U6552 ( .DIN1(n6580), .DIN2(n4812), .Q(n6577) );
  nnd2s1 U6553 ( .DIN1(n5223), .DIN2(n6581), .Q(n6572) );
  nnd2s1 U6554 ( .DIN1(n6582), .DIN2(n6583), .Q(n6581) );
  nnd2s1 U6555 ( .DIN1(n4812), .DIN2(n6579), .Q(n6583) );
  and2s1 U6556 ( .DIN1(n4996), .DIN2(n1643), .Q(n4812) );
  nnd2s1 U6557 ( .DIN1(n6580), .DIN2(n4810), .Q(n6582) );
  nor2s1 U6558 ( .DIN1(n4996), .DIN2(n1594), .Q(n4810) );
  xor2s1 U6559 ( .DIN1(n4827), .DIN2(n4923), .Q(n4996) );
  or3s1 U6560 ( .DIN1(n6584), .DIN2(n6585), .DIN3(n6586), .Q(n4923) );
  nnd4s1 U6561 ( .DIN1(n6587), .DIN2(n6588), .DIN3(n6589), .DIN4(n6590), 
        .Q(n6586) );
  and3s1 U6562 ( .DIN1(n6591), .DIN2(n6592), .DIN3(n6593), .Q(n6590) );
  nnd2s1 U6563 ( .DIN1(n5510), .DIN2(n5525), .Q(n6588) );
  nnd2s1 U6564 ( .DIN1(n5884), .DIN2(n5511), .Q(n6587) );
  nnd3s1 U6565 ( .DIN1(n6594), .DIN2(n6595), .DIN3(n6596), .Q(n6585) );
  nnd2s1 U6566 ( .DIN1(n5283), .DIN2(n5509), .Q(n6596) );
  or2s1 U6567 ( .DIN1(n5822), .DIN2(n6597), .Q(n6595) );
  nnd2s1 U6568 ( .DIN1(n5840), .DIN2(n5542), .Q(n6594) );
  nnd4s1 U6569 ( .DIN1(n6598), .DIN2(n6599), .DIN3(n6600), .DIN4(n6601), 
        .Q(n6584) );
  nnd2s1 U6570 ( .DIN1(n6352), .DIN2(n6602), .Q(n6601) );
  nnd2s1 U6571 ( .DIN1(n6389), .DIN2(n5857), .Q(n6602) );
  nnd2s1 U6572 ( .DIN1(n5286), .DIN2(n6603), .Q(n6600) );
  nnd2s1 U6573 ( .DIN1(n5824), .DIN2(n5302), .Q(n6603) );
  nor2s1 U6574 ( .DIN1(n5816), .DIN2(n6347), .Q(n5824) );
  nnd2s1 U6575 ( .DIN1(n5307), .DIN2(n6604), .Q(n6599) );
  nnd2s1 U6576 ( .DIN1(n5498), .DIN2(n6605), .Q(n6598) );
  or3s1 U6577 ( .DIN1(n6606), .DIN2(n6607), .DIN3(n6608), .Q(n4827) );
  nnd4s1 U6578 ( .DIN1(n6609), .DIN2(n6610), .DIN3(n5133), .DIN4(n6611), 
        .Q(n6608) );
  and3s1 U6579 ( .DIN1(n6612), .DIN2(n6613), .DIN3(n6614), .Q(n6611) );
  nor3s1 U6580 ( .DIN1(n6615), .DIN2(n6616), .DIN3(n6617), .Q(n5133) );
  nnd4s1 U6581 ( .DIN1(n6618), .DIN2(n6619), .DIN3(n6620), .DIN4(n6621), 
        .Q(n6617) );
  and3s1 U6582 ( .DIN1(n6622), .DIN2(n6623), .DIN3(n6624), .Q(n6621) );
  nnd2s1 U6583 ( .DIN1(n5261), .DIN2(n5140), .Q(n6624) );
  nnd2s1 U6584 ( .DIN1(n5106), .DIN2(n5440), .Q(n6623) );
  nnd2s1 U6585 ( .DIN1(n5120), .DIN2(n5451), .Q(n6622) );
  nnd3s1 U6586 ( .DIN1(n6625), .DIN2(n6626), .DIN3(n6228), .Q(n6616) );
  nnd2s1 U6587 ( .DIN1(n5442), .DIN2(n6204), .Q(n6228) );
  or2s1 U6588 ( .DIN1(n5126), .DIN2(n6236), .Q(n6626) );
  nor2s1 U6589 ( .DIN1(n5137), .DIN2(n5109), .Q(n6236) );
  nnd2s1 U6590 ( .DIN1(n5475), .DIN2(n5272), .Q(n6625) );
  nnd2s1 U6591 ( .DIN1(n5466), .DIN2(n5263), .Q(n5272) );
  nnd4s1 U6592 ( .DIN1(n6627), .DIN2(n6628), .DIN3(n6629), .DIN4(n6630), 
        .Q(n6615) );
  nnd2s1 U6593 ( .DIN1(n5731), .DIN2(n6631), .Q(n6630) );
  nnd2s1 U6594 ( .DIN1(n5139), .DIN2(n6632), .Q(n6629) );
  nnd2s1 U6595 ( .DIN1(n5263), .DIN2(n5481), .Q(n6632) );
  nnd2s1 U6596 ( .DIN1(n5441), .DIN2(n6633), .Q(n6628) );
  nnd2s1 U6597 ( .DIN1(n5464), .DIN2(n5119), .Q(n6633) );
  nnd2s1 U6598 ( .DIN1(n5124), .DIN2(n6634), .Q(n6627) );
  nnd2s1 U6599 ( .DIN1(n6244), .DIN2(n6138), .Q(n6634) );
  hi1s1 U6600 ( .DIN(n5474), .Q(n6244) );
  nnd2s1 U6601 ( .DIN1(n5771), .DIN2(n5485), .Q(n5474) );
  nnd2s1 U6602 ( .DIN1(n5120), .DIN2(n5111), .Q(n6610) );
  nnd2s1 U6603 ( .DIN1(n5116), .DIN2(n5452), .Q(n6609) );
  nnd3s1 U6604 ( .DIN1(n6635), .DIN2(n6636), .DIN3(n6637), .Q(n6607) );
  nnd2s1 U6605 ( .DIN1(n5440), .DIN2(n5108), .Q(n6637) );
  or2s1 U6606 ( .DIN1(n5122), .DIN2(n5118), .Q(n6636) );
  nor2s1 U6607 ( .DIN1(n5261), .DIN2(n5265), .Q(n5118) );
  nnd2s1 U6608 ( .DIN1(n5754), .DIN2(n5128), .Q(n6635) );
  nnd4s1 U6609 ( .DIN1(n6638), .DIN2(n6639), .DIN3(n6640), .DIN4(n6641), 
        .Q(n6606) );
  nnd2s1 U6610 ( .DIN1(n6209), .DIN2(n6642), .Q(n6641) );
  nnd2s1 U6611 ( .DIN1(n6245), .DIN2(n5771), .Q(n6642) );
  nnd2s1 U6612 ( .DIN1(n5138), .DIN2(n6643), .Q(n6640) );
  nnd2s1 U6613 ( .DIN1(n5738), .DIN2(n5264), .Q(n6643) );
  nor2s1 U6614 ( .DIN1(n5107), .DIN2(n6204), .Q(n5738) );
  nnd2s1 U6615 ( .DIN1(n5139), .DIN2(n6644), .Q(n6639) );
  nnd2s1 U6616 ( .DIN1(n5140), .DIN2(n6631), .Q(n6638) );
  nnd2s1 U6617 ( .DIN1(n5775), .DIN2(n5119), .Q(n6631) );
  hi1s1 U6618 ( .DIN(n6579), .Q(n6580) );
  xor2s1 U6619 ( .DIN1(n4997), .DIN2(n6645), .Q(n6579) );
  xor2s1 U6620 ( .DIN1(n1369), .DIN2(n4910), .Q(n6645) );
  or3s1 U6621 ( .DIN1(n6646), .DIN2(n6647), .DIN3(n6648), .Q(n4910) );
  nnd4s1 U6622 ( .DIN1(n6649), .DIN2(n6650), .DIN3(n5178), .DIN4(n6651), 
        .Q(n6648) );
  and3s1 U6623 ( .DIN1(n6652), .DIN2(n6653), .DIN3(n6654), .Q(n6651) );
  nor3s1 U6624 ( .DIN1(n6655), .DIN2(n6656), .DIN3(n6657), .Q(n5178) );
  nnd4s1 U6625 ( .DIN1(n6658), .DIN2(n6659), .DIN3(n6660), .DIN4(n6661), 
        .Q(n6657) );
  and3s1 U6626 ( .DIN1(n6662), .DIN2(n6663), .DIN3(n6664), .Q(n6661) );
  nnd2s1 U6627 ( .DIN1(n5335), .DIN2(n5185), .Q(n6664) );
  nnd2s1 U6628 ( .DIN1(n5151), .DIN2(n5650), .Q(n6663) );
  nnd2s1 U6629 ( .DIN1(n5165), .DIN2(n5661), .Q(n6662) );
  nnd3s1 U6630 ( .DIN1(n6665), .DIN2(n6666), .DIN3(n6536), .Q(n6656) );
  nnd2s1 U6631 ( .DIN1(n5652), .DIN2(n6512), .Q(n6536) );
  or2s1 U6632 ( .DIN1(n5171), .DIN2(n6544), .Q(n6666) );
  nor2s1 U6633 ( .DIN1(n5182), .DIN2(n5154), .Q(n6544) );
  nnd2s1 U6634 ( .DIN1(n5685), .DIN2(n5346), .Q(n6665) );
  nnd2s1 U6635 ( .DIN1(n5676), .DIN2(n5337), .Q(n5346) );
  nnd4s1 U6636 ( .DIN1(n6667), .DIN2(n6668), .DIN3(n6669), .DIN4(n6670), 
        .Q(n6655) );
  nnd2s1 U6637 ( .DIN1(n6046), .DIN2(n6671), .Q(n6670) );
  nnd2s1 U6638 ( .DIN1(n5184), .DIN2(n6672), .Q(n6669) );
  nnd2s1 U6639 ( .DIN1(n5337), .DIN2(n5691), .Q(n6672) );
  nnd2s1 U6640 ( .DIN1(n5651), .DIN2(n6673), .Q(n6668) );
  nnd2s1 U6641 ( .DIN1(n5674), .DIN2(n5164), .Q(n6673) );
  nnd2s1 U6642 ( .DIN1(n5169), .DIN2(n6674), .Q(n6667) );
  nnd2s1 U6643 ( .DIN1(n6552), .DIN2(n6446), .Q(n6674) );
  hi1s1 U6644 ( .DIN(n5684), .Q(n6552) );
  nnd2s1 U6645 ( .DIN1(n6086), .DIN2(n5695), .Q(n5684) );
  nnd2s1 U6646 ( .DIN1(n5165), .DIN2(n5156), .Q(n6650) );
  nnd2s1 U6647 ( .DIN1(n5161), .DIN2(n5662), .Q(n6649) );
  nnd3s1 U6648 ( .DIN1(n6675), .DIN2(n6676), .DIN3(n6677), .Q(n6647) );
  nnd2s1 U6649 ( .DIN1(n5650), .DIN2(n5153), .Q(n6677) );
  or2s1 U6650 ( .DIN1(n5167), .DIN2(n5163), .Q(n6676) );
  nor2s1 U6651 ( .DIN1(n5335), .DIN2(n5339), .Q(n5163) );
  nnd2s1 U6652 ( .DIN1(n6069), .DIN2(n5173), .Q(n6675) );
  nnd4s1 U6653 ( .DIN1(n6678), .DIN2(n6679), .DIN3(n6680), .DIN4(n6681), 
        .Q(n6646) );
  nnd2s1 U6654 ( .DIN1(n6517), .DIN2(n6682), .Q(n6681) );
  nnd2s1 U6655 ( .DIN1(n6553), .DIN2(n6086), .Q(n6682) );
  nnd2s1 U6656 ( .DIN1(n5183), .DIN2(n6683), .Q(n6680) );
  nnd2s1 U6657 ( .DIN1(n6053), .DIN2(n5338), .Q(n6683) );
  nor2s1 U6658 ( .DIN1(n5152), .DIN2(n6512), .Q(n6053) );
  nnd2s1 U6659 ( .DIN1(n5184), .DIN2(n6684), .Q(n6679) );
  nnd2s1 U6660 ( .DIN1(n5185), .DIN2(n6671), .Q(n6678) );
  nnd2s1 U6661 ( .DIN1(n6090), .DIN2(n5164), .Q(n6671) );
  or3s1 U6662 ( .DIN1(n6685), .DIN2(n6686), .DIN3(n6687), .Q(n4997) );
  nnd4s1 U6663 ( .DIN1(n6416), .DIN2(n6688), .DIN3(n6689), .DIN4(n6690), 
        .Q(n6687) );
  and4s1 U6664 ( .DIN1(n6691), .DIN2(n6692), .DIN3(n6693), .DIN4(n6694), 
        .Q(n6690) );
  nnd2s1 U6665 ( .DIN1(n6020), .DIN2(n5372), .Q(n6694) );
  nnd2s1 U6666 ( .DIN1(n5627), .DIN2(n5205), .Q(n6693) );
  nnd2s1 U6667 ( .DIN1(n5388), .DIN2(n5583), .Q(n6692) );
  nor4s1 U6668 ( .DIN1(n6695), .DIN2(n6696), .DIN3(n6697), .DIN4(n6698), 
        .Q(n6416) );
  nnd4s1 U6669 ( .DIN1(n6699), .DIN2(n6700), .DIN3(n5993), .DIN4(n6701), 
        .Q(n6698) );
  nnd2s1 U6670 ( .DIN1(n5414), .DIN2(n5988), .Q(n6701) );
  nnd2s1 U6671 ( .DIN1(n5388), .DIN2(n5970), .Q(n5993) );
  nnd2s1 U6672 ( .DIN1(n5400), .DIN2(n5399), .Q(n6700) );
  nnd2s1 U6673 ( .DIN1(n5210), .DIN2(n6020), .Q(n6699) );
  nnd3s1 U6674 ( .DIN1(n6702), .DIN2(n6703), .DIN3(n6704), .Q(n6697) );
  nnd2s1 U6675 ( .DIN1(n5565), .DIN2(n6705), .Q(n6704) );
  nnd2s1 U6676 ( .DIN1(n5212), .DIN2(n5222), .Q(n6705) );
  nnd2s1 U6677 ( .DIN1(n5370), .DIN2(n6706), .Q(n6703) );
  nnd2s1 U6678 ( .DIN1(n5588), .DIN2(n5592), .Q(n6706) );
  nnd2s1 U6679 ( .DIN1(n5378), .DIN2(n6707), .Q(n6702) );
  nnd2s1 U6680 ( .DIN1(n5202), .DIN2(n5903), .Q(n6707) );
  nor2s1 U6681 ( .DIN1(n5908), .DIN2(n5390), .Q(n6696) );
  nor2s1 U6682 ( .DIN1(n5405), .DIN2(n5399), .Q(n5908) );
  nor2s1 U6683 ( .DIN1(n6708), .DIN2(n5368), .Q(n6695) );
  nor2s1 U6684 ( .DIN1(n5372), .DIN2(n5214), .Q(n6708) );
  nnd3s1 U6685 ( .DIN1(n5637), .DIN2(n6709), .DIN3(n6710), .Q(n6686) );
  nnd2s1 U6686 ( .DIN1(n5385), .DIN2(n5582), .Q(n6710) );
  nnd2s1 U6687 ( .DIN1(n5399), .DIN2(n5359), .Q(n6709) );
  nnd2s1 U6688 ( .DIN1(n5373), .DIN2(n5414), .Q(n5637) );
  nnd4s1 U6689 ( .DIN1(n6711), .DIN2(n6712), .DIN3(n6713), .DIN4(n6714), 
        .Q(n6685) );
  nnd2s1 U6690 ( .DIN1(n5210), .DIN2(n6715), .Q(n6714) );
  nnd2s1 U6691 ( .DIN1(n5588), .DIN2(n5212), .Q(n6715) );
  nnd2s1 U6692 ( .DIN1(n5568), .DIN2(n6716), .Q(n6713) );
  nnd2s1 U6693 ( .DIN1(n5564), .DIN2(n5595), .Q(n6716) );
  nnd2s1 U6694 ( .DIN1(n5358), .DIN2(n6717), .Q(n6712) );
  nnd3s1 U6695 ( .DIN1(n5571), .DIN2(n5395), .DIN3(n5202), .Q(n6717) );
  nor2s1 U6696 ( .DIN1(n5408), .DIN2(n5399), .Q(n5202) );
  nnd2s1 U6697 ( .DIN1(n5214), .DIN2(n6718), .Q(n6711) );
  nnd2s1 U6698 ( .DIN1(n6719), .DIN2(n6720), .Q(N35) );
  nnd2s1 U6699 ( .DIN1(n6721), .DIN2(n1615), .Q(n6720) );
  xor2s1 U6700 ( .DIN1(n6722), .DIN2(n6723), .Q(n6721) );
  xor2s1 U6701 ( .DIN1(n6724), .DIN2(n6725), .Q(n6723) );
  xor2s1 U6702 ( .DIN1(n5013), .DIN2(n1552), .Q(n6725) );
  hi1s1 U6703 ( .DIN(n4933), .Q(n5223) );
  or3s1 U6704 ( .DIN1(n6726), .DIN2(n6727), .DIN3(n6728), .Q(n4933) );
  nnd4s1 U6705 ( .DIN1(n6593), .DIN2(n6729), .DIN3(n6730), .DIN4(n6731), 
        .Q(n6728) );
  and3s1 U6706 ( .DIN1(n6732), .DIN2(n5803), .DIN3(n6733), .Q(n6731) );
  nnd2s1 U6707 ( .DIN1(n5510), .DIN2(n5533), .Q(n5803) );
  nnd2s1 U6708 ( .DIN1(n5841), .DIN2(n5294), .Q(n6732) );
  nor4s1 U6709 ( .DIN1(n6734), .DIN2(n6735), .DIN3(n6736), .DIN4(n6737), 
        .Q(n6593) );
  nnd4s1 U6710 ( .DIN1(n6738), .DIN2(n6370), .DIN3(n6739), .DIN4(n6740), 
        .Q(n6737) );
  nnd2s1 U6711 ( .DIN1(n5533), .DIN2(n6367), .Q(n6740) );
  nnd2s1 U6712 ( .DIN1(n5536), .DIN2(n5498), .Q(n6739) );
  nnd2s1 U6713 ( .DIN1(n6352), .DIN2(n5516), .Q(n6370) );
  nnd2s1 U6714 ( .DIN1(n5299), .DIN2(n5815), .Q(n6738) );
  nnd3s1 U6715 ( .DIN1(n6741), .DIN2(n6742), .DIN3(n6743), .Q(n6736) );
  nnd2s1 U6716 ( .DIN1(n5884), .DIN2(n6744), .Q(n6743) );
  nnd2s1 U6717 ( .DIN1(n5814), .DIN2(n6745), .Q(n6742) );
  nnd2s1 U6718 ( .DIN1(n5305), .DIN2(n5302), .Q(n6745) );
  nnd2s1 U6719 ( .DIN1(n5285), .DIN2(n6746), .Q(n6741) );
  nnd2s1 U6720 ( .DIN1(n5291), .DIN2(n6346), .Q(n6746) );
  nor2s1 U6721 ( .DIN1(n6287), .DIN2(n5518), .Q(n6735) );
  nor2s1 U6722 ( .DIN1(n5545), .DIN2(n5536), .Q(n6287) );
  nor2s1 U6723 ( .DIN1(n6747), .DIN2(n6280), .Q(n6734) );
  nor2s1 U6724 ( .DIN1(n5497), .DIN2(n5509), .Q(n6747) );
  nnd3s1 U6725 ( .DIN1(n6748), .DIN2(n6749), .DIN3(n6750), .Q(n6727) );
  nnd2s1 U6726 ( .DIN1(n5508), .DIN2(n5299), .Q(n6750) );
  nnd2s1 U6727 ( .DIN1(n5816), .DIN2(n5516), .Q(n6749) );
  nnd2s1 U6728 ( .DIN1(n5815), .DIN2(n5286), .Q(n6748) );
  nnd4s1 U6729 ( .DIN1(n6751), .DIN2(n6752), .DIN3(n6753), .DIN4(n6754), 
        .Q(n6726) );
  nnd2s1 U6730 ( .DIN1(n6347), .DIN2(n6755), .Q(n6754) );
  nnd2s1 U6731 ( .DIN1(n5857), .DIN2(n5826), .Q(n6755) );
  nnd2s1 U6732 ( .DIN1(n5884), .DIN2(n6756), .Q(n6753) );
  nnd2s1 U6733 ( .DIN1(n6280), .DIN2(n5862), .Q(n6756) );
  nnd2s1 U6734 ( .DIN1(n5509), .DIN2(n6757), .Q(n6752) );
  nnd2s1 U6735 ( .DIN1(n5507), .DIN2(n5886), .Q(n6757) );
  nor2s1 U6736 ( .DIN1(n5307), .DIN2(n5536), .Q(n5507) );
  nnd2s1 U6737 ( .DIN1(n5497), .DIN2(n6758), .Q(n6751) );
  nnd3s1 U6738 ( .DIN1(n5858), .DIN2(n5861), .DIN3(n5291), .Q(n6758) );
  nor2s1 U6739 ( .DIN1(n5542), .DIN2(n5536), .Q(n5291) );
  hi1s1 U6740 ( .DIN(n4921), .Q(n4837) );
  or3s1 U6741 ( .DIN1(n6759), .DIN2(n6760), .DIN3(n6761), .Q(n4921) );
  nnd4s1 U6742 ( .DIN1(n6614), .DIN2(n5130), .DIN3(n6762), .DIN4(n6763), 
        .Q(n6761) );
  and3s1 U6743 ( .DIN1(n6764), .DIN2(n5720), .DIN3(n6619), .Q(n6763) );
  nor2s1 U6744 ( .DIN1(n6765), .DIN2(n6766), .Q(n6619) );
  nnd4s1 U6745 ( .DIN1(n6767), .DIN2(n6768), .DIN3(n6252), .DIN4(n6769), 
        .Q(n6766) );
  nnd2s1 U6746 ( .DIN1(n5250), .DIN2(n5257), .Q(n6769) );
  nnd2s1 U6747 ( .DIN1(n5797), .DIN2(n5127), .Q(n5257) );
  nnd2s1 U6748 ( .DIN1(n5261), .DIN2(n5109), .Q(n6252) );
  nnd2s1 U6749 ( .DIN1(n5755), .DIN2(n5731), .Q(n6768) );
  nnd2s1 U6750 ( .DIN1(n5140), .DIN2(n5265), .Q(n6767) );
  nnd4s1 U6751 ( .DIN1(n6770), .DIN2(n6771), .DIN3(n6772), .DIN4(n6773), 
        .Q(n6765) );
  nnd2s1 U6752 ( .DIN1(n5110), .DIN2(n6774), .Q(n6773) );
  nnd2s1 U6753 ( .DIN1(n6146), .DIN2(n5741), .Q(n6774) );
  nnd2s1 U6754 ( .DIN1(n5472), .DIN2(n6775), .Q(n6772) );
  nnd2s1 U6755 ( .DIN1(n5466), .DIN2(n5481), .Q(n6775) );
  nnd2s1 U6756 ( .DIN1(n5442), .DIN2(n6776), .Q(n6771) );
  nnd3s1 U6757 ( .DIN1(n5254), .DIN2(n5268), .DIN3(n5264), .Q(n6776) );
  nnd2s1 U6758 ( .DIN1(n5459), .DIN2(n6777), .Q(n6770) );
  nnd4s1 U6759 ( .DIN1(n5267), .DIN2(n5449), .DIN3(n5744), .DIN4(n5466), 
        .Q(n6777) );
  nnd2s1 U6760 ( .DIN1(n5111), .DIN2(n5472), .Q(n5720) );
  nnd2s1 U6761 ( .DIN1(n5755), .DIN2(n5124), .Q(n6764) );
  nor2s1 U6762 ( .DIN1(n6778), .DIN2(n6779), .Q(n5130) );
  nnd4s1 U6763 ( .DIN1(n6780), .DIN2(n6781), .DIN3(n6782), .DIN4(n6783), 
        .Q(n6779) );
  nnd2s1 U6764 ( .DIN1(n5111), .DIN2(n5763), .Q(n6783) );
  nnd2s1 U6765 ( .DIN1(n5464), .DIN2(n5126), .Q(n5763) );
  nnd2s1 U6766 ( .DIN1(n5107), .DIN2(n5108), .Q(n6782) );
  nnd2s1 U6767 ( .DIN1(n5139), .DIN2(n5441), .Q(n6781) );
  nnd2s1 U6768 ( .DIN1(n5754), .DIN2(n5482), .Q(n6780) );
  nnd4s1 U6769 ( .DIN1(n6784), .DIN2(n6785), .DIN3(n6786), .DIN4(n6787), 
        .Q(n6778) );
  nnd2s1 U6770 ( .DIN1(n5249), .DIN2(n6788), .Q(n6787) );
  or2s1 U6771 ( .DIN1(n6255), .DIN2(n5110), .Q(n6788) );
  nnd2s1 U6772 ( .DIN1(n5452), .DIN2(n6789), .Q(n6786) );
  nnd2s1 U6773 ( .DIN1(n5254), .DIN2(n5461), .Q(n6789) );
  nnd2s1 U6774 ( .DIN1(n5140), .DIN2(n6790), .Q(n6785) );
  nnd2s1 U6775 ( .DIN1(n5779), .DIN2(n5127), .Q(n6790) );
  nnd2s1 U6776 ( .DIN1(n5124), .DIN2(n6791), .Q(n6784) );
  nnd3s1 U6777 ( .DIN1(n5775), .DIN2(n5779), .DIN3(n6792), .Q(n6791) );
  nor4s1 U6778 ( .DIN1(n6793), .DIN2(n6794), .DIN3(n6795), .DIN4(n6796), 
        .Q(n6614) );
  nnd4s1 U6779 ( .DIN1(n6797), .DIN2(n6226), .DIN3(n6798), .DIN4(n6799), 
        .Q(n6796) );
  nnd2s1 U6780 ( .DIN1(n5472), .DIN2(n5129), .Q(n6799) );
  nnd2s1 U6781 ( .DIN1(n5475), .DIN2(n5140), .Q(n6798) );
  nnd2s1 U6782 ( .DIN1(n5110), .DIN2(n6209), .Q(n6226) );
  nnd2s1 U6783 ( .DIN1(n5261), .DIN2(n5731), .Q(n6797) );
  nnd3s1 U6784 ( .DIN1(n6800), .DIN2(n6801), .DIN3(n6802), .Q(n6795) );
  nnd2s1 U6785 ( .DIN1(n5116), .DIN2(n6803), .Q(n6802) );
  nnd2s1 U6786 ( .DIN1(n5106), .DIN2(n6804), .Q(n6801) );
  nnd2s1 U6787 ( .DIN1(n5267), .DIN2(n5264), .Q(n6804) );
  nnd2s1 U6788 ( .DIN1(n5250), .DIN2(n6805), .Q(n6800) );
  nnd2s1 U6789 ( .DIN1(n5255), .DIN2(n5126), .Q(n6805) );
  nor2s1 U6790 ( .DIN1(n6145), .DIN2(n5458), .Q(n6794) );
  nor2s1 U6791 ( .DIN1(n5482), .DIN2(n5475), .Q(n6145) );
  nor2s1 U6792 ( .DIN1(n6806), .DIN2(n6139), .Q(n6793) );
  nor2s1 U6793 ( .DIN1(n5441), .DIN2(n5440), .Q(n6806) );
  nnd3s1 U6794 ( .DIN1(n6807), .DIN2(n6808), .DIN3(n6809), .Q(n6760) );
  nnd2s1 U6795 ( .DIN1(n5261), .DIN2(n5451), .Q(n6809) );
  nnd2s1 U6796 ( .DIN1(n5110), .DIN2(n5107), .Q(n6808) );
  nnd2s1 U6797 ( .DIN1(n5731), .DIN2(n5138), .Q(n6807) );
  nnd4s1 U6798 ( .DIN1(n6810), .DIN2(n6811), .DIN3(n6812), .DIN4(n6813), 
        .Q(n6759) );
  nnd2s1 U6799 ( .DIN1(n6204), .DIN2(n6814), .Q(n6813) );
  nnd2s1 U6800 ( .DIN1(n5771), .DIN2(n5740), .Q(n6814) );
  nnd2s1 U6801 ( .DIN1(n5116), .DIN2(n6815), .Q(n6812) );
  nnd2s1 U6802 ( .DIN1(n6139), .DIN2(n5775), .Q(n6815) );
  nnd2s1 U6803 ( .DIN1(n5440), .DIN2(n6816), .Q(n6811) );
  nnd2s1 U6804 ( .DIN1(n5450), .DIN2(n5797), .Q(n6816) );
  nor2s1 U6805 ( .DIN1(n5139), .DIN2(n5475), .Q(n5450) );
  nnd2s1 U6806 ( .DIN1(n5441), .DIN2(n6817), .Q(n6810) );
  nnd3s1 U6807 ( .DIN1(n5772), .DIN2(n5774), .DIN3(n5255), .Q(n6817) );
  nor2s1 U6808 ( .DIN1(n5128), .DIN2(n5475), .Q(n5255) );
  or3s1 U6809 ( .DIN1(n6818), .DIN2(n6819), .DIN3(n6820), .Q(n5013) );
  nnd4s1 U6810 ( .DIN1(n6415), .DIN2(n6821), .DIN3(n6689), .DIN4(n6822), 
        .Q(n6820) );
  and4s1 U6811 ( .DIN1(n6823), .DIN2(n6824), .DIN3(n6825), .DIN4(n6826), 
        .Q(n6822) );
  nnd2s1 U6812 ( .DIN1(n5398), .DIN2(n5385), .Q(n6826) );
  nnd2s1 U6813 ( .DIN1(n5621), .DIN2(n5414), .Q(n6825) );
  nnd2s1 U6814 ( .DIN1(n5582), .DIN2(n5357), .Q(n6824) );
  nor3s1 U6815 ( .DIN1(n6827), .DIN2(n6828), .DIN3(n6829), .Q(n6689) );
  nnd4s1 U6816 ( .DIN1(n6830), .DIN2(n6831), .DIN3(n6414), .DIN4(n6832), 
        .Q(n6829) );
  and3s1 U6817 ( .DIN1(n6833), .DIN2(n6834), .DIN3(n6835), .Q(n6832) );
  nnd2s1 U6818 ( .DIN1(n5210), .DIN2(n5583), .Q(n6835) );
  nnd2s1 U6819 ( .DIN1(n5627), .DIN2(n5568), .Q(n6834) );
  nnd2s1 U6820 ( .DIN1(n5400), .DIN2(n5385), .Q(n6833) );
  nor2s1 U6821 ( .DIN1(n6836), .DIN2(n6837), .Q(n6414) );
  nnd4s1 U6822 ( .DIN1(n6838), .DIN2(n6839), .DIN3(n6840), .DIN4(n6841), 
        .Q(n6837) );
  nnd2s1 U6823 ( .DIN1(n5210), .DIN2(n6842), .Q(n6841) );
  nnd2s1 U6824 ( .DIN1(n5904), .DIN2(n5222), .Q(n6842) );
  nnd2s1 U6825 ( .DIN1(n5357), .DIN2(n6843), .Q(n6840) );
  nnd3s1 U6826 ( .DIN1(n5221), .DIN2(n5212), .DIN3(n5203), .Q(n6843) );
  nnd2s1 U6827 ( .DIN1(n5370), .DIN2(n5398), .Q(n6839) );
  nnd2s1 U6828 ( .DIN1(n5627), .DIN2(n5359), .Q(n6838) );
  nnd4s1 U6829 ( .DIN1(n6844), .DIN2(n6845), .DIN3(n6846), .DIN4(n6847), 
        .Q(n6836) );
  nnd2s1 U6830 ( .DIN1(n5970), .DIN2(n6848), .Q(n6847) );
  nnd2s1 U6831 ( .DIN1(n5903), .DIN2(n5564), .Q(n6848) );
  nnd2s1 U6832 ( .DIN1(n5373), .DIN2(n6849), .Q(n6846) );
  nnd2s1 U6833 ( .DIN1(n5380), .DIN2(n5413), .Q(n6849) );
  nnd2s1 U6834 ( .DIN1(n5197), .DIN2(n6850), .Q(n6845) );
  nnd2s1 U6835 ( .DIN1(n5948), .DIN2(n5368), .Q(n6850) );
  nor2s1 U6836 ( .DIN1(n6020), .DIN2(n5621), .Q(n5948) );
  nnd2s1 U6837 ( .DIN1(n5388), .DIN2(n6851), .Q(n6844) );
  nnd2s1 U6838 ( .DIN1(n5222), .DIN2(n5589), .Q(n6851) );
  nnd3s1 U6839 ( .DIN1(n6852), .DIN2(n6853), .DIN3(n6854), .Q(n6828) );
  nnd2s1 U6840 ( .DIN1(n5359), .DIN2(n5414), .Q(n6854) );
  nnd2s1 U6841 ( .DIN1(n5970), .DIN2(n5565), .Q(n6853) );
  nnd2s1 U6842 ( .DIN1(n5370), .DIN2(n5378), .Q(n6852) );
  nnd4s1 U6843 ( .DIN1(n6855), .DIN2(n6856), .DIN3(n6857), .DIN4(n6858), 
        .Q(n6827) );
  nnd2s1 U6844 ( .DIN1(n5582), .DIN2(n6859), .Q(n6858) );
  nnd2s1 U6845 ( .DIN1(n5903), .DIN2(n5629), .Q(n6859) );
  nnd2s1 U6846 ( .DIN1(n5621), .DIN2(n6860), .Q(n6857) );
  nnd4s1 U6847 ( .DIN1(n5381), .DIN2(n5595), .DIN3(n5571), .DIN4(n5629), 
        .Q(n6860) );
  nnd2s1 U6848 ( .DIN1(n5405), .DIN2(n5945), .Q(n6856) );
  nnd2s1 U6849 ( .DIN1(n5588), .DIN2(n5203), .Q(n5945) );
  nnd2s1 U6850 ( .DIN1(n5197), .DIN2(n5572), .Q(n6855) );
  nnd2s1 U6851 ( .DIN1(n5201), .DIN2(n5213), .Q(n5572) );
  nor4s1 U6852 ( .DIN1(n6861), .DIN2(n6862), .DIN3(n6863), .DIN4(n6864), 
        .Q(n6415) );
  nnd4s1 U6853 ( .DIN1(n6865), .DIN2(n6866), .DIN3(n6867), .DIN4(n6868), 
        .Q(n6864) );
  nor2s1 U6854 ( .DIN1(n6869), .DIN2(n6870), .Q(n6868) );
  nor2s1 U6855 ( .DIN1(n5395), .DIN2(n5221), .Q(n6870) );
  nor2s1 U6856 ( .DIN1(n5387), .DIN2(n5563), .Q(n6869) );
  nnd2s1 U6857 ( .DIN1(n5565), .DIN2(n5398), .Q(n6867) );
  or2s1 U6858 ( .DIN1(n5381), .DIN2(n5591), .Q(n6866) );
  nor2s1 U6859 ( .DIN1(n5205), .DIN2(n6020), .Q(n5591) );
  nnd2s1 U6860 ( .DIN1(n5970), .DIN2(n5357), .Q(n6865) );
  nnd3s1 U6861 ( .DIN1(n6871), .DIN2(n6872), .DIN3(n6873), .Q(n6863) );
  nnd2s1 U6862 ( .DIN1(n5583), .DIN2(n6874), .Q(n6873) );
  nnd2s1 U6863 ( .DIN1(n5380), .DIN2(n5595), .Q(n6874) );
  nnd2s1 U6864 ( .DIN1(n5372), .DIN2(n5567), .Q(n6872) );
  nnd2s1 U6865 ( .DIN1(n5597), .DIN2(n5213), .Q(n5567) );
  nnd2s1 U6866 ( .DIN1(n5378), .DIN2(n6875), .Q(n6871) );
  nnd2s1 U6867 ( .DIN1(n5384), .DIN2(n5912), .Q(n6875) );
  nor2s1 U6868 ( .DIN1(n6876), .DIN2(n5201), .Q(n6862) );
  nor2s1 U6869 ( .DIN1(n5565), .DIN2(n5210), .Q(n6876) );
  nor2s1 U6870 ( .DIN1(n6877), .DIN2(n5212), .Q(n6861) );
  nor2s1 U6871 ( .DIN1(n5399), .DIN2(n5388), .Q(n6877) );
  nnd4s1 U6872 ( .DIN1(n5972), .DIN2(n5638), .DIN3(n6878), .DIN4(n6879), 
        .Q(n6819) );
  nnd2s1 U6873 ( .DIN1(n5358), .DIN2(n6021), .Q(n6879) );
  nnd2s1 U6874 ( .DIN1(n5405), .DIN2(n5988), .Q(n6878) );
  nnd2s1 U6875 ( .DIN1(n5399), .DIN2(n5910), .Q(n5638) );
  nnd2s1 U6876 ( .DIN1(n5370), .DIN2(n5205), .Q(n5972) );
  nnd4s1 U6877 ( .DIN1(n6880), .DIN2(n6881), .DIN3(n6882), .DIN4(n6883), 
        .Q(n6818) );
  nnd2s1 U6878 ( .DIN1(n5214), .DIN2(n6884), .Q(n6883) );
  nnd2s1 U6879 ( .DIN1(n5212), .DIN2(n5589), .Q(n6884) );
  nnd2s1 U6880 ( .DIN1(n5359), .DIN2(n6885), .Q(n6882) );
  nnd2s1 U6881 ( .DIN1(n5563), .DIN2(n5629), .Q(n6885) );
  nnd2s1 U6882 ( .DIN1(n5627), .DIN2(n5415), .Q(n6881) );
  nnd2s1 U6883 ( .DIN1(n5390), .DIN2(n5213), .Q(n5415) );
  or2s1 U6884 ( .DIN1(n5410), .DIN2(n5383), .Q(n6880) );
  nor2s1 U6885 ( .DIN1(n5366), .DIN2(n5357), .Q(n5383) );
  xor2s1 U6886 ( .DIN1(n4919), .DIN2(n6886), .Q(n6722) );
  xor2s1 U6887 ( .DIN1(n1411), .DIN2(n6887), .Q(n6886) );
  or3s1 U6888 ( .DIN1(n6888), .DIN2(n6889), .DIN3(n6890), .Q(n4919) );
  nnd4s1 U6889 ( .DIN1(n6654), .DIN2(n5175), .DIN3(n6891), .DIN4(n6892), 
        .Q(n6890) );
  and3s1 U6890 ( .DIN1(n6893), .DIN2(n6035), .DIN3(n6659), .Q(n6892) );
  nor2s1 U6891 ( .DIN1(n6894), .DIN2(n6895), .Q(n6659) );
  nnd4s1 U6892 ( .DIN1(n6896), .DIN2(n6897), .DIN3(n6560), .DIN4(n6898), 
        .Q(n6895) );
  nnd2s1 U6893 ( .DIN1(n5324), .DIN2(n5331), .Q(n6898) );
  nnd2s1 U6894 ( .DIN1(n6112), .DIN2(n5172), .Q(n5331) );
  nnd2s1 U6895 ( .DIN1(n5335), .DIN2(n5154), .Q(n6560) );
  nnd2s1 U6896 ( .DIN1(n6070), .DIN2(n6046), .Q(n6897) );
  nnd2s1 U6897 ( .DIN1(n5185), .DIN2(n5339), .Q(n6896) );
  nnd4s1 U6898 ( .DIN1(n6899), .DIN2(n6900), .DIN3(n6901), .DIN4(n6902), 
        .Q(n6894) );
  nnd2s1 U6899 ( .DIN1(n5155), .DIN2(n6903), .Q(n6902) );
  nnd2s1 U6900 ( .DIN1(n6454), .DIN2(n6056), .Q(n6903) );
  nnd2s1 U6901 ( .DIN1(n5682), .DIN2(n6904), .Q(n6901) );
  nnd2s1 U6902 ( .DIN1(n5676), .DIN2(n5691), .Q(n6904) );
  nnd2s1 U6903 ( .DIN1(n5652), .DIN2(n6905), .Q(n6900) );
  nnd3s1 U6904 ( .DIN1(n5328), .DIN2(n5342), .DIN3(n5338), .Q(n6905) );
  nnd2s1 U6905 ( .DIN1(n5669), .DIN2(n6906), .Q(n6899) );
  nnd4s1 U6906 ( .DIN1(n5341), .DIN2(n5659), .DIN3(n6059), .DIN4(n5676), 
        .Q(n6906) );
  nnd2s1 U6907 ( .DIN1(n5156), .DIN2(n5682), .Q(n6035) );
  nnd2s1 U6908 ( .DIN1(n6070), .DIN2(n5169), .Q(n6893) );
  nor2s1 U6909 ( .DIN1(n6907), .DIN2(n6908), .Q(n5175) );
  nnd4s1 U6910 ( .DIN1(n6909), .DIN2(n6910), .DIN3(n6911), .DIN4(n6912), 
        .Q(n6908) );
  nnd2s1 U6911 ( .DIN1(n5156), .DIN2(n6078), .Q(n6912) );
  nnd2s1 U6912 ( .DIN1(n5674), .DIN2(n5171), .Q(n6078) );
  nnd2s1 U6913 ( .DIN1(n5152), .DIN2(n5153), .Q(n6911) );
  nnd2s1 U6914 ( .DIN1(n5184), .DIN2(n5651), .Q(n6910) );
  nnd2s1 U6915 ( .DIN1(n6069), .DIN2(n5692), .Q(n6909) );
  nnd4s1 U6916 ( .DIN1(n6913), .DIN2(n6914), .DIN3(n6915), .DIN4(n6916), 
        .Q(n6907) );
  nnd2s1 U6917 ( .DIN1(n5323), .DIN2(n6917), .Q(n6916) );
  or2s1 U6918 ( .DIN1(n6563), .DIN2(n5155), .Q(n6917) );
  nnd2s1 U6919 ( .DIN1(n5662), .DIN2(n6918), .Q(n6915) );
  nnd2s1 U6920 ( .DIN1(n5328), .DIN2(n5671), .Q(n6918) );
  nnd2s1 U6921 ( .DIN1(n5185), .DIN2(n6919), .Q(n6914) );
  nnd2s1 U6922 ( .DIN1(n6094), .DIN2(n5172), .Q(n6919) );
  nnd2s1 U6923 ( .DIN1(n5169), .DIN2(n6920), .Q(n6913) );
  nnd3s1 U6924 ( .DIN1(n6090), .DIN2(n6094), .DIN3(n6921), .Q(n6920) );
  nor4s1 U6925 ( .DIN1(n6922), .DIN2(n6923), .DIN3(n6924), .DIN4(n6925), 
        .Q(n6654) );
  nnd4s1 U6926 ( .DIN1(n6926), .DIN2(n6534), .DIN3(n6927), .DIN4(n6928), 
        .Q(n6925) );
  nnd2s1 U6927 ( .DIN1(n5682), .DIN2(n5174), .Q(n6928) );
  nnd2s1 U6928 ( .DIN1(n5685), .DIN2(n5185), .Q(n6927) );
  nnd2s1 U6929 ( .DIN1(n5155), .DIN2(n6517), .Q(n6534) );
  nnd2s1 U6930 ( .DIN1(n5335), .DIN2(n6046), .Q(n6926) );
  nnd3s1 U6931 ( .DIN1(n6929), .DIN2(n6930), .DIN3(n6931), .Q(n6924) );
  nnd2s1 U6932 ( .DIN1(n5161), .DIN2(n6932), .Q(n6931) );
  nnd2s1 U6933 ( .DIN1(n5151), .DIN2(n6933), .Q(n6930) );
  nnd2s1 U6934 ( .DIN1(n5341), .DIN2(n5338), .Q(n6933) );
  nnd2s1 U6935 ( .DIN1(n5324), .DIN2(n6934), .Q(n6929) );
  nnd2s1 U6936 ( .DIN1(n5329), .DIN2(n5171), .Q(n6934) );
  nor2s1 U6937 ( .DIN1(n6453), .DIN2(n5668), .Q(n6923) );
  nor2s1 U6938 ( .DIN1(n5692), .DIN2(n5685), .Q(n6453) );
  nor2s1 U6939 ( .DIN1(n6935), .DIN2(n6447), .Q(n6922) );
  nor2s1 U6940 ( .DIN1(n5651), .DIN2(n5650), .Q(n6935) );
  nnd3s1 U6941 ( .DIN1(n6936), .DIN2(n6937), .DIN3(n6938), .Q(n6889) );
  nnd2s1 U6942 ( .DIN1(n5335), .DIN2(n5661), .Q(n6938) );
  nnd2s1 U6943 ( .DIN1(n5155), .DIN2(n5152), .Q(n6937) );
  nnd2s1 U6944 ( .DIN1(n6046), .DIN2(n5183), .Q(n6936) );
  nnd4s1 U6945 ( .DIN1(n6939), .DIN2(n6940), .DIN3(n6941), .DIN4(n6942), 
        .Q(n6888) );
  nnd2s1 U6946 ( .DIN1(n6512), .DIN2(n6943), .Q(n6942) );
  nnd2s1 U6947 ( .DIN1(n6086), .DIN2(n6055), .Q(n6943) );
  nnd2s1 U6948 ( .DIN1(n5161), .DIN2(n6944), .Q(n6941) );
  nnd2s1 U6949 ( .DIN1(n6447), .DIN2(n6090), .Q(n6944) );
  nnd2s1 U6950 ( .DIN1(n5650), .DIN2(n6945), .Q(n6940) );
  nnd2s1 U6951 ( .DIN1(n5660), .DIN2(n6112), .Q(n6945) );
  nor2s1 U6952 ( .DIN1(n5184), .DIN2(n5685), .Q(n5660) );
  nnd2s1 U6953 ( .DIN1(n5651), .DIN2(n6946), .Q(n6939) );
  nnd3s1 U6954 ( .DIN1(n6087), .DIN2(n6089), .DIN3(n5329), .Q(n6946) );
  nor2s1 U6955 ( .DIN1(n5173), .DIN2(n5685), .Q(n5329) );
  nnd2s1 U6956 ( .DIN1(n6947), .DIN2(n1605), .Q(n6719) );
  xor2s1 U6957 ( .DIN1(w3[1]), .DIN2(text_in_r[1]), .Q(n6947) );
  nnd2s1 U6958 ( .DIN1(n6948), .DIN2(n6949), .Q(N34) );
  nnd2s1 U6959 ( .DIN1(n6950), .DIN2(n1616), .Q(n6949) );
  xor2s1 U6960 ( .DIN1(n6951), .DIN2(n6952), .Q(n6950) );
  xor2s1 U6961 ( .DIN1(n1546), .DIN2(n5713), .Q(n6952) );
  hi1s1 U6962 ( .DIN(n6724), .Q(n5713) );
  xnr2s1 U6963 ( .DIN1(n4852), .DIN2(n4949), .Q(n6724) );
  nor3s1 U6964 ( .DIN1(n6953), .DIN2(n6954), .DIN3(n6955), .Q(n4949) );
  nnd4s1 U6965 ( .DIN1(n6956), .DIN2(n6957), .DIN3(n6958), .DIN4(n6959), 
        .Q(n6955) );
  and4s1 U6966 ( .DIN1(n6960), .DIN2(n6961), .DIN3(n6962), .DIN4(n6963), 
        .Q(n6959) );
  nnd2s1 U6967 ( .DIN1(n5565), .DIN2(n6964), .Q(n6963) );
  nnd2s1 U6968 ( .DIN1(n5904), .DIN2(n5203), .Q(n6964) );
  nnd2s1 U6969 ( .DIN1(n5366), .DIN2(n6965), .Q(n6962) );
  nnd2s1 U6970 ( .DIN1(n5203), .DIN2(n5592), .Q(n6965) );
  nnd2s1 U6971 ( .DIN1(n5219), .DIN2(n6966), .Q(n6961) );
  nnd2s1 U6972 ( .DIN1(n5904), .DIN2(n5588), .Q(n6966) );
  nnd2s1 U6973 ( .DIN1(n5568), .DIN2(n6967), .Q(n6960) );
  nnd2s1 U6974 ( .DIN1(n6420), .DIN2(n5412), .Q(n6967) );
  nor2s1 U6975 ( .DIN1(n5210), .DIN2(n5219), .Q(n6420) );
  nnd2s1 U6976 ( .DIN1(n5400), .DIN2(n5214), .Q(n6958) );
  nnd2s1 U6977 ( .DIN1(n5408), .DIN2(n5988), .Q(n6957) );
  nnd2s1 U6978 ( .DIN1(n5597), .DIN2(n5387), .Q(n5988) );
  nnd2s1 U6979 ( .DIN1(n5398), .DIN2(n5372), .Q(n6956) );
  nnd3s1 U6980 ( .DIN1(n6830), .DIN2(n6688), .DIN3(n6821), .Q(n6954) );
  nor4s1 U6981 ( .DIN1(n6968), .DIN2(n6969), .DIN3(n6970), .DIN4(n6971), 
        .Q(n6821) );
  nnd4s1 U6982 ( .DIN1(n6972), .DIN2(n6973), .DIN3(n6974), .DIN4(n6975), 
        .Q(n6971) );
  nor2s1 U6983 ( .DIN1(n6976), .DIN2(n6977), .Q(n6975) );
  nor2s1 U6984 ( .DIN1(n5912), .DIN2(n5203), .Q(n6977) );
  nor2s1 U6985 ( .DIN1(n6010), .DIN2(n5407), .Q(n6976) );
  nor2s1 U6986 ( .DIN1(n5210), .DIN2(n5408), .Q(n6010) );
  nnd2s1 U6987 ( .DIN1(n5357), .DIN2(n5613), .Q(n6974) );
  nnd2s1 U6988 ( .DIN1(n5589), .DIN2(n5390), .Q(n5613) );
  nnd2s1 U6989 ( .DIN1(n5371), .DIN2(n6978), .Q(n6973) );
  nnd3s1 U6990 ( .DIN1(n6979), .DIN2(n5395), .DIN3(n5912), .Q(n6978) );
  nnd2s1 U6991 ( .DIN1(n5910), .DIN2(n6980), .Q(n6972) );
  nnd3s1 U6992 ( .DIN1(n5571), .DIN2(n5629), .DIN3(n5595), .Q(n6980) );
  nnd3s1 U6993 ( .DIN1(n5939), .DIN2(n5190), .DIN3(n6981), .Q(n6970) );
  nnd2s1 U6994 ( .DIN1(n5385), .DIN2(n5358), .Q(n6981) );
  nnd2s1 U6995 ( .DIN1(n5372), .DIN2(n5378), .Q(n5190) );
  nnd2s1 U6996 ( .DIN1(n5219), .DIN2(n6020), .Q(n5939) );
  nor2s1 U6997 ( .DIN1(n5904), .DIN2(n5395), .Q(n6969) );
  nor2s1 U6998 ( .DIN1(n6979), .DIN2(n5368), .Q(n6968) );
  nor2s1 U6999 ( .DIN1(n6982), .DIN2(n6983), .Q(n6688) );
  nnd4s1 U7000 ( .DIN1(n6984), .DIN2(n6985), .DIN3(n6986), .DIN4(n6987), 
        .Q(n6983) );
  nnd2s1 U7001 ( .DIN1(n5621), .DIN2(n5405), .Q(n6987) );
  nnd2s1 U7002 ( .DIN1(n6020), .DIN2(n5357), .Q(n6986) );
  nnd2s1 U7003 ( .DIN1(n5214), .DIN2(n5358), .Q(n6985) );
  nnd2s1 U7004 ( .DIN1(n5197), .DIN2(n5583), .Q(n6984) );
  nnd4s1 U7005 ( .DIN1(n6988), .DIN2(n6989), .DIN3(n6990), .DIN4(n6991), 
        .Q(n6982) );
  nnd2s1 U7006 ( .DIN1(n5400), .DIN2(n6992), .Q(n6991) );
  nnd2s1 U7007 ( .DIN1(n5629), .DIN2(n5623), .Q(n6992) );
  nnd2s1 U7008 ( .DIN1(n5196), .DIN2(n6993), .Q(n6990) );
  or2s1 U7009 ( .DIN1(n6021), .DIN2(n5388), .Q(n6993) );
  nnd2s1 U7010 ( .DIN1(n5623), .DIN2(n5564), .Q(n6021) );
  nnd2s1 U7011 ( .DIN1(n5373), .DIN2(n6994), .Q(n6989) );
  or2s1 U7012 ( .DIN1(n5614), .DIN2(n5357), .Q(n6994) );
  hi1s1 U7013 ( .DIN(n5571), .Q(n5357) );
  nnd2s1 U7014 ( .DIN1(n5903), .DIN2(n5384), .Q(n5614) );
  nnd2s1 U7015 ( .DIN1(n5205), .DIN2(n6995), .Q(n6988) );
  nnd3s1 U7016 ( .DIN1(n5564), .DIN2(n5629), .DIN3(n6996), .Q(n6995) );
  and4s1 U7017 ( .DIN1(n6997), .DIN2(n6998), .DIN3(n6999), .DIN4(n7000), 
        .Q(n6830) );
  and4s1 U7018 ( .DIN1(n7001), .DIN2(n7002), .DIN3(n7003), .DIN4(n7004), 
        .Q(n7000) );
  nnd2s1 U7019 ( .DIN1(n5398), .DIN2(n5197), .Q(n7004) );
  nnd2s1 U7020 ( .DIN1(n5196), .DIN2(n5408), .Q(n7003) );
  nnd2s1 U7021 ( .DIN1(n5214), .DIN2(n5910), .Q(n7002) );
  nnd2s1 U7022 ( .DIN1(n5565), .DIN2(n5568), .Q(n7001) );
  hi1s1 U7023 ( .DIN(n5368), .Q(n5568) );
  and3s1 U7024 ( .DIN1(n7005), .DIN2(n7006), .DIN3(n7007), .Q(n6999) );
  nnd2s1 U7025 ( .DIN1(n5359), .DIN2(n7008), .Q(n7007) );
  nnd3s1 U7026 ( .DIN1(n5413), .DIN2(n6979), .DIN3(n5571), .Q(n7008) );
  nnd2s1 U7027 ( .DIN1(n5414), .DIN2(n5964), .Q(n7006) );
  nnd2s1 U7028 ( .DIN1(n5592), .DIN2(n5407), .Q(n5964) );
  nnd2s1 U7029 ( .DIN1(n5373), .DIN2(n7009), .Q(n7005) );
  nnd2s1 U7030 ( .DIN1(n5563), .DIN2(n5381), .Q(n7009) );
  nnd2s1 U7031 ( .DIN1(n5627), .DIN2(n7010), .Q(n6998) );
  nnd4s1 U7032 ( .DIN1(n5222), .DIN2(n5410), .DIN3(n5221), .DIN4(n5212), 
        .Q(n7010) );
  nnd2s1 U7033 ( .DIN1(n5399), .DIN2(n5583), .Q(n6997) );
  nnd4s1 U7034 ( .DIN1(n6412), .DIN2(n7011), .DIN3(n7012), .DIN4(n5606), 
        .Q(n6953) );
  nnd2s1 U7035 ( .DIN1(n5385), .DIN2(n5371), .Q(n5606) );
  nnd2s1 U7036 ( .DIN1(n5388), .DIN2(n5373), .Q(n7012) );
  hi1s1 U7037 ( .DIN(n5201), .Q(n5373) );
  nnd2s1 U7038 ( .DIN1(n5197), .DIN2(n5910), .Q(n7011) );
  nor3s1 U7039 ( .DIN1(n7013), .DIN2(n7014), .DIN3(n7015), .Q(n6412) );
  nnd4s1 U7040 ( .DIN1(n6691), .DIN2(n6831), .DIN3(n6823), .DIN4(n7016), 
        .Q(n7015) );
  and4s1 U7041 ( .DIN1(n7017), .DIN2(n7018), .DIN3(n7019), .DIN4(n7020), 
        .Q(n7016) );
  nnd2s1 U7042 ( .DIN1(n5405), .DIN2(n6020), .Q(n7020) );
  hi1s1 U7043 ( .DIN(n5564), .Q(n5405) );
  nnd2s1 U7044 ( .DIN1(n5210), .DIN2(n5400), .Q(n7019) );
  nnd2s1 U7045 ( .DIN1(n5565), .DIN2(n5359), .Q(n7018) );
  hi1s1 U7046 ( .DIN(n5588), .Q(n5359) );
  nnd2s1 U7047 ( .DIN1(n5366), .DIN2(n5371), .Q(n7017) );
  hi1s1 U7048 ( .DIN(n5212), .Q(n5371) );
  nor4s1 U7049 ( .DIN1(n7021), .DIN2(n7022), .DIN3(n7023), .DIN4(n7024), 
        .Q(n6823) );
  nnd4s1 U7050 ( .DIN1(n7025), .DIN2(n7026), .DIN3(n7027), .DIN4(n7028), 
        .Q(n7024) );
  nnd2s1 U7051 ( .DIN1(n5399), .DIN2(n5582), .Q(n7028) );
  nnd2s1 U7052 ( .DIN1(n5358), .DIN2(n5372), .Q(n7027) );
  nnd2s1 U7053 ( .DIN1(n5197), .DIN2(n5378), .Q(n7026) );
  hi1s1 U7054 ( .DIN(n5395), .Q(n5197) );
  nnd2s1 U7055 ( .DIN1(n7029), .DIN2(n7030), .Q(n5395) );
  nnd2s1 U7056 ( .DIN1(n5214), .DIN2(n5205), .Q(n7025) );
  nnd3s1 U7057 ( .DIN1(n7031), .DIN2(n7032), .DIN3(n7033), .Q(n7023) );
  nnd2s1 U7058 ( .DIN1(n5400), .DIN2(n7034), .Q(n7033) );
  nnd2s1 U7059 ( .DIN1(n5413), .DIN2(n5912), .Q(n7034) );
  nnd2s1 U7060 ( .DIN1(n5370), .DIN2(n6000), .Q(n7032) );
  nnd2s1 U7061 ( .DIN1(n5410), .DIN2(n5387), .Q(n6000) );
  nnd2s1 U7062 ( .DIN1(n5398), .DIN2(n7035), .Q(n7031) );
  nnd2s1 U7063 ( .DIN1(n6996), .DIN2(n5912), .Q(n7035) );
  nor2s1 U7064 ( .DIN1(n5388), .DIN2(n5408), .Q(n6996) );
  nor2s1 U7065 ( .DIN1(n5213), .DIN2(n5629), .Q(n7022) );
  and2s1 U7066 ( .DIN1(n5219), .DIN2(n7036), .Q(n7021) );
  nnd3s1 U7067 ( .DIN1(n5410), .DIN2(n5203), .DIN3(n5222), .Q(n7036) );
  nor4s1 U7068 ( .DIN1(n7037), .DIN2(n7038), .DIN3(n7039), .DIN4(n7040), 
        .Q(n6831) );
  nnd4s1 U7069 ( .DIN1(n7041), .DIN2(n7042), .DIN3(n7043), .DIN4(n7044), 
        .Q(n7040) );
  and3s1 U7070 ( .DIN1(n7045), .DIN2(n7046), .DIN3(n7047), .Q(n7044) );
  nnd2s1 U7071 ( .DIN1(n5366), .DIN2(n6428), .Q(n7047) );
  nnd2s1 U7072 ( .DIN1(n5387), .DIN2(n5390), .Q(n6428) );
  hi1s1 U7073 ( .DIN(n5629), .Q(n5366) );
  nnd2s1 U7074 ( .DIN1(n7048), .DIN2(n7030), .Q(n5629) );
  nnd2s1 U7075 ( .DIN1(n5970), .DIN2(n7049), .Q(n7046) );
  nnd2s1 U7076 ( .DIN1(n5912), .DIN2(n5595), .Q(n7049) );
  hi1s1 U7077 ( .DIN(n5213), .Q(n5970) );
  nnd2s1 U7078 ( .DIN1(n5196), .DIN2(n7050), .Q(n7045) );
  nnd2s1 U7079 ( .DIN1(n5413), .DIN2(n5381), .Q(n7050) );
  hi1s1 U7080 ( .DIN(n5410), .Q(n5196) );
  nnd2s1 U7081 ( .DIN1(n5210), .DIN2(n5398), .Q(n7043) );
  nnd2s1 U7082 ( .DIN1(n5408), .DIN2(n7051), .Q(n7042) );
  nnd2s1 U7083 ( .DIN1(n5201), .DIN2(n5203), .Q(n7051) );
  hi1s1 U7084 ( .DIN(n6979), .Q(n5408) );
  nnd2s1 U7085 ( .DIN1(n7048), .DIN2(n7052), .Q(n6979) );
  nnd2s1 U7086 ( .DIN1(n5910), .DIN2(n7053), .Q(n7041) );
  nnd2s1 U7087 ( .DIN1(n5412), .DIN2(n5623), .Q(n7053) );
  nnd3s1 U7088 ( .DIN1(n7054), .DIN2(n7055), .DIN3(n7056), .Q(n7039) );
  nnd2s1 U7089 ( .DIN1(n5627), .DIN2(n5583), .Q(n7056) );
  hi1s1 U7090 ( .DIN(n5203), .Q(n5583) );
  nnd2s1 U7091 ( .DIN1(n7057), .DIN2(n7058), .Q(n5203) );
  nnd2s1 U7092 ( .DIN1(n5565), .DIN2(n5582), .Q(n7055) );
  hi1s1 U7093 ( .DIN(n5623), .Q(n5565) );
  nnd2s1 U7094 ( .DIN1(n5621), .DIN2(n5372), .Q(n7054) );
  hi1s1 U7095 ( .DIN(n5413), .Q(n5372) );
  hi1s1 U7096 ( .DIN(n5222), .Q(n5621) );
  nor2s1 U7097 ( .DIN1(n5212), .DIN2(n5564), .Q(n7038) );
  nnd2s1 U7098 ( .DIN1(n7059), .DIN2(n7048), .Q(n5564) );
  nor2s1 U7099 ( .DIN1(n5571), .DIN2(n5904), .Q(n7037) );
  nnd2s1 U7100 ( .DIN1(n7060), .DIN2(n7052), .Q(n5571) );
  nor2s1 U7101 ( .DIN1(n7061), .DIN2(n7062), .Q(n6691) );
  nnd4s1 U7102 ( .DIN1(n5890), .DIN2(n7063), .DIN3(n7064), .DIN4(n7065), 
        .Q(n7062) );
  nnd2s1 U7103 ( .DIN1(n5388), .DIN2(n6718), .Q(n7065) );
  nnd2s1 U7104 ( .DIN1(n5588), .DIN2(n5407), .Q(n6718) );
  nnd2s1 U7105 ( .DIN1(n7066), .DIN2(n7057), .Q(n5588) );
  nnd2s1 U7106 ( .DIN1(n5627), .DIN2(n6020), .Q(n7064) );
  hi1s1 U7107 ( .DIN(n5387), .Q(n6020) );
  nnd2s1 U7108 ( .DIN1(n5400), .DIN2(n5219), .Q(n7063) );
  hi1s1 U7109 ( .DIN(n5903), .Q(n5219) );
  hi1s1 U7110 ( .DIN(n5221), .Q(n5400) );
  nnd2s1 U7111 ( .DIN1(n5210), .DIN2(n5910), .Q(n5890) );
  hi1s1 U7112 ( .DIN(n5570), .Q(n5210) );
  nnd4s1 U7113 ( .DIN1(n7067), .DIN2(n7068), .DIN3(n7069), .DIN4(n7070), 
        .Q(n7061) );
  nnd2s1 U7114 ( .DIN1(n5414), .DIN2(n7071), .Q(n7070) );
  nnd2s1 U7115 ( .DIN1(n5368), .DIN2(n5410), .Q(n7071) );
  hi1s1 U7116 ( .DIN(n5912), .Q(n5414) );
  nnd2s1 U7117 ( .DIN1(n5370), .DIN2(n7072), .Q(n7069) );
  nnd3s1 U7118 ( .DIN1(n5212), .DIN2(n5201), .DIN3(n5221), .Q(n7072) );
  nnd3s1 U7119 ( .DIN1(sa32[6]), .DIN2(sa32[7]), .DIN3(n7066), .Q(n5221) );
  nnd3s1 U7120 ( .DIN1(sa32[5]), .DIN2(sa32[4]), .DIN3(n7073), .Q(n5201) );
  nnd3s1 U7121 ( .DIN1(sa32[5]), .DIN2(n7074), .DIN3(sa32[6]), .Q(n5212) );
  nnd2s1 U7122 ( .DIN1(n5385), .DIN2(n7075), .Q(n7068) );
  nnd4s1 U7123 ( .DIN1(n5222), .DIN2(n5589), .DIN3(n5597), .DIN4(n5368), 
        .Q(n7075) );
  nnd2s1 U7124 ( .DIN1(n7066), .DIN2(n7073), .Q(n5222) );
  hi1s1 U7125 ( .DIN(n5563), .Q(n5385) );
  nnd2s1 U7126 ( .DIN1(n5378), .DIN2(n5206), .Q(n7067) );
  nnd2s1 U7127 ( .DIN1(n5570), .DIN2(n5623), .Q(n5206) );
  nnd2s1 U7128 ( .DIN1(n7076), .DIN2(n7060), .Q(n5623) );
  nnd2s1 U7129 ( .DIN1(n7059), .DIN2(n7029), .Q(n5570) );
  hi1s1 U7130 ( .DIN(n5589), .Q(n5378) );
  nnd3s1 U7131 ( .DIN1(n7074), .DIN2(n1381), .DIN3(sa32[6]), .Q(n5589) );
  nnd3s1 U7132 ( .DIN1(n5992), .DIN2(n7077), .DIN3(n7078), .Q(n7014) );
  nnd2s1 U7133 ( .DIN1(n5627), .DIN2(n5358), .Q(n7078) );
  hi1s1 U7134 ( .DIN(n5592), .Q(n5358) );
  hi1s1 U7135 ( .DIN(n5384), .Q(n5627) );
  nnd2s1 U7136 ( .DIN1(n7059), .DIN2(n7060), .Q(n5384) );
  nnd2s1 U7137 ( .DIN1(n5399), .DIN2(n5218), .Q(n7077) );
  nnd2s1 U7138 ( .DIN1(n5368), .DIN2(n5213), .Q(n5218) );
  nnd3s1 U7139 ( .DIN1(n1381), .DIN2(n1425), .DIN3(n7074), .Q(n5368) );
  hi1s1 U7140 ( .DIN(n5381), .Q(n5399) );
  nnd2s1 U7141 ( .DIN1(n7052), .DIN2(n7029), .Q(n5381) );
  nnd2s1 U7142 ( .DIN1(n5370), .DIN2(n5582), .Q(n5992) );
  hi1s1 U7143 ( .DIN(n5407), .Q(n5582) );
  nnd3s1 U7144 ( .DIN1(sa32[4]), .DIN2(n1381), .DIN3(n7057), .Q(n5407) );
  hi1s1 U7145 ( .DIN(n5595), .Q(n5370) );
  nnd2s1 U7146 ( .DIN1(n7076), .DIN2(n7048), .Q(n5595) );
  nor2s1 U7147 ( .DIN1(sa32[3]), .DIN2(sa32[1]), .Q(n7048) );
  nnd4s1 U7148 ( .DIN1(n7079), .DIN2(n7080), .DIN3(n7081), .DIN4(n7082), 
        .Q(n7013) );
  nnd2s1 U7149 ( .DIN1(n5214), .DIN2(n7083), .Q(n7082) );
  nnd2s1 U7150 ( .DIN1(n5410), .DIN2(n5213), .Q(n7083) );
  nnd3s1 U7151 ( .DIN1(sa32[7]), .DIN2(n1425), .DIN3(n7066), .Q(n5213) );
  nor2s1 U7152 ( .DIN1(sa32[5]), .DIN2(sa32[4]), .Q(n7066) );
  nnd3s1 U7153 ( .DIN1(sa32[5]), .DIN2(sa32[4]), .DIN3(n7057), .Q(n5410) );
  nor2s1 U7154 ( .DIN1(n1425), .DIN2(sa32[7]), .Q(n7057) );
  hi1s1 U7155 ( .DIN(n5380), .Q(n5214) );
  nnd2s1 U7156 ( .DIN1(n7084), .DIN2(n7030), .Q(n5380) );
  nnd2s1 U7157 ( .DIN1(n5205), .DIN2(n7085), .Q(n7081) );
  nnd2s1 U7158 ( .DIN1(n6009), .DIN2(n5912), .Q(n7085) );
  nnd2s1 U7159 ( .DIN1(n7084), .DIN2(n7052), .Q(n5912) );
  nor2s1 U7160 ( .DIN1(n1395), .DIN2(sa32[2]), .Q(n7052) );
  hi1s1 U7161 ( .DIN(n5397), .Q(n6009) );
  nnd2s1 U7162 ( .DIN1(n5563), .DIN2(n5413), .Q(n5397) );
  nnd2s1 U7163 ( .DIN1(n7076), .DIN2(n7084), .Q(n5413) );
  nnd2s1 U7164 ( .DIN1(n7059), .DIN2(n7084), .Q(n5563) );
  nor2s1 U7165 ( .DIN1(n1512), .DIN2(sa32[1]), .Q(n7084) );
  nor2s1 U7166 ( .DIN1(n1513), .DIN2(sa32[0]), .Q(n7059) );
  hi1s1 U7167 ( .DIN(n5904), .Q(n5205) );
  nnd3s1 U7168 ( .DIN1(sa32[4]), .DIN2(n1381), .DIN3(n7073), .Q(n5904) );
  nnd2s1 U7169 ( .DIN1(n5388), .DIN2(n7086), .Q(n7080) );
  nnd2s1 U7170 ( .DIN1(n5592), .DIN2(n5387), .Q(n7086) );
  nnd3s1 U7171 ( .DIN1(n7074), .DIN2(n1425), .DIN3(sa32[5]), .Q(n5387) );
  and2s1 U7172 ( .DIN1(sa32[7]), .DIN2(sa32[4]), .Q(n7074) );
  nnd3s1 U7173 ( .DIN1(sa32[7]), .DIN2(n1425), .DIN3(n7058), .Q(n5592) );
  hi1s1 U7174 ( .DIN(n5412), .Q(n5388) );
  nnd2s1 U7175 ( .DIN1(n7060), .DIN2(n7030), .Q(n5412) );
  nor2s1 U7176 ( .DIN1(sa32[2]), .DIN2(sa32[0]), .Q(n7030) );
  nor2s1 U7177 ( .DIN1(n1512), .DIN2(n1394), .Q(n7060) );
  or2s1 U7178 ( .DIN1(n5903), .DIN2(n6003), .Q(n7079) );
  nor2s1 U7179 ( .DIN1(n5910), .DIN2(n5398), .Q(n6003) );
  hi1s1 U7180 ( .DIN(n5390), .Q(n5398) );
  nnd2s1 U7181 ( .DIN1(n7073), .DIN2(n7058), .Q(n5390) );
  nor2s1 U7182 ( .DIN1(sa32[7]), .DIN2(sa32[6]), .Q(n7073) );
  hi1s1 U7183 ( .DIN(n5597), .Q(n5910) );
  nnd3s1 U7184 ( .DIN1(sa32[6]), .DIN2(sa32[7]), .DIN3(n7058), .Q(n5597) );
  nor2s1 U7185 ( .DIN1(n1381), .DIN2(sa32[4]), .Q(n7058) );
  nnd2s1 U7186 ( .DIN1(n7076), .DIN2(n7029), .Q(n5903) );
  nor2s1 U7187 ( .DIN1(n1394), .DIN2(sa32[3]), .Q(n7029) );
  nor2s1 U7188 ( .DIN1(n1513), .DIN2(n1395), .Q(n7076) );
  nor4s1 U7189 ( .DIN1(n7087), .DIN2(n7088), .DIN3(n7089), .DIN4(n7090), 
        .Q(n4852) );
  nnd4s1 U7190 ( .DIN1(n5865), .DIN2(n7091), .DIN3(n7092), .DIN4(n7093), 
        .Q(n7090) );
  nnd2s1 U7191 ( .DIN1(n5816), .DIN2(n5814), .Q(n7093) );
  nnd2s1 U7192 ( .DIN1(n5283), .DIN2(n6284), .Q(n7092) );
  nnd2s1 U7193 ( .DIN1(n5510), .DIN2(n5516), .Q(n7091) );
  nnd2s1 U7194 ( .DIN1(n5508), .DIN2(n5519), .Q(n5865) );
  nnd4s1 U7195 ( .DIN1(n7094), .DIN2(n7095), .DIN3(n7096), .DIN4(n7097), 
        .Q(n7089) );
  nnd2s1 U7196 ( .DIN1(n5884), .DIN2(n7098), .Q(n7097) );
  nnd2s1 U7197 ( .DIN1(n6597), .DIN2(n5549), .Q(n7098) );
  nor2s1 U7198 ( .DIN1(n5299), .DIN2(n5303), .Q(n6597) );
  nnd2s1 U7199 ( .DIN1(n5525), .DIN2(n7099), .Q(n7096) );
  nnd2s1 U7200 ( .DIN1(n5822), .DIN2(n5292), .Q(n7099) );
  nnd2s1 U7201 ( .DIN1(n5294), .DIN2(n7100), .Q(n7095) );
  nnd2s1 U7202 ( .DIN1(n6346), .DIN2(n5860), .Q(n7100) );
  nnd2s1 U7203 ( .DIN1(n5542), .DIN2(n6367), .Q(n7094) );
  nnd3s1 U7204 ( .DIN1(n7101), .DIN2(n6729), .DIN3(n7102), .Q(n7088) );
  nor2s1 U7205 ( .DIN1(n7103), .DIN2(n7104), .Q(n6729) );
  nnd4s1 U7206 ( .DIN1(n7105), .DIN2(n7106), .DIN3(n7107), .DIN4(n7108), 
        .Q(n7104) );
  nnd2s1 U7207 ( .DIN1(n5510), .DIN2(n5849), .Q(n7108) );
  nnd2s1 U7208 ( .DIN1(n5524), .DIN2(n6346), .Q(n5849) );
  nnd2s1 U7209 ( .DIN1(n5283), .DIN2(n5816), .Q(n7107) );
  nnd2s1 U7210 ( .DIN1(n5307), .DIN2(n5497), .Q(n7106) );
  nnd2s1 U7211 ( .DIN1(n5545), .DIN2(n5840), .Q(n7105) );
  nnd4s1 U7212 ( .DIN1(n7109), .DIN2(n7110), .DIN3(n7111), .DIN4(n7112), 
        .Q(n7103) );
  nnd2s1 U7213 ( .DIN1(n5284), .DIN2(n7113), .Q(n7112) );
  or2s1 U7214 ( .DIN1(n6399), .DIN2(n5516), .Q(n7113) );
  nnd2s1 U7215 ( .DIN1(n5511), .DIN2(n7114), .Q(n7111) );
  nnd2s1 U7216 ( .DIN1(n5290), .DIN2(n5521), .Q(n7114) );
  nnd2s1 U7217 ( .DIN1(n5498), .DIN2(n7115), .Q(n7110) );
  nnd2s1 U7218 ( .DIN1(n5867), .DIN2(n5860), .Q(n7115) );
  nnd2s1 U7219 ( .DIN1(n5294), .DIN2(n7116), .Q(n7109) );
  nnd3s1 U7220 ( .DIN1(n5862), .DIN2(n5867), .DIN3(n7117), .Q(n7116) );
  nnd4s1 U7221 ( .DIN1(n6589), .DIN2(n7118), .DIN3(n7119), .DIN4(n5496), 
        .Q(n7087) );
  nnd2s1 U7222 ( .DIN1(n5303), .DIN2(n5509), .Q(n5496) );
  nnd2s1 U7223 ( .DIN1(n5537), .DIN2(n5286), .Q(n7119) );
  nnd2s1 U7224 ( .DIN1(n5307), .DIN2(n5498), .Q(n7118) );
  nor3s1 U7225 ( .DIN1(n7120), .DIN2(n7121), .DIN3(n7122), .Q(n6589) );
  nnd4s1 U7226 ( .DIN1(n7123), .DIN2(n6733), .DIN3(n7124), .DIN4(n7125), 
        .Q(n7122) );
  and3s1 U7227 ( .DIN1(n7126), .DIN2(n7127), .DIN3(n7128), .Q(n7125) );
  nnd2s1 U7228 ( .DIN1(n5498), .DIN2(n5299), .Q(n7128) );
  nnd2s1 U7229 ( .DIN1(n5814), .DIN2(n5509), .Q(n7127) );
  nnd2s1 U7230 ( .DIN1(n5508), .DIN2(n5525), .Q(n7126) );
  nor2s1 U7231 ( .DIN1(n7129), .DIN2(n7130), .Q(n6733) );
  nnd4s1 U7232 ( .DIN1(n7131), .DIN2(n7132), .DIN3(n6396), .DIN4(n7133), 
        .Q(n7130) );
  nnd2s1 U7233 ( .DIN1(n5285), .DIN2(n5295), .Q(n7133) );
  nnd2s1 U7234 ( .DIN1(n5886), .DIN2(n5860), .Q(n5295) );
  nnd2s1 U7235 ( .DIN1(n6284), .DIN2(n5299), .Q(n6396) );
  nnd2s1 U7236 ( .DIN1(n5841), .DIN2(n5815), .Q(n7132) );
  nnd2s1 U7237 ( .DIN1(n5498), .DIN2(n5303), .Q(n7131) );
  nnd4s1 U7238 ( .DIN1(n7134), .DIN2(n7135), .DIN3(n7136), .DIN4(n7137), 
        .Q(n7129) );
  nnd2s1 U7239 ( .DIN1(n5516), .DIN2(n7138), .Q(n7137) );
  nnd2s1 U7240 ( .DIN1(n6288), .DIN2(n5827), .Q(n7138) );
  nnd2s1 U7241 ( .DIN1(n5533), .DIN2(n7139), .Q(n7136) );
  nnd2s1 U7242 ( .DIN1(n5527), .DIN2(n5544), .Q(n7139) );
  nnd2s1 U7243 ( .DIN1(n5499), .DIN2(n7140), .Q(n7135) );
  nnd3s1 U7244 ( .DIN1(n5302), .DIN2(n5290), .DIN3(n5306), .Q(n7140) );
  nnd2s1 U7245 ( .DIN1(n5519), .DIN2(n7141), .Q(n7134) );
  nnd4s1 U7246 ( .DIN1(n5527), .DIN2(n5830), .DIN3(n5305), .DIN4(n5506), 
        .Q(n7141) );
  nnd3s1 U7247 ( .DIN1(n7142), .DIN2(n7143), .DIN3(n6372), .Q(n7121) );
  nnd2s1 U7248 ( .DIN1(n5499), .DIN2(n6347), .Q(n6372) );
  or2s1 U7249 ( .DIN1(n6346), .DIN2(n6380), .Q(n7143) );
  nor2s1 U7250 ( .DIN1(n5537), .DIN2(n6284), .Q(n6380) );
  nnd2s1 U7251 ( .DIN1(n5536), .DIN2(n5311), .Q(n7142) );
  nnd2s1 U7252 ( .DIN1(n5527), .DIN2(n5301), .Q(n5311) );
  nnd4s1 U7253 ( .DIN1(n7144), .DIN2(n7145), .DIN3(n7146), .DIN4(n7147), 
        .Q(n7120) );
  nnd2s1 U7254 ( .DIN1(n5815), .DIN2(n6605), .Q(n7147) );
  nnd2s1 U7255 ( .DIN1(n5862), .DIN2(n5549), .Q(n6605) );
  nnd2s1 U7256 ( .DIN1(n5307), .DIN2(n7148), .Q(n7146) );
  nnd2s1 U7257 ( .DIN1(n5301), .DIN2(n5544), .Q(n7148) );
  nnd2s1 U7258 ( .DIN1(n5497), .DIN2(n7149), .Q(n7145) );
  nnd2s1 U7259 ( .DIN1(n5524), .DIN2(n5549), .Q(n7149) );
  nnd2s1 U7260 ( .DIN1(n5294), .DIN2(n7150), .Q(n7144) );
  nnd2s1 U7261 ( .DIN1(n6388), .DIN2(n6279), .Q(n7150) );
  hi1s1 U7262 ( .DIN(n5535), .Q(n6388) );
  nnd2s1 U7263 ( .DIN1(n5857), .DIN2(n5548), .Q(n5535) );
  hi1s1 U7264 ( .DIN(n6887), .Q(n4941) );
  or3s1 U7265 ( .DIN1(n7151), .DIN2(n7152), .DIN3(n7153), .Q(n6887) );
  nnd4s1 U7266 ( .DIN1(n6592), .DIN2(n7102), .DIN3(n6730), .DIN4(n7154), 
        .Q(n7153) );
  and4s1 U7267 ( .DIN1(n7124), .DIN2(n7155), .DIN3(n7156), .DIN4(n7157), 
        .Q(n7154) );
  nnd2s1 U7268 ( .DIN1(n5537), .DIN2(n5519), .Q(n7157) );
  nnd2s1 U7269 ( .DIN1(n5294), .DIN2(n5499), .Q(n7156) );
  nnd2s1 U7270 ( .DIN1(n5840), .DIN2(n5533), .Q(n7155) );
  and4s1 U7271 ( .DIN1(n7158), .DIN2(n7159), .DIN3(n7160), .DIN4(n7161), 
        .Q(n7124) );
  and4s1 U7272 ( .DIN1(n7162), .DIN2(n6330), .DIN3(n7163), .DIN4(n7164), 
        .Q(n7161) );
  nnd2s1 U7273 ( .DIN1(n5536), .DIN2(n6347), .Q(n7164) );
  nnd2s1 U7274 ( .DIN1(n5283), .DIN2(n5285), .Q(n7163) );
  nnd2s1 U7275 ( .DIN1(n6352), .DIN2(n5525), .Q(n6330) );
  nnd2s1 U7276 ( .DIN1(n5307), .DIN2(n5294), .Q(n7162) );
  and3s1 U7277 ( .DIN1(n7165), .DIN2(n7166), .DIN3(n7167), .Q(n7160) );
  nnd2s1 U7278 ( .DIN1(n5533), .DIN2(n7168), .Q(n7167) );
  nnd2s1 U7279 ( .DIN1(n5306), .DIN2(n5518), .Q(n7168) );
  nnd2s1 U7280 ( .DIN1(n5286), .DIN2(n7169), .Q(n7166) );
  nnd2s1 U7281 ( .DIN1(n5822), .DIN2(n5306), .Q(n7169) );
  nnd2s1 U7282 ( .DIN1(n5499), .DIN2(n6381), .Q(n7165) );
  nnd2s1 U7283 ( .DIN1(n5521), .DIN2(n5544), .Q(n6381) );
  nnd2s1 U7284 ( .DIN1(n5303), .DIN2(n7170), .Q(n7159) );
  nnd3s1 U7285 ( .DIN1(n5544), .DIN2(n5292), .DIN3(n5305), .Q(n7170) );
  hi1s1 U7286 ( .DIN(n6346), .Q(n5303) );
  or2s1 U7287 ( .DIN1(n5518), .DIN2(n7117), .Q(n7158) );
  nor2s1 U7288 ( .DIN1(n5516), .DIN2(n5542), .Q(n7117) );
  nor3s1 U7289 ( .DIN1(n7171), .DIN2(n7172), .DIN3(n7173), .Q(n6730) );
  nnd4s1 U7290 ( .DIN1(n7101), .DIN2(n7123), .DIN3(n6591), .DIN4(n7174), 
        .Q(n7173) );
  and3s1 U7291 ( .DIN1(n7175), .DIN2(n7176), .DIN3(n7177), .Q(n7174) );
  nnd2s1 U7292 ( .DIN1(n5533), .DIN2(n5509), .Q(n7177) );
  nnd2s1 U7293 ( .DIN1(n5498), .DIN2(n5519), .Q(n7176) );
  hi1s1 U7294 ( .DIN(n5306), .Q(n5498) );
  nnd2s1 U7295 ( .DIN1(n5841), .DIN2(n5884), .Q(n7175) );
  hi1s1 U7296 ( .DIN(n5527), .Q(n5884) );
  nor4s1 U7297 ( .DIN1(n7178), .DIN2(n7179), .DIN3(n7180), .DIN4(n7181), 
        .Q(n6591) );
  nnd4s1 U7298 ( .DIN1(n7182), .DIN2(n7183), .DIN3(n6295), .DIN4(n5812), 
        .Q(n7181) );
  nnd2s1 U7299 ( .DIN1(n5285), .DIN2(n5516), .Q(n5812) );
  nnd2s1 U7300 ( .DIN1(n5537), .DIN2(n5499), .Q(n6295) );
  nnd2s1 U7301 ( .DIN1(n5294), .DIN2(n5299), .Q(n7183) );
  nnd2s1 U7302 ( .DIN1(n5841), .DIN2(n5509), .Q(n7182) );
  nnd3s1 U7303 ( .DIN1(n7184), .DIN2(n7185), .DIN3(n7186), .Q(n7180) );
  nnd2s1 U7304 ( .DIN1(n5510), .DIN2(n6744), .Q(n7186) );
  nnd2s1 U7305 ( .DIN1(n5826), .DIN2(n5548), .Q(n6744) );
  nnd2s1 U7306 ( .DIN1(n5283), .DIN2(n7187), .Q(n7185) );
  nnd2s1 U7307 ( .DIN1(n6324), .DIN2(n5527), .Q(n7187) );
  nor2s1 U7308 ( .DIN1(n5840), .DIN2(n5815), .Q(n6324) );
  nnd2s1 U7309 ( .DIN1(n6352), .DIN2(n7188), .Q(n7184) );
  nnd2s1 U7310 ( .DIN1(n5862), .DIN2(n6346), .Q(n7188) );
  and2s1 U7311 ( .DIN1(n5511), .DIN2(n7189), .Q(n7179) );
  nnd3s1 U7312 ( .DIN1(n5302), .DIN2(n5292), .DIN3(n5306), .Q(n7189) );
  nor2s1 U7313 ( .DIN1(n7190), .DIN2(n5305), .Q(n7178) );
  nor2s1 U7314 ( .DIN1(n5516), .DIN2(n5299), .Q(n7190) );
  hi1s1 U7315 ( .DIN(n5549), .Q(n5516) );
  nor4s1 U7316 ( .DIN1(n7191), .DIN2(n7192), .DIN3(n7193), .DIN4(n7194), 
        .Q(n7123) );
  nnd4s1 U7317 ( .DIN1(n7195), .DIN2(n7196), .DIN3(n7197), .DIN4(n7198), 
        .Q(n7194) );
  and3s1 U7318 ( .DIN1(n7199), .DIN2(n7200), .DIN3(n7201), .Q(n7198) );
  nnd2s1 U7319 ( .DIN1(n5814), .DIN2(n6347), .Q(n7201) );
  nnd2s1 U7320 ( .DIN1(n5816), .DIN2(n7202), .Q(n7200) );
  nnd2s1 U7321 ( .DIN1(n5524), .DIN2(n5828), .Q(n7202) );
  nnd2s1 U7322 ( .DIN1(n5525), .DIN2(n6604), .Q(n7199) );
  nnd2s1 U7323 ( .DIN1(n5518), .DIN2(n5521), .Q(n6604) );
  nnd2s1 U7324 ( .DIN1(n5286), .DIN2(n7203), .Q(n7197) );
  nnd2s1 U7325 ( .DIN1(n5305), .DIN2(n5544), .Q(n7203) );
  nnd2s1 U7326 ( .DIN1(n6284), .DIN2(n7204), .Q(n7196) );
  nnd2s1 U7327 ( .DIN1(n5549), .DIN2(n5860), .Q(n7204) );
  nnd2s1 U7328 ( .DIN1(n6352), .DIN2(n7205), .Q(n7195) );
  nnd2s1 U7329 ( .DIN1(n6279), .DIN2(n6280), .Q(n7205) );
  nnd3s1 U7330 ( .DIN1(n7206), .DIN2(n7207), .DIN3(n7208), .Q(n7193) );
  nnd2s1 U7331 ( .DIN1(n5545), .DIN2(n5508), .Q(n7208) );
  nnd2s1 U7332 ( .DIN1(n5536), .DIN2(n5284), .Q(n7207) );
  nnd2s1 U7333 ( .DIN1(n5510), .DIN2(n5542), .Q(n7206) );
  nor2s1 U7334 ( .DIN1(n6341), .DIN2(n5858), .Q(n7192) );
  nor2s1 U7335 ( .DIN1(n5518), .DIN2(n5886), .Q(n7191) );
  nor4s1 U7336 ( .DIN1(n7209), .DIN2(n7210), .DIN3(n7211), .DIN4(n7212), 
        .Q(n7101) );
  nnd4s1 U7337 ( .DIN1(n7213), .DIN2(n7214), .DIN3(n7215), .DIN4(n7216), 
        .Q(n7212) );
  nnd2s1 U7338 ( .DIN1(n5536), .DIN2(n5816), .Q(n7216) );
  nnd2s1 U7339 ( .DIN1(n5307), .DIN2(n6284), .Q(n7215) );
  nnd2s1 U7340 ( .DIN1(n5284), .DIN2(n5542), .Q(n7214) );
  hi1s1 U7341 ( .DIN(n5544), .Q(n5284) );
  nnd2s1 U7342 ( .DIN1(n5283), .DIN2(n5537), .Q(n7213) );
  nnd3s1 U7343 ( .DIN1(n7217), .DIN2(n7218), .DIN3(n7219), .Q(n7211) );
  nnd2s1 U7344 ( .DIN1(n5509), .DIN2(n7220), .Q(n7219) );
  nnd3s1 U7345 ( .DIN1(n5828), .DIN2(n5548), .DIN3(n5858), .Q(n7220) );
  nnd2s1 U7346 ( .DIN1(n5510), .DIN2(n7221), .Q(n7218) );
  nnd2s1 U7347 ( .DIN1(n5857), .DIN2(n6317), .Q(n7221) );
  hi1s1 U7348 ( .DIN(n5290), .Q(n5510) );
  nnd2s1 U7349 ( .DIN1(n5533), .DIN2(n7222), .Q(n7217) );
  nnd2s1 U7350 ( .DIN1(n5822), .DIN2(n5827), .Q(n7222) );
  nor2s1 U7351 ( .DIN1(n5860), .DIN2(n5527), .Q(n7210) );
  and2s1 U7352 ( .DIN1(n5841), .DIN2(n7223), .Q(n7209) );
  nnd4s1 U7353 ( .DIN1(n5306), .DIN2(n5302), .DIN3(n5305), .DIN4(n5544), 
        .Q(n7223) );
  nnd3s1 U7354 ( .DIN1(n7224), .DIN2(n7225), .DIN3(n7226), .Q(n7172) );
  nnd2s1 U7355 ( .DIN1(n5299), .DIN2(n5816), .Q(n7226) );
  nnd2s1 U7356 ( .DIN1(n6352), .DIN2(n5814), .Q(n7225) );
  hi1s1 U7357 ( .DIN(n5301), .Q(n6352) );
  nnd2s1 U7358 ( .DIN1(n5499), .DIN2(n5285), .Q(n7224) );
  nnd4s1 U7359 ( .DIN1(n7227), .DIN2(n7228), .DIN3(n7229), .DIN4(n7230), 
        .Q(n7171) );
  nnd2s1 U7360 ( .DIN1(n6347), .DIN2(n7231), .Q(n7230) );
  nnd2s1 U7361 ( .DIN1(n5867), .DIN2(n6346), .Q(n7231) );
  nnd2s1 U7362 ( .DIN1(n5840), .DIN2(n7232), .Q(n7229) );
  nnd4s1 U7363 ( .DIN1(n6317), .DIN2(n5858), .DIN3(n5867), .DIN4(n6280), 
        .Q(n7232) );
  hi1s1 U7364 ( .DIN(n5305), .Q(n5840) );
  nnd2s1 U7365 ( .DIN1(n7233), .DIN2(n7234), .Q(n5305) );
  nnd2s1 U7366 ( .DIN1(n5545), .DIN2(n6321), .Q(n7228) );
  nnd2s1 U7367 ( .DIN1(n6288), .DIN2(n5292), .Q(n6321) );
  nnd2s1 U7368 ( .DIN1(n5283), .DIN2(n5850), .Q(n7227) );
  nnd2s1 U7369 ( .DIN1(n5290), .DIN2(n5301), .Q(n5850) );
  nor4s1 U7370 ( .DIN1(n7235), .DIN2(n7236), .DIN3(n7237), .DIN4(n7238), 
        .Q(n7102) );
  nnd4s1 U7371 ( .DIN1(n7239), .DIN2(n7240), .DIN3(n7241), .DIN4(n7242), 
        .Q(n7238) );
  nnd2s1 U7372 ( .DIN1(n5283), .DIN2(n5294), .Q(n7242) );
  hi1s1 U7373 ( .DIN(n5861), .Q(n5283) );
  nor2s1 U7374 ( .DIN1(n7243), .DIN2(n6316), .Q(n7241) );
  nor2s1 U7375 ( .DIN1(n5521), .DIN2(n6346), .Q(n6316) );
  nnd3s1 U7376 ( .DIN1(sa03[2]), .DIN2(sa03[0]), .DIN3(n7244), .Q(n6346) );
  nor2s1 U7377 ( .DIN1(n5548), .DIN2(n5506), .Q(n7243) );
  nnd2s1 U7378 ( .DIN1(n5816), .DIN2(n5533), .Q(n7240) );
  hi1s1 U7379 ( .DIN(n6279), .Q(n5533) );
  hi1s1 U7380 ( .DIN(n5292), .Q(n5816) );
  nnd2s1 U7381 ( .DIN1(n5497), .DIN2(n5519), .Q(n7239) );
  nnd3s1 U7382 ( .DIN1(n7245), .DIN2(n7246), .DIN3(n7247), .Q(n7237) );
  nnd2s1 U7383 ( .DIN1(n5511), .DIN2(n5848), .Q(n7247) );
  nnd2s1 U7384 ( .DIN1(n5518), .DIN2(n5506), .Q(n5848) );
  nnd2s1 U7385 ( .DIN1(n6284), .DIN2(n7248), .Q(n7246) );
  nnd3s1 U7386 ( .DIN1(n5867), .DIN2(n6280), .DIN3(n5858), .Q(n7248) );
  nnd2s1 U7387 ( .DIN1(n5508), .DIN2(n7249), .Q(n7245) );
  nnd3s1 U7388 ( .DIN1(n6279), .DIN2(n5861), .DIN3(n5828), .Q(n7249) );
  nor2s1 U7389 ( .DIN1(n5828), .DIN2(n5527), .Q(n7236) );
  nnd2s1 U7390 ( .DIN1(n7250), .DIN2(n7251), .Q(n5527) );
  nor2s1 U7391 ( .DIN1(n6389), .DIN2(n5827), .Q(n7235) );
  nor2s1 U7392 ( .DIN1(n5299), .DIN2(n5542), .Q(n6389) );
  hi1s1 U7393 ( .DIN(n5828), .Q(n5542) );
  nnd3s1 U7394 ( .DIN1(n7252), .DIN2(n1388), .DIN3(sa03[0]), .Q(n5828) );
  nor4s1 U7395 ( .DIN1(n7253), .DIN2(n7254), .DIN3(n7255), .DIN4(n7256), 
        .Q(n6592) );
  nnd4s1 U7396 ( .DIN1(n7257), .DIN2(n7258), .DIN3(n7259), .DIN4(n7260), 
        .Q(n7256) );
  nor2s1 U7397 ( .DIN1(n7261), .DIN2(n7262), .Q(n7260) );
  nor2s1 U7398 ( .DIN1(n5858), .DIN2(n5301), .Q(n7262) );
  nor2s1 U7399 ( .DIN1(n5306), .DIN2(n5861), .Q(n7261) );
  nnd3s1 U7400 ( .DIN1(n1355), .DIN2(n1388), .DIN3(n7244), .Q(n5861) );
  nnd2s1 U7401 ( .DIN1(n7250), .DIN2(n7263), .Q(n5306) );
  nnd2s1 U7402 ( .DIN1(n5519), .DIN2(n5815), .Q(n7259) );
  hi1s1 U7403 ( .DIN(n5857), .Q(n5519) );
  or2s1 U7404 ( .DIN1(n6317), .DIN2(n5821), .Q(n7258) );
  nor2s1 U7405 ( .DIN1(n5294), .DIN2(n5815), .Q(n5821) );
  hi1s1 U7406 ( .DIN(n5521), .Q(n5815) );
  hi1s1 U7407 ( .DIN(n6341), .Q(n5294) );
  nnd2s1 U7408 ( .DIN1(n7251), .DIN2(n7234), .Q(n6341) );
  nnd2s1 U7409 ( .DIN1(n5537), .DIN2(n5814), .Q(n7257) );
  hi1s1 U7410 ( .DIN(n5518), .Q(n5537) );
  nnd3s1 U7411 ( .DIN1(n7264), .DIN2(n7265), .DIN3(n7266), .Q(n7255) );
  nnd2s1 U7412 ( .DIN1(n5286), .DIN2(n5883), .Q(n7266) );
  nnd2s1 U7413 ( .DIN1(n5301), .DIN2(n5830), .Q(n5883) );
  hi1s1 U7414 ( .DIN(n5548), .Q(n5286) );
  nnd3s1 U7415 ( .DIN1(sa03[0]), .DIN2(n1424), .DIN3(n7267), .Q(n5548) );
  nnd2s1 U7416 ( .DIN1(n5285), .DIN2(n7268), .Q(n7265) );
  nnd2s1 U7417 ( .DIN1(n6279), .DIN2(n5524), .Q(n7268) );
  nnd3s1 U7418 ( .DIN1(n7269), .DIN2(n1424), .DIN3(sa03[0]), .Q(n6279) );
  hi1s1 U7419 ( .DIN(n5506), .Q(n5285) );
  nnd2s1 U7420 ( .DIN1(n5508), .DIN2(n7270), .Q(n7264) );
  nnd2s1 U7421 ( .DIN1(n5549), .DIN2(n6317), .Q(n7270) );
  nnd3s1 U7422 ( .DIN1(n7269), .DIN2(n1355), .DIN3(sa03[1]), .Q(n5549) );
  hi1s1 U7423 ( .DIN(n5302), .Q(n5508) );
  nor2s1 U7424 ( .DIN1(n7271), .DIN2(n5292), .Q(n7254) );
  nnd2s1 U7425 ( .DIN1(n7263), .DIN2(n7272), .Q(n5292) );
  nor2s1 U7426 ( .DIN1(n5307), .DIN2(n5499), .Q(n7271) );
  hi1s1 U7427 ( .DIN(n6280), .Q(n5499) );
  nnd3s1 U7428 ( .DIN1(sa03[0]), .DIN2(n7252), .DIN3(sa03[2]), .Q(n6280) );
  nor2s1 U7429 ( .DIN1(n7273), .DIN2(n5290), .Q(n7253) );
  nnd2s1 U7430 ( .DIN1(n7251), .DIN2(n7272), .Q(n5290) );
  nor2s1 U7431 ( .DIN1(n5814), .DIN2(n5299), .Q(n7273) );
  hi1s1 U7432 ( .DIN(n5886), .Q(n5299) );
  nnd3s1 U7433 ( .DIN1(sa03[2]), .DIN2(n1355), .DIN3(n7244), .Q(n5886) );
  hi1s1 U7434 ( .DIN(n5860), .Q(n5814) );
  nnd4s1 U7435 ( .DIN1(n5804), .DIN2(n7274), .DIN3(n7275), .DIN4(n7276), 
        .Q(n7152) );
  nnd2s1 U7436 ( .DIN1(n5497), .DIN2(n6399), .Q(n7276) );
  nnd2s1 U7437 ( .DIN1(n5862), .DIN2(n5860), .Q(n6399) );
  nnd3s1 U7438 ( .DIN1(sa03[0]), .DIN2(sa03[1]), .DIN3(n7267), .Q(n5860) );
  hi1s1 U7439 ( .DIN(n5822), .Q(n5497) );
  nnd2s1 U7440 ( .DIN1(n7277), .DIN2(n7233), .Q(n5822) );
  nnd2s1 U7441 ( .DIN1(n5545), .DIN2(n6367), .Q(n7275) );
  nnd2s1 U7442 ( .DIN1(n5521), .DIN2(n5830), .Q(n6367) );
  nnd2s1 U7443 ( .DIN1(n7251), .DIN2(n7277), .Q(n5521) );
  nor2s1 U7444 ( .DIN1(n1396), .DIN2(sa03[6]), .Q(n7251) );
  hi1s1 U7445 ( .DIN(n5862), .Q(n5545) );
  nnd3s1 U7446 ( .DIN1(n7252), .DIN2(n1355), .DIN3(sa03[2]), .Q(n5862) );
  nnd2s1 U7447 ( .DIN1(n5511), .DIN2(n6347), .Q(n7274) );
  hi1s1 U7448 ( .DIN(n5827), .Q(n6347) );
  nnd2s1 U7449 ( .DIN1(n7234), .DIN2(n7278), .Q(n5827) );
  nnd2s1 U7450 ( .DIN1(n5536), .DIN2(n6284), .Q(n5804) );
  hi1s1 U7451 ( .DIN(n5830), .Q(n6284) );
  nnd2s1 U7452 ( .DIN1(n7277), .DIN2(n7263), .Q(n5830) );
  hi1s1 U7453 ( .DIN(n6317), .Q(n5536) );
  nnd3s1 U7454 ( .DIN1(sa03[0]), .DIN2(n1388), .DIN3(n7244), .Q(n6317) );
  nor2s1 U7455 ( .DIN1(n1424), .DIN2(sa03[3]), .Q(n7244) );
  nnd4s1 U7456 ( .DIN1(n7279), .DIN2(n7280), .DIN3(n7281), .DIN4(n7282), 
        .Q(n7151) );
  nnd2s1 U7457 ( .DIN1(n5307), .DIN2(n7283), .Q(n7282) );
  nnd2s1 U7458 ( .DIN1(n5302), .DIN2(n5506), .Q(n7283) );
  nnd2s1 U7459 ( .DIN1(n7250), .DIN2(n7278), .Q(n5506) );
  nnd2s1 U7460 ( .DIN1(n7277), .DIN2(n7278), .Q(n5302) );
  nor2s1 U7461 ( .DIN1(n1515), .DIN2(n1397), .Q(n7277) );
  hi1s1 U7462 ( .DIN(n5826), .Q(n5307) );
  nnd3s1 U7463 ( .DIN1(n1355), .DIN2(n1424), .DIN3(n7269), .Q(n5826) );
  nnd2s1 U7464 ( .DIN1(n5509), .DIN2(n7284), .Q(n7281) );
  nnd2s1 U7465 ( .DIN1(n5867), .DIN2(n5857), .Q(n7284) );
  nnd3s1 U7466 ( .DIN1(n1355), .DIN2(n1424), .DIN3(n7267), .Q(n5857) );
  hi1s1 U7467 ( .DIN(n6288), .Q(n5509) );
  nnd2s1 U7468 ( .DIN1(n7263), .DIN2(n7234), .Q(n6288) );
  nor2s1 U7469 ( .DIN1(sa03[7]), .DIN2(sa03[5]), .Q(n7234) );
  nor2s1 U7470 ( .DIN1(n1514), .DIN2(sa03[4]), .Q(n7263) );
  or2s1 U7471 ( .DIN1(n5544), .DIN2(n5523), .Q(n7280) );
  nor2s1 U7472 ( .DIN1(n5525), .DIN2(n5511), .Q(n5523) );
  hi1s1 U7473 ( .DIN(n5858), .Q(n5511) );
  nnd3s1 U7474 ( .DIN1(sa03[1]), .DIN2(n7269), .DIN3(sa03[0]), .Q(n5858) );
  nor2s1 U7475 ( .DIN1(n1508), .DIN2(sa03[2]), .Q(n7269) );
  hi1s1 U7476 ( .DIN(n5867), .Q(n5525) );
  nnd3s1 U7477 ( .DIN1(n1355), .DIN2(n1388), .DIN3(n7252), .Q(n5867) );
  nor2s1 U7478 ( .DIN1(sa03[3]), .DIN2(sa03[1]), .Q(n7252) );
  nnd2s1 U7479 ( .DIN1(n7272), .DIN2(n7278), .Q(n5544) );
  nor2s1 U7480 ( .DIN1(n1514), .DIN2(n1396), .Q(n7278) );
  nnd2s1 U7481 ( .DIN1(n5841), .DIN2(n5534), .Q(n7279) );
  nnd2s1 U7482 ( .DIN1(n5518), .DIN2(n5301), .Q(n5534) );
  nnd2s1 U7483 ( .DIN1(n7250), .DIN2(n7233), .Q(n5301) );
  nor2s1 U7484 ( .DIN1(n1515), .DIN2(sa03[5]), .Q(n7250) );
  nnd2s1 U7485 ( .DIN1(n7233), .DIN2(n7272), .Q(n5518) );
  nor2s1 U7486 ( .DIN1(n1397), .DIN2(sa03[7]), .Q(n7272) );
  nor2s1 U7487 ( .DIN1(sa03[6]), .DIN2(sa03[4]), .Q(n7233) );
  hi1s1 U7488 ( .DIN(n5524), .Q(n5841) );
  nnd3s1 U7489 ( .DIN1(sa03[1]), .DIN2(n1355), .DIN3(n7267), .Q(n5524) );
  nor2s1 U7490 ( .DIN1(n1388), .DIN2(n1508), .Q(n7267) );
  nor3s1 U7491 ( .DIN1(n7285), .DIN2(n7286), .DIN3(n7287), .Q(n4845) );
  nnd4s1 U7492 ( .DIN1(n6613), .DIN2(n5132), .DIN3(n6762), .DIN4(n7288), 
        .Q(n7287) );
  and4s1 U7493 ( .DIN1(n6620), .DIN2(n7289), .DIN3(n7290), .DIN4(n7291), 
        .Q(n7288) );
  nnd2s1 U7494 ( .DIN1(n5137), .DIN2(n5459), .Q(n7291) );
  nnd2s1 U7495 ( .DIN1(n5442), .DIN2(n5124), .Q(n7290) );
  nnd2s1 U7496 ( .DIN1(n5754), .DIN2(n5472), .Q(n7289) );
  and4s1 U7497 ( .DIN1(n7292), .DIN2(n7293), .DIN3(n7294), .DIN4(n7295), 
        .Q(n6620) );
  and4s1 U7498 ( .DIN1(n7296), .DIN2(n6188), .DIN3(n7297), .DIN4(n7298), 
        .Q(n7295) );
  nnd2s1 U7499 ( .DIN1(n5475), .DIN2(n6204), .Q(n7298) );
  nnd2s1 U7500 ( .DIN1(n5108), .DIN2(n5250), .Q(n7297) );
  nnd2s1 U7501 ( .DIN1(n5120), .DIN2(n6209), .Q(n6188) );
  nnd2s1 U7502 ( .DIN1(n5139), .DIN2(n5124), .Q(n7296) );
  and3s1 U7503 ( .DIN1(n7299), .DIN2(n7300), .DIN3(n7301), .Q(n7294) );
  nnd2s1 U7504 ( .DIN1(n5472), .DIN2(n7302), .Q(n7301) );
  nnd2s1 U7505 ( .DIN1(n5268), .DIN2(n5458), .Q(n7302) );
  nnd2s1 U7506 ( .DIN1(n5138), .DIN2(n7303), .Q(n7300) );
  nnd2s1 U7507 ( .DIN1(n5122), .DIN2(n5268), .Q(n7303) );
  nnd2s1 U7508 ( .DIN1(n5442), .DIN2(n6237), .Q(n7299) );
  nnd2s1 U7509 ( .DIN1(n5461), .DIN2(n5481), .Q(n6237) );
  nnd2s1 U7510 ( .DIN1(n5265), .DIN2(n7304), .Q(n7293) );
  nnd3s1 U7511 ( .DIN1(n5267), .DIN2(n5123), .DIN3(n5481), .Q(n7304) );
  hi1s1 U7512 ( .DIN(n5126), .Q(n5265) );
  or2s1 U7513 ( .DIN1(n5458), .DIN2(n6792), .Q(n7292) );
  nor2s1 U7514 ( .DIN1(n5110), .DIN2(n5128), .Q(n6792) );
  nor3s1 U7515 ( .DIN1(n7305), .DIN2(n7306), .DIN3(n7307), .Q(n6762) );
  nnd4s1 U7516 ( .DIN1(n5131), .DIN2(n6618), .DIN3(n6612), .DIN4(n7308), 
        .Q(n7307) );
  and3s1 U7517 ( .DIN1(n7309), .DIN2(n7310), .DIN3(n7311), .Q(n7308) );
  nnd2s1 U7518 ( .DIN1(n5440), .DIN2(n5472), .Q(n7311) );
  nnd2s1 U7519 ( .DIN1(n5140), .DIN2(n5459), .Q(n7310) );
  nnd2s1 U7520 ( .DIN1(n5755), .DIN2(n5116), .Q(n7309) );
  hi1s1 U7521 ( .DIN(n5466), .Q(n5116) );
  nor4s1 U7522 ( .DIN1(n7312), .DIN2(n7313), .DIN3(n7314), .DIN4(n7315), 
        .Q(n6612) );
  nnd4s1 U7523 ( .DIN1(n7316), .DIN2(n7317), .DIN3(n6153), .DIN4(n5729), 
        .Q(n7315) );
  nnd2s1 U7524 ( .DIN1(n5110), .DIN2(n5250), .Q(n5729) );
  nnd2s1 U7525 ( .DIN1(n5442), .DIN2(n5137), .Q(n6153) );
  nnd2s1 U7526 ( .DIN1(n5261), .DIN2(n5124), .Q(n7317) );
  nnd2s1 U7527 ( .DIN1(n5755), .DIN2(n5440), .Q(n7316) );
  nnd3s1 U7528 ( .DIN1(n7318), .DIN2(n7319), .DIN3(n7320), .Q(n7314) );
  nnd2s1 U7529 ( .DIN1(n5111), .DIN2(n6803), .Q(n7320) );
  nnd2s1 U7530 ( .DIN1(n5740), .DIN2(n5485), .Q(n6803) );
  nnd2s1 U7531 ( .DIN1(n5108), .DIN2(n7321), .Q(n7319) );
  nnd2s1 U7532 ( .DIN1(n6182), .DIN2(n5466), .Q(n7321) );
  nor2s1 U7533 ( .DIN1(n5754), .DIN2(n5731), .Q(n6182) );
  nnd2s1 U7534 ( .DIN1(n6209), .DIN2(n7322), .Q(n7318) );
  nnd2s1 U7535 ( .DIN1(n5775), .DIN2(n5126), .Q(n7322) );
  and2s1 U7536 ( .DIN1(n5452), .DIN2(n7323), .Q(n7313) );
  nnd3s1 U7537 ( .DIN1(n5123), .DIN2(n5268), .DIN3(n5264), .Q(n7323) );
  nor2s1 U7538 ( .DIN1(n7324), .DIN2(n5267), .Q(n7312) );
  nor2s1 U7539 ( .DIN1(n5110), .DIN2(n5261), .Q(n7324) );
  hi1s1 U7540 ( .DIN(n5119), .Q(n5110) );
  nor4s1 U7541 ( .DIN1(n7325), .DIN2(n7326), .DIN3(n7327), .DIN4(n7328), 
        .Q(n6618) );
  nnd4s1 U7542 ( .DIN1(n7329), .DIN2(n7330), .DIN3(n7331), .DIN4(n7332), 
        .Q(n7328) );
  and3s1 U7543 ( .DIN1(n7333), .DIN2(n7334), .DIN3(n7335), .Q(n7332) );
  nnd2s1 U7544 ( .DIN1(n5106), .DIN2(n6204), .Q(n7335) );
  nnd2s1 U7545 ( .DIN1(n5107), .DIN2(n7336), .Q(n7334) );
  nnd2s1 U7546 ( .DIN1(n5464), .DIN2(n5742), .Q(n7336) );
  nnd2s1 U7547 ( .DIN1(n5120), .DIN2(n6644), .Q(n7333) );
  nnd2s1 U7548 ( .DIN1(n5458), .DIN2(n5461), .Q(n6644) );
  nnd2s1 U7549 ( .DIN1(n5138), .DIN2(n7337), .Q(n7331) );
  nnd2s1 U7550 ( .DIN1(n5267), .DIN2(n5481), .Q(n7337) );
  nnd2s1 U7551 ( .DIN1(n5109), .DIN2(n7338), .Q(n7330) );
  nnd2s1 U7552 ( .DIN1(n5119), .DIN2(n5127), .Q(n7338) );
  nnd2s1 U7553 ( .DIN1(n6209), .DIN2(n7339), .Q(n7329) );
  nnd2s1 U7554 ( .DIN1(n6138), .DIN2(n6139), .Q(n7339) );
  nnd3s1 U7555 ( .DIN1(n7340), .DIN2(n7341), .DIN3(n7342), .Q(n7327) );
  nnd2s1 U7556 ( .DIN1(n5482), .DIN2(n5451), .Q(n7342) );
  nnd2s1 U7557 ( .DIN1(n5475), .DIN2(n5249), .Q(n7341) );
  nnd2s1 U7558 ( .DIN1(n5111), .DIN2(n5128), .Q(n7340) );
  nor2s1 U7559 ( .DIN1(n5772), .DIN2(n6199), .Q(n7326) );
  nor2s1 U7560 ( .DIN1(n5458), .DIN2(n5797), .Q(n7325) );
  nor4s1 U7561 ( .DIN1(n7343), .DIN2(n7344), .DIN3(n7345), .DIN4(n7346), 
        .Q(n5131) );
  nnd4s1 U7562 ( .DIN1(n7347), .DIN2(n7348), .DIN3(n7349), .DIN4(n7350), 
        .Q(n7346) );
  nnd2s1 U7563 ( .DIN1(n5475), .DIN2(n5107), .Q(n7350) );
  nnd2s1 U7564 ( .DIN1(n5139), .DIN2(n5109), .Q(n7349) );
  nnd2s1 U7565 ( .DIN1(n5249), .DIN2(n5128), .Q(n7348) );
  hi1s1 U7566 ( .DIN(n5481), .Q(n5249) );
  nnd2s1 U7567 ( .DIN1(n5137), .DIN2(n5108), .Q(n7347) );
  hi1s1 U7568 ( .DIN(n5458), .Q(n5137) );
  nnd3s1 U7569 ( .DIN1(n7351), .DIN2(n7352), .DIN3(n7353), .Q(n7345) );
  nnd2s1 U7570 ( .DIN1(n5440), .DIN2(n7354), .Q(n7353) );
  nnd3s1 U7571 ( .DIN1(n5742), .DIN2(n5485), .DIN3(n5772), .Q(n7354) );
  nnd2s1 U7572 ( .DIN1(n5111), .DIN2(n7355), .Q(n7352) );
  nnd2s1 U7573 ( .DIN1(n5771), .DIN2(n6175), .Q(n7355) );
  hi1s1 U7574 ( .DIN(n5254), .Q(n5111) );
  nnd2s1 U7575 ( .DIN1(n5472), .DIN2(n7356), .Q(n7351) );
  nnd2s1 U7576 ( .DIN1(n5122), .DIN2(n5741), .Q(n7356) );
  nor2s1 U7577 ( .DIN1(n5466), .DIN2(n5127), .Q(n7344) );
  and2s1 U7578 ( .DIN1(n5755), .DIN2(n7357), .Q(n7343) );
  nnd4s1 U7579 ( .DIN1(n5481), .DIN2(n5267), .DIN3(n5264), .DIN4(n5268), 
        .Q(n7357) );
  nnd3s1 U7580 ( .DIN1(n7358), .DIN2(n7359), .DIN3(n7360), .Q(n7306) );
  nnd2s1 U7581 ( .DIN1(n5261), .DIN2(n5107), .Q(n7360) );
  nnd2s1 U7582 ( .DIN1(n6209), .DIN2(n5106), .Q(n7359) );
  nnd2s1 U7583 ( .DIN1(n5442), .DIN2(n5250), .Q(n7358) );
  nnd4s1 U7584 ( .DIN1(n7361), .DIN2(n7362), .DIN3(n7363), .DIN4(n7364), 
        .Q(n7305) );
  nnd2s1 U7585 ( .DIN1(n6204), .DIN2(n7365), .Q(n7364) );
  nnd2s1 U7586 ( .DIN1(n5779), .DIN2(n5126), .Q(n7365) );
  nnd2s1 U7587 ( .DIN1(n5754), .DIN2(n7366), .Q(n7363) );
  nnd4s1 U7588 ( .DIN1(n6175), .DIN2(n6139), .DIN3(n5772), .DIN4(n5779), 
        .Q(n7366) );
  hi1s1 U7589 ( .DIN(n5267), .Q(n5754) );
  nnd2s1 U7590 ( .DIN1(n7367), .DIN2(n7368), .Q(n5267) );
  nnd2s1 U7591 ( .DIN1(n5482), .DIN2(n6179), .Q(n7362) );
  nnd2s1 U7592 ( .DIN1(n6146), .DIN2(n5123), .Q(n6179) );
  nnd2s1 U7593 ( .DIN1(n5108), .DIN2(n5764), .Q(n7361) );
  nnd2s1 U7594 ( .DIN1(n5254), .DIN2(n5263), .Q(n5764) );
  nor4s1 U7595 ( .DIN1(n7369), .DIN2(n7370), .DIN3(n7371), .DIN4(n7372), 
        .Q(n5132) );
  nnd4s1 U7596 ( .DIN1(n7373), .DIN2(n7374), .DIN3(n7375), .DIN4(n7376), 
        .Q(n7372) );
  nnd2s1 U7597 ( .DIN1(n5124), .DIN2(n5108), .Q(n7376) );
  nor2s1 U7598 ( .DIN1(n7377), .DIN2(n6174), .Q(n7375) );
  nor2s1 U7599 ( .DIN1(n5461), .DIN2(n5126), .Q(n6174) );
  nnd3s1 U7600 ( .DIN1(sa10[2]), .DIN2(sa10[0]), .DIN3(n7378), .Q(n5126) );
  nor2s1 U7601 ( .DIN1(n5449), .DIN2(n5485), .Q(n7377) );
  nnd2s1 U7602 ( .DIN1(n5107), .DIN2(n5472), .Q(n7374) );
  hi1s1 U7603 ( .DIN(n6138), .Q(n5472) );
  hi1s1 U7604 ( .DIN(n5123), .Q(n5107) );
  nnd2s1 U7605 ( .DIN1(n5459), .DIN2(n5441), .Q(n7373) );
  nnd3s1 U7606 ( .DIN1(n7379), .DIN2(n7380), .DIN3(n7381), .Q(n7371) );
  nnd2s1 U7607 ( .DIN1(n5452), .DIN2(n5762), .Q(n7381) );
  nnd2s1 U7608 ( .DIN1(n5458), .DIN2(n5449), .Q(n5762) );
  nnd2s1 U7609 ( .DIN1(n5109), .DIN2(n7382), .Q(n7380) );
  nnd3s1 U7610 ( .DIN1(n5772), .DIN2(n5779), .DIN3(n6139), .Q(n7382) );
  nnd2s1 U7611 ( .DIN1(n5451), .DIN2(n7383), .Q(n7379) );
  nnd3s1 U7612 ( .DIN1(n5742), .DIN2(n5774), .DIN3(n6138), .Q(n7383) );
  nor2s1 U7613 ( .DIN1(n5742), .DIN2(n5466), .Q(n7370) );
  nnd2s1 U7614 ( .DIN1(n7384), .DIN2(n7385), .Q(n5466) );
  nor2s1 U7615 ( .DIN1(n6245), .DIN2(n5741), .Q(n7369) );
  nor2s1 U7616 ( .DIN1(n5261), .DIN2(n5128), .Q(n6245) );
  hi1s1 U7617 ( .DIN(n5742), .Q(n5128) );
  nnd3s1 U7618 ( .DIN1(n7386), .DIN2(n1389), .DIN3(sa10[0]), .Q(n5742) );
  nor4s1 U7619 ( .DIN1(n7387), .DIN2(n7388), .DIN3(n7389), .DIN4(n7390), 
        .Q(n6613) );
  nnd4s1 U7620 ( .DIN1(n7391), .DIN2(n7392), .DIN3(n7393), .DIN4(n7394), 
        .Q(n7390) );
  nnd2s1 U7621 ( .DIN1(n5459), .DIN2(n5731), .Q(n7394) );
  hi1s1 U7622 ( .DIN(n5771), .Q(n5459) );
  nor2s1 U7623 ( .DIN1(n7395), .DIN2(n7396), .Q(n7393) );
  nor2s1 U7624 ( .DIN1(n5127), .DIN2(n5458), .Q(n7396) );
  nor2s1 U7625 ( .DIN1(n5736), .DIN2(n6175), .Q(n7395) );
  nor2s1 U7626 ( .DIN1(n5124), .DIN2(n5731), .Q(n5736) );
  hi1s1 U7627 ( .DIN(n5461), .Q(n5731) );
  hi1s1 U7628 ( .DIN(n6199), .Q(n5124) );
  nnd2s1 U7629 ( .DIN1(n7384), .DIN2(n7367), .Q(n6199) );
  nnd2s1 U7630 ( .DIN1(n5140), .DIN2(n5108), .Q(n7392) );
  hi1s1 U7631 ( .DIN(n5774), .Q(n5108) );
  nnd3s1 U7632 ( .DIN1(n1356), .DIN2(n1389), .DIN3(n7378), .Q(n5774) );
  hi1s1 U7633 ( .DIN(n5268), .Q(n5140) );
  nnd2s1 U7634 ( .DIN1(n7385), .DIN2(n7397), .Q(n5268) );
  nnd2s1 U7635 ( .DIN1(n6209), .DIN2(n5452), .Q(n7391) );
  hi1s1 U7636 ( .DIN(n5263), .Q(n6209) );
  nnd3s1 U7637 ( .DIN1(n7398), .DIN2(n7399), .DIN3(n7400), .Q(n7389) );
  nnd2s1 U7638 ( .DIN1(n5138), .DIN2(n5795), .Q(n7400) );
  nnd2s1 U7639 ( .DIN1(n5263), .DIN2(n5744), .Q(n5795) );
  hi1s1 U7640 ( .DIN(n5485), .Q(n5138) );
  nnd3s1 U7641 ( .DIN1(sa10[0]), .DIN2(n1426), .DIN3(n7401), .Q(n5485) );
  nnd2s1 U7642 ( .DIN1(n5250), .DIN2(n7402), .Q(n7399) );
  nnd2s1 U7643 ( .DIN1(n6138), .DIN2(n5464), .Q(n7402) );
  nnd3s1 U7644 ( .DIN1(n7403), .DIN2(n1426), .DIN3(sa10[0]), .Q(n6138) );
  hi1s1 U7645 ( .DIN(n5449), .Q(n5250) );
  nnd2s1 U7646 ( .DIN1(n5451), .DIN2(n7404), .Q(n7398) );
  nnd2s1 U7647 ( .DIN1(n5119), .DIN2(n6175), .Q(n7404) );
  nnd3s1 U7648 ( .DIN1(n7403), .DIN2(n1356), .DIN3(sa10[1]), .Q(n5119) );
  hi1s1 U7649 ( .DIN(n5264), .Q(n5451) );
  nor2s1 U7650 ( .DIN1(n7405), .DIN2(n5123), .Q(n7388) );
  nnd2s1 U7651 ( .DIN1(n7406), .DIN2(n7397), .Q(n5123) );
  nor2s1 U7652 ( .DIN1(n5139), .DIN2(n5442), .Q(n7405) );
  hi1s1 U7653 ( .DIN(n6139), .Q(n5442) );
  nnd3s1 U7654 ( .DIN1(sa10[0]), .DIN2(n7386), .DIN3(sa10[2]), .Q(n6139) );
  nor2s1 U7655 ( .DIN1(n7407), .DIN2(n5254), .Q(n7387) );
  nnd2s1 U7656 ( .DIN1(n7384), .DIN2(n7406), .Q(n5254) );
  nor2s1 U7657 ( .DIN1(n5106), .DIN2(n5261), .Q(n7407) );
  hi1s1 U7658 ( .DIN(n5797), .Q(n5261) );
  nnd3s1 U7659 ( .DIN1(sa10[2]), .DIN2(n1356), .DIN3(n7378), .Q(n5797) );
  hi1s1 U7660 ( .DIN(n5127), .Q(n5106) );
  nnd4s1 U7661 ( .DIN1(n5721), .DIN2(n7408), .DIN3(n7409), .DIN4(n7410), 
        .Q(n7286) );
  nnd2s1 U7662 ( .DIN1(n5441), .DIN2(n6255), .Q(n7410) );
  nnd2s1 U7663 ( .DIN1(n5775), .DIN2(n5127), .Q(n6255) );
  nnd3s1 U7664 ( .DIN1(sa10[1]), .DIN2(sa10[0]), .DIN3(n7401), .Q(n5127) );
  hi1s1 U7665 ( .DIN(n5122), .Q(n5441) );
  nnd2s1 U7666 ( .DIN1(n7368), .DIN2(n7411), .Q(n5122) );
  nnd2s1 U7667 ( .DIN1(n5482), .DIN2(n5129), .Q(n7409) );
  nnd2s1 U7668 ( .DIN1(n5461), .DIN2(n5744), .Q(n5129) );
  nnd2s1 U7669 ( .DIN1(n7384), .DIN2(n7411), .Q(n5461) );
  nor2s1 U7670 ( .DIN1(n1527), .DIN2(sa10[6]), .Q(n7384) );
  hi1s1 U7671 ( .DIN(n5775), .Q(n5482) );
  nnd3s1 U7672 ( .DIN1(n7386), .DIN2(n1356), .DIN3(sa10[2]), .Q(n5775) );
  nnd2s1 U7673 ( .DIN1(n6204), .DIN2(n5452), .Q(n7408) );
  hi1s1 U7674 ( .DIN(n5741), .Q(n6204) );
  nnd2s1 U7675 ( .DIN1(n7367), .DIN2(n7412), .Q(n5741) );
  nnd2s1 U7676 ( .DIN1(n5475), .DIN2(n5109), .Q(n5721) );
  hi1s1 U7677 ( .DIN(n5744), .Q(n5109) );
  nnd2s1 U7678 ( .DIN1(n7397), .DIN2(n7411), .Q(n5744) );
  hi1s1 U7679 ( .DIN(n6175), .Q(n5475) );
  nnd3s1 U7680 ( .DIN1(sa10[0]), .DIN2(n1389), .DIN3(n7378), .Q(n6175) );
  nor2s1 U7681 ( .DIN1(n1426), .DIN2(sa10[3]), .Q(n7378) );
  nnd4s1 U7682 ( .DIN1(n7413), .DIN2(n7414), .DIN3(n7415), .DIN4(n7416), 
        .Q(n7285) );
  nnd2s1 U7683 ( .DIN1(n5139), .DIN2(n7417), .Q(n7416) );
  nnd2s1 U7684 ( .DIN1(n5264), .DIN2(n5449), .Q(n7417) );
  nnd2s1 U7685 ( .DIN1(n7385), .DIN2(n7412), .Q(n5449) );
  nnd2s1 U7686 ( .DIN1(n7412), .DIN2(n7411), .Q(n5264) );
  nor2s1 U7687 ( .DIN1(n1516), .DIN2(n1398), .Q(n7411) );
  hi1s1 U7688 ( .DIN(n5740), .Q(n5139) );
  nnd3s1 U7689 ( .DIN1(n1356), .DIN2(n1426), .DIN3(n7403), .Q(n5740) );
  nnd2s1 U7690 ( .DIN1(n5440), .DIN2(n7418), .Q(n7415) );
  nnd2s1 U7691 ( .DIN1(n5779), .DIN2(n5771), .Q(n7418) );
  nnd3s1 U7692 ( .DIN1(n1356), .DIN2(n1426), .DIN3(n7401), .Q(n5771) );
  hi1s1 U7693 ( .DIN(n6146), .Q(n5440) );
  nnd2s1 U7694 ( .DIN1(n7367), .DIN2(n7397), .Q(n6146) );
  and2s1 U7695 ( .DIN1(sa10[6]), .DIN2(n1527), .Q(n7397) );
  nor2s1 U7696 ( .DIN1(sa10[7]), .DIN2(sa10[5]), .Q(n7367) );
  or2s1 U7697 ( .DIN1(n5481), .DIN2(n5463), .Q(n7414) );
  nor2s1 U7698 ( .DIN1(n5120), .DIN2(n5452), .Q(n5463) );
  hi1s1 U7699 ( .DIN(n5772), .Q(n5452) );
  nnd3s1 U7700 ( .DIN1(sa10[0]), .DIN2(n7403), .DIN3(sa10[1]), .Q(n5772) );
  nor2s1 U7701 ( .DIN1(n1509), .DIN2(sa10[2]), .Q(n7403) );
  hi1s1 U7702 ( .DIN(n5779), .Q(n5120) );
  nnd3s1 U7703 ( .DIN1(n1356), .DIN2(n1389), .DIN3(n7386), .Q(n5779) );
  nor2s1 U7704 ( .DIN1(sa10[3]), .DIN2(sa10[1]), .Q(n7386) );
  nnd2s1 U7705 ( .DIN1(n7406), .DIN2(n7412), .Q(n5481) );
  and2s1 U7706 ( .DIN1(sa10[4]), .DIN2(sa10[6]), .Q(n7412) );
  nnd2s1 U7707 ( .DIN1(n5755), .DIN2(n5473), .Q(n7413) );
  nnd2s1 U7708 ( .DIN1(n5458), .DIN2(n5263), .Q(n5473) );
  nnd2s1 U7709 ( .DIN1(n7368), .DIN2(n7385), .Q(n5263) );
  nor2s1 U7710 ( .DIN1(n1516), .DIN2(sa10[5]), .Q(n7385) );
  nnd2s1 U7711 ( .DIN1(n7406), .DIN2(n7368), .Q(n5458) );
  nor2s1 U7712 ( .DIN1(sa10[6]), .DIN2(sa10[4]), .Q(n7368) );
  nor2s1 U7713 ( .DIN1(n1398), .DIN2(sa10[7]), .Q(n7406) );
  hi1s1 U7714 ( .DIN(n5464), .Q(n5755) );
  nnd3s1 U7715 ( .DIN1(sa10[1]), .DIN2(n1356), .DIN3(n7401), .Q(n5464) );
  nor2s1 U7716 ( .DIN1(n1389), .DIN2(n1509), .Q(n7401) );
  xor2s1 U7717 ( .DIN1(n1556), .DIN2(n4931), .Q(n6951) );
  nor3s1 U7718 ( .DIN1(n7419), .DIN2(n7420), .DIN3(n7421), .Q(n4931) );
  nnd4s1 U7719 ( .DIN1(n6653), .DIN2(n5177), .DIN3(n6891), .DIN4(n7422), 
        .Q(n7421) );
  and4s1 U7720 ( .DIN1(n6660), .DIN2(n7423), .DIN3(n7424), .DIN4(n7425), 
        .Q(n7422) );
  nnd2s1 U7721 ( .DIN1(n5182), .DIN2(n5669), .Q(n7425) );
  nnd2s1 U7722 ( .DIN1(n5652), .DIN2(n5169), .Q(n7424) );
  nnd2s1 U7723 ( .DIN1(n6069), .DIN2(n5682), .Q(n7423) );
  and4s1 U7724 ( .DIN1(n7426), .DIN2(n7427), .DIN3(n7428), .DIN4(n7429), 
        .Q(n6660) );
  and4s1 U7725 ( .DIN1(n7430), .DIN2(n6496), .DIN3(n7431), .DIN4(n7432), 
        .Q(n7429) );
  nnd2s1 U7726 ( .DIN1(n5685), .DIN2(n6512), .Q(n7432) );
  nnd2s1 U7727 ( .DIN1(n5153), .DIN2(n5324), .Q(n7431) );
  nnd2s1 U7728 ( .DIN1(n5165), .DIN2(n6517), .Q(n6496) );
  nnd2s1 U7729 ( .DIN1(n5184), .DIN2(n5169), .Q(n7430) );
  and3s1 U7730 ( .DIN1(n7433), .DIN2(n7434), .DIN3(n7435), .Q(n7428) );
  nnd2s1 U7731 ( .DIN1(n5682), .DIN2(n7436), .Q(n7435) );
  nnd2s1 U7732 ( .DIN1(n5342), .DIN2(n5668), .Q(n7436) );
  nnd2s1 U7733 ( .DIN1(n5183), .DIN2(n7437), .Q(n7434) );
  nnd2s1 U7734 ( .DIN1(n5167), .DIN2(n5342), .Q(n7437) );
  nnd2s1 U7735 ( .DIN1(n5652), .DIN2(n6545), .Q(n7433) );
  nnd2s1 U7736 ( .DIN1(n5671), .DIN2(n5691), .Q(n6545) );
  nnd2s1 U7737 ( .DIN1(n5339), .DIN2(n7438), .Q(n7427) );
  nnd3s1 U7738 ( .DIN1(n5341), .DIN2(n5168), .DIN3(n5691), .Q(n7438) );
  hi1s1 U7739 ( .DIN(n5171), .Q(n5339) );
  or2s1 U7740 ( .DIN1(n5668), .DIN2(n6921), .Q(n7426) );
  nor2s1 U7741 ( .DIN1(n5155), .DIN2(n5173), .Q(n6921) );
  nor3s1 U7742 ( .DIN1(n7439), .DIN2(n7440), .DIN3(n7441), .Q(n6891) );
  nnd4s1 U7743 ( .DIN1(n5176), .DIN2(n6658), .DIN3(n6652), .DIN4(n7442), 
        .Q(n7441) );
  and3s1 U7744 ( .DIN1(n7443), .DIN2(n7444), .DIN3(n7445), .Q(n7442) );
  nnd2s1 U7745 ( .DIN1(n5650), .DIN2(n5682), .Q(n7445) );
  nnd2s1 U7746 ( .DIN1(n5185), .DIN2(n5669), .Q(n7444) );
  nnd2s1 U7747 ( .DIN1(n6070), .DIN2(n5161), .Q(n7443) );
  hi1s1 U7748 ( .DIN(n5676), .Q(n5161) );
  nor4s1 U7749 ( .DIN1(n7446), .DIN2(n7447), .DIN3(n7448), .DIN4(n7449), 
        .Q(n6652) );
  nnd4s1 U7750 ( .DIN1(n7450), .DIN2(n7451), .DIN3(n6461), .DIN4(n6044), 
        .Q(n7449) );
  nnd2s1 U7751 ( .DIN1(n5155), .DIN2(n5324), .Q(n6044) );
  nnd2s1 U7752 ( .DIN1(n5652), .DIN2(n5182), .Q(n6461) );
  nnd2s1 U7753 ( .DIN1(n5335), .DIN2(n5169), .Q(n7451) );
  nnd2s1 U7754 ( .DIN1(n6070), .DIN2(n5650), .Q(n7450) );
  nnd3s1 U7755 ( .DIN1(n7452), .DIN2(n7453), .DIN3(n7454), .Q(n7448) );
  nnd2s1 U7756 ( .DIN1(n5156), .DIN2(n6932), .Q(n7454) );
  nnd2s1 U7757 ( .DIN1(n6055), .DIN2(n5695), .Q(n6932) );
  nnd2s1 U7758 ( .DIN1(n5153), .DIN2(n7455), .Q(n7453) );
  nnd2s1 U7759 ( .DIN1(n6490), .DIN2(n5676), .Q(n7455) );
  nor2s1 U7760 ( .DIN1(n6069), .DIN2(n6046), .Q(n6490) );
  nnd2s1 U7761 ( .DIN1(n6517), .DIN2(n7456), .Q(n7452) );
  nnd2s1 U7762 ( .DIN1(n6090), .DIN2(n5171), .Q(n7456) );
  and2s1 U7763 ( .DIN1(n5662), .DIN2(n7457), .Q(n7447) );
  nnd3s1 U7764 ( .DIN1(n5168), .DIN2(n5342), .DIN3(n5338), .Q(n7457) );
  nor2s1 U7765 ( .DIN1(n7458), .DIN2(n5341), .Q(n7446) );
  nor2s1 U7766 ( .DIN1(n5155), .DIN2(n5335), .Q(n7458) );
  hi1s1 U7767 ( .DIN(n5164), .Q(n5155) );
  nor4s1 U7768 ( .DIN1(n7459), .DIN2(n7460), .DIN3(n7461), .DIN4(n7462), 
        .Q(n6658) );
  nnd4s1 U7769 ( .DIN1(n7463), .DIN2(n7464), .DIN3(n7465), .DIN4(n7466), 
        .Q(n7462) );
  and3s1 U7770 ( .DIN1(n7467), .DIN2(n7468), .DIN3(n7469), .Q(n7466) );
  nnd2s1 U7771 ( .DIN1(n5151), .DIN2(n6512), .Q(n7469) );
  nnd2s1 U7772 ( .DIN1(n5152), .DIN2(n7470), .Q(n7468) );
  nnd2s1 U7773 ( .DIN1(n5674), .DIN2(n6057), .Q(n7470) );
  nnd2s1 U7774 ( .DIN1(n5165), .DIN2(n6684), .Q(n7467) );
  nnd2s1 U7775 ( .DIN1(n5668), .DIN2(n5671), .Q(n6684) );
  nnd2s1 U7776 ( .DIN1(n5183), .DIN2(n7471), .Q(n7465) );
  nnd2s1 U7777 ( .DIN1(n5341), .DIN2(n5691), .Q(n7471) );
  nnd2s1 U7778 ( .DIN1(n5154), .DIN2(n7472), .Q(n7464) );
  nnd2s1 U7779 ( .DIN1(n5164), .DIN2(n5172), .Q(n7472) );
  nnd2s1 U7780 ( .DIN1(n6517), .DIN2(n7473), .Q(n7463) );
  nnd2s1 U7781 ( .DIN1(n6446), .DIN2(n6447), .Q(n7473) );
  nnd3s1 U7782 ( .DIN1(n7474), .DIN2(n7475), .DIN3(n7476), .Q(n7461) );
  nnd2s1 U7783 ( .DIN1(n5692), .DIN2(n5661), .Q(n7476) );
  nnd2s1 U7784 ( .DIN1(n5685), .DIN2(n5323), .Q(n7475) );
  nnd2s1 U7785 ( .DIN1(n5156), .DIN2(n5173), .Q(n7474) );
  nor2s1 U7786 ( .DIN1(n6087), .DIN2(n6507), .Q(n7460) );
  nor2s1 U7787 ( .DIN1(n5668), .DIN2(n6112), .Q(n7459) );
  nor4s1 U7788 ( .DIN1(n7477), .DIN2(n7478), .DIN3(n7479), .DIN4(n7480), 
        .Q(n5176) );
  nnd4s1 U7789 ( .DIN1(n7481), .DIN2(n7482), .DIN3(n7483), .DIN4(n7484), 
        .Q(n7480) );
  nnd2s1 U7790 ( .DIN1(n5685), .DIN2(n5152), .Q(n7484) );
  nnd2s1 U7791 ( .DIN1(n5184), .DIN2(n5154), .Q(n7483) );
  nnd2s1 U7792 ( .DIN1(n5323), .DIN2(n5173), .Q(n7482) );
  hi1s1 U7793 ( .DIN(n5691), .Q(n5323) );
  nnd2s1 U7794 ( .DIN1(n5182), .DIN2(n5153), .Q(n7481) );
  hi1s1 U7795 ( .DIN(n5668), .Q(n5182) );
  nnd3s1 U7796 ( .DIN1(n7485), .DIN2(n7486), .DIN3(n7487), .Q(n7479) );
  nnd2s1 U7797 ( .DIN1(n5650), .DIN2(n7488), .Q(n7487) );
  nnd3s1 U7798 ( .DIN1(n6057), .DIN2(n5695), .DIN3(n6087), .Q(n7488) );
  nnd2s1 U7799 ( .DIN1(n5156), .DIN2(n7489), .Q(n7486) );
  nnd2s1 U7800 ( .DIN1(n6086), .DIN2(n6483), .Q(n7489) );
  hi1s1 U7801 ( .DIN(n5328), .Q(n5156) );
  nnd2s1 U7802 ( .DIN1(n5682), .DIN2(n7490), .Q(n7485) );
  nnd2s1 U7803 ( .DIN1(n5167), .DIN2(n6056), .Q(n7490) );
  nor2s1 U7804 ( .DIN1(n5676), .DIN2(n5172), .Q(n7478) );
  and2s1 U7805 ( .DIN1(n6070), .DIN2(n7491), .Q(n7477) );
  nnd4s1 U7806 ( .DIN1(n5691), .DIN2(n5341), .DIN3(n5338), .DIN4(n5342), 
        .Q(n7491) );
  nnd3s1 U7807 ( .DIN1(n7492), .DIN2(n7493), .DIN3(n7494), .Q(n7440) );
  nnd2s1 U7808 ( .DIN1(n5335), .DIN2(n5152), .Q(n7494) );
  nnd2s1 U7809 ( .DIN1(n6517), .DIN2(n5151), .Q(n7493) );
  nnd2s1 U7810 ( .DIN1(n5652), .DIN2(n5324), .Q(n7492) );
  nnd4s1 U7811 ( .DIN1(n7495), .DIN2(n7496), .DIN3(n7497), .DIN4(n7498), 
        .Q(n7439) );
  nnd2s1 U7812 ( .DIN1(n6512), .DIN2(n7499), .Q(n7498) );
  nnd2s1 U7813 ( .DIN1(n6094), .DIN2(n5171), .Q(n7499) );
  nnd2s1 U7814 ( .DIN1(n6069), .DIN2(n7500), .Q(n7497) );
  nnd4s1 U7815 ( .DIN1(n6483), .DIN2(n6447), .DIN3(n6087), .DIN4(n6094), 
        .Q(n7500) );
  hi1s1 U7816 ( .DIN(n5341), .Q(n6069) );
  nnd2s1 U7817 ( .DIN1(n7501), .DIN2(n7502), .Q(n5341) );
  nnd2s1 U7818 ( .DIN1(n5692), .DIN2(n6487), .Q(n7496) );
  nnd2s1 U7819 ( .DIN1(n6454), .DIN2(n5168), .Q(n6487) );
  nnd2s1 U7820 ( .DIN1(n5153), .DIN2(n6079), .Q(n7495) );
  nnd2s1 U7821 ( .DIN1(n5328), .DIN2(n5337), .Q(n6079) );
  nor4s1 U7822 ( .DIN1(n7503), .DIN2(n7504), .DIN3(n7505), .DIN4(n7506), 
        .Q(n5177) );
  nnd4s1 U7823 ( .DIN1(n7507), .DIN2(n7508), .DIN3(n7509), .DIN4(n7510), 
        .Q(n7506) );
  nnd2s1 U7824 ( .DIN1(n5169), .DIN2(n5153), .Q(n7510) );
  nor2s1 U7825 ( .DIN1(n7511), .DIN2(n6482), .Q(n7509) );
  nor2s1 U7826 ( .DIN1(n5671), .DIN2(n5171), .Q(n6482) );
  nnd3s1 U7827 ( .DIN1(sa21[2]), .DIN2(sa21[0]), .DIN3(n7512), .Q(n5171) );
  nor2s1 U7828 ( .DIN1(n5659), .DIN2(n5695), .Q(n7511) );
  nnd2s1 U7829 ( .DIN1(n5152), .DIN2(n5682), .Q(n7508) );
  hi1s1 U7830 ( .DIN(n6446), .Q(n5682) );
  hi1s1 U7831 ( .DIN(n5168), .Q(n5152) );
  nnd2s1 U7832 ( .DIN1(n5669), .DIN2(n5651), .Q(n7507) );
  nnd3s1 U7833 ( .DIN1(n7513), .DIN2(n7514), .DIN3(n7515), .Q(n7505) );
  nnd2s1 U7834 ( .DIN1(n5662), .DIN2(n6077), .Q(n7515) );
  nnd2s1 U7835 ( .DIN1(n5668), .DIN2(n5659), .Q(n6077) );
  nnd2s1 U7836 ( .DIN1(n5154), .DIN2(n7516), .Q(n7514) );
  nnd3s1 U7837 ( .DIN1(n6087), .DIN2(n6094), .DIN3(n6447), .Q(n7516) );
  nnd2s1 U7838 ( .DIN1(n5661), .DIN2(n7517), .Q(n7513) );
  nnd3s1 U7839 ( .DIN1(n6057), .DIN2(n6089), .DIN3(n6446), .Q(n7517) );
  nor2s1 U7840 ( .DIN1(n6057), .DIN2(n5676), .Q(n7504) );
  nnd2s1 U7841 ( .DIN1(n7518), .DIN2(n7519), .Q(n5676) );
  nor2s1 U7842 ( .DIN1(n6553), .DIN2(n6056), .Q(n7503) );
  nor2s1 U7843 ( .DIN1(n5335), .DIN2(n5173), .Q(n6553) );
  hi1s1 U7844 ( .DIN(n6057), .Q(n5173) );
  nnd3s1 U7845 ( .DIN1(n7520), .DIN2(n1390), .DIN3(sa21[0]), .Q(n6057) );
  nor4s1 U7846 ( .DIN1(n7521), .DIN2(n7522), .DIN3(n7523), .DIN4(n7524), 
        .Q(n6653) );
  nnd4s1 U7847 ( .DIN1(n7525), .DIN2(n7526), .DIN3(n7527), .DIN4(n7528), 
        .Q(n7524) );
  nnd2s1 U7848 ( .DIN1(n5669), .DIN2(n6046), .Q(n7528) );
  hi1s1 U7849 ( .DIN(n6086), .Q(n5669) );
  nor2s1 U7850 ( .DIN1(n7529), .DIN2(n7530), .Q(n7527) );
  nor2s1 U7851 ( .DIN1(n5172), .DIN2(n5668), .Q(n7530) );
  nor2s1 U7852 ( .DIN1(n6051), .DIN2(n6483), .Q(n7529) );
  nor2s1 U7853 ( .DIN1(n5169), .DIN2(n6046), .Q(n6051) );
  hi1s1 U7854 ( .DIN(n5671), .Q(n6046) );
  hi1s1 U7855 ( .DIN(n6507), .Q(n5169) );
  nnd2s1 U7856 ( .DIN1(n7518), .DIN2(n7501), .Q(n6507) );
  nnd2s1 U7857 ( .DIN1(n5185), .DIN2(n5153), .Q(n7526) );
  hi1s1 U7858 ( .DIN(n6089), .Q(n5153) );
  nnd3s1 U7859 ( .DIN1(n1357), .DIN2(n1390), .DIN3(n7512), .Q(n6089) );
  hi1s1 U7860 ( .DIN(n5342), .Q(n5185) );
  nnd2s1 U7861 ( .DIN1(n7519), .DIN2(n7531), .Q(n5342) );
  nnd2s1 U7862 ( .DIN1(n6517), .DIN2(n5662), .Q(n7525) );
  hi1s1 U7863 ( .DIN(n5337), .Q(n6517) );
  nnd3s1 U7864 ( .DIN1(n7532), .DIN2(n7533), .DIN3(n7534), .Q(n7523) );
  nnd2s1 U7865 ( .DIN1(n5183), .DIN2(n6110), .Q(n7534) );
  nnd2s1 U7866 ( .DIN1(n5337), .DIN2(n6059), .Q(n6110) );
  hi1s1 U7867 ( .DIN(n5695), .Q(n5183) );
  nnd3s1 U7868 ( .DIN1(sa21[0]), .DIN2(n1427), .DIN3(n7535), .Q(n5695) );
  nnd2s1 U7869 ( .DIN1(n5324), .DIN2(n7536), .Q(n7533) );
  nnd2s1 U7870 ( .DIN1(n6446), .DIN2(n5674), .Q(n7536) );
  nnd3s1 U7871 ( .DIN1(n7537), .DIN2(n1427), .DIN3(sa21[0]), .Q(n6446) );
  hi1s1 U7872 ( .DIN(n5659), .Q(n5324) );
  nnd2s1 U7873 ( .DIN1(n5661), .DIN2(n7538), .Q(n7532) );
  nnd2s1 U7874 ( .DIN1(n5164), .DIN2(n6483), .Q(n7538) );
  nnd3s1 U7875 ( .DIN1(n7537), .DIN2(n1357), .DIN3(sa21[1]), .Q(n5164) );
  hi1s1 U7876 ( .DIN(n5338), .Q(n5661) );
  nor2s1 U7877 ( .DIN1(n7539), .DIN2(n5168), .Q(n7522) );
  nnd2s1 U7878 ( .DIN1(n7540), .DIN2(n7531), .Q(n5168) );
  nor2s1 U7879 ( .DIN1(n5184), .DIN2(n5652), .Q(n7539) );
  hi1s1 U7880 ( .DIN(n6447), .Q(n5652) );
  nnd3s1 U7881 ( .DIN1(sa21[0]), .DIN2(n7520), .DIN3(sa21[2]), .Q(n6447) );
  nor2s1 U7882 ( .DIN1(n7541), .DIN2(n5328), .Q(n7521) );
  nnd2s1 U7883 ( .DIN1(n7518), .DIN2(n7540), .Q(n5328) );
  nor2s1 U7884 ( .DIN1(n5151), .DIN2(n5335), .Q(n7541) );
  hi1s1 U7885 ( .DIN(n6112), .Q(n5335) );
  nnd3s1 U7886 ( .DIN1(sa21[2]), .DIN2(n1357), .DIN3(n7512), .Q(n6112) );
  hi1s1 U7887 ( .DIN(n5172), .Q(n5151) );
  nnd4s1 U7888 ( .DIN1(n6036), .DIN2(n7542), .DIN3(n7543), .DIN4(n7544), 
        .Q(n7420) );
  nnd2s1 U7889 ( .DIN1(n5651), .DIN2(n6563), .Q(n7544) );
  nnd2s1 U7890 ( .DIN1(n6090), .DIN2(n5172), .Q(n6563) );
  nnd3s1 U7891 ( .DIN1(sa21[1]), .DIN2(sa21[0]), .DIN3(n7535), .Q(n5172) );
  hi1s1 U7892 ( .DIN(n5167), .Q(n5651) );
  nnd2s1 U7893 ( .DIN1(n7502), .DIN2(n7545), .Q(n5167) );
  nnd2s1 U7894 ( .DIN1(n5692), .DIN2(n5174), .Q(n7543) );
  nnd2s1 U7895 ( .DIN1(n5671), .DIN2(n6059), .Q(n5174) );
  nnd2s1 U7896 ( .DIN1(n7518), .DIN2(n7545), .Q(n5671) );
  nor2s1 U7897 ( .DIN1(n1528), .DIN2(sa21[6]), .Q(n7518) );
  hi1s1 U7898 ( .DIN(n6090), .Q(n5692) );
  nnd3s1 U7899 ( .DIN1(n7520), .DIN2(n1357), .DIN3(sa21[2]), .Q(n6090) );
  nnd2s1 U7900 ( .DIN1(n6512), .DIN2(n5662), .Q(n7542) );
  hi1s1 U7901 ( .DIN(n6056), .Q(n6512) );
  nnd2s1 U7902 ( .DIN1(n7501), .DIN2(n7546), .Q(n6056) );
  nnd2s1 U7903 ( .DIN1(n5685), .DIN2(n5154), .Q(n6036) );
  hi1s1 U7904 ( .DIN(n6059), .Q(n5154) );
  nnd2s1 U7905 ( .DIN1(n7531), .DIN2(n7545), .Q(n6059) );
  hi1s1 U7906 ( .DIN(n6483), .Q(n5685) );
  nnd3s1 U7907 ( .DIN1(sa21[0]), .DIN2(n1390), .DIN3(n7512), .Q(n6483) );
  nor2s1 U7908 ( .DIN1(n1427), .DIN2(sa21[3]), .Q(n7512) );
  nnd4s1 U7909 ( .DIN1(n7547), .DIN2(n7548), .DIN3(n7549), .DIN4(n7550), 
        .Q(n7419) );
  nnd2s1 U7910 ( .DIN1(n5184), .DIN2(n7551), .Q(n7550) );
  nnd2s1 U7911 ( .DIN1(n5338), .DIN2(n5659), .Q(n7551) );
  nnd2s1 U7912 ( .DIN1(n7519), .DIN2(n7546), .Q(n5659) );
  nnd2s1 U7913 ( .DIN1(n7546), .DIN2(n7545), .Q(n5338) );
  nor2s1 U7914 ( .DIN1(n1517), .DIN2(n1399), .Q(n7545) );
  hi1s1 U7915 ( .DIN(n6055), .Q(n5184) );
  nnd3s1 U7916 ( .DIN1(n1357), .DIN2(n1427), .DIN3(n7537), .Q(n6055) );
  nnd2s1 U7917 ( .DIN1(n5650), .DIN2(n7552), .Q(n7549) );
  nnd2s1 U7918 ( .DIN1(n6094), .DIN2(n6086), .Q(n7552) );
  nnd3s1 U7919 ( .DIN1(n1357), .DIN2(n1427), .DIN3(n7535), .Q(n6086) );
  hi1s1 U7920 ( .DIN(n6454), .Q(n5650) );
  nnd2s1 U7921 ( .DIN1(n7501), .DIN2(n7531), .Q(n6454) );
  and2s1 U7922 ( .DIN1(sa21[6]), .DIN2(n1528), .Q(n7531) );
  nor2s1 U7923 ( .DIN1(sa21[7]), .DIN2(sa21[5]), .Q(n7501) );
  or2s1 U7924 ( .DIN1(n5691), .DIN2(n5673), .Q(n7548) );
  nor2s1 U7925 ( .DIN1(n5165), .DIN2(n5662), .Q(n5673) );
  hi1s1 U7926 ( .DIN(n6087), .Q(n5662) );
  nnd3s1 U7927 ( .DIN1(sa21[0]), .DIN2(n7537), .DIN3(sa21[1]), .Q(n6087) );
  nor2s1 U7928 ( .DIN1(n1510), .DIN2(sa21[2]), .Q(n7537) );
  hi1s1 U7929 ( .DIN(n6094), .Q(n5165) );
  nnd3s1 U7930 ( .DIN1(n1357), .DIN2(n1390), .DIN3(n7520), .Q(n6094) );
  nor2s1 U7931 ( .DIN1(sa21[3]), .DIN2(sa21[1]), .Q(n7520) );
  nnd2s1 U7932 ( .DIN1(n7540), .DIN2(n7546), .Q(n5691) );
  and2s1 U7933 ( .DIN1(sa21[4]), .DIN2(sa21[6]), .Q(n7546) );
  nnd2s1 U7934 ( .DIN1(n6070), .DIN2(n5683), .Q(n7547) );
  nnd2s1 U7935 ( .DIN1(n5668), .DIN2(n5337), .Q(n5683) );
  nnd2s1 U7936 ( .DIN1(n7502), .DIN2(n7519), .Q(n5337) );
  nor2s1 U7937 ( .DIN1(n1517), .DIN2(sa21[5]), .Q(n7519) );
  nnd2s1 U7938 ( .DIN1(n7540), .DIN2(n7502), .Q(n5668) );
  nor2s1 U7939 ( .DIN1(sa21[6]), .DIN2(sa21[4]), .Q(n7502) );
  nor2s1 U7940 ( .DIN1(n1399), .DIN2(sa21[7]), .Q(n7540) );
  hi1s1 U7941 ( .DIN(n5674), .Q(n6070) );
  nnd3s1 U7942 ( .DIN1(sa21[1]), .DIN2(n1357), .DIN3(n7535), .Q(n5674) );
  nor2s1 U7943 ( .DIN1(n1390), .DIN2(n1510), .Q(n7535) );
  nnd2s1 U7944 ( .DIN1(n7553), .DIN2(n1605), .Q(n6948) );
  xor2s1 U7945 ( .DIN1(n1557), .DIN2(text_in_r[0]), .Q(n7553) );
  nnd2s1 U7946 ( .DIN1(n7554), .DIN2(n7555), .Q(N281) );
  nnd2s1 U7947 ( .DIN1(n7556), .DIN2(n1616), .Q(n7555) );
  xor2s1 U7948 ( .DIN1(n7557), .DIN2(n7558), .Q(n7556) );
  xor2s1 U7949 ( .DIN1(n7559), .DIN2(n7560), .Q(n7558) );
  xor2s1 U7950 ( .DIN1(w0[31]), .DIN2(n7561), .Q(n7557) );
  nnd2s1 U7951 ( .DIN1(n7562), .DIN2(n1605), .Q(n7554) );
  xor2s1 U7952 ( .DIN1(w0[31]), .DIN2(text_in_r[127]), .Q(n7562) );
  nnd2s1 U7953 ( .DIN1(n7563), .DIN2(n7564), .Q(N280) );
  nnd2s1 U7954 ( .DIN1(n7565), .DIN2(n1616), .Q(n7564) );
  xor2s1 U7955 ( .DIN1(n7566), .DIN2(n7567), .Q(n7565) );
  xor2s1 U7956 ( .DIN1(n7568), .DIN2(n7569), .Q(n7567) );
  xor2s1 U7957 ( .DIN1(n5083), .DIN2(w0[30]), .Q(n7566) );
  nnd2s1 U7958 ( .DIN1(n7570), .DIN2(n1605), .Q(n7563) );
  xor2s1 U7959 ( .DIN1(w0[30]), .DIN2(text_in_r[126]), .Q(n7570) );
  nnd2s1 U7960 ( .DIN1(n7571), .DIN2(n7572), .Q(N279) );
  nnd2s1 U7961 ( .DIN1(n7573), .DIN2(n1617), .Q(n7572) );
  xor2s1 U7962 ( .DIN1(n7574), .DIN2(n7575), .Q(n7573) );
  xor2s1 U7963 ( .DIN1(n7576), .DIN2(n7577), .Q(n7575) );
  xor2s1 U7964 ( .DIN1(n1480), .DIN2(n5082), .Q(n7574) );
  nnd2s1 U7965 ( .DIN1(n7578), .DIN2(n1605), .Q(n7571) );
  xor2s1 U7966 ( .DIN1(w0[29]), .DIN2(text_in_r[125]), .Q(n7578) );
  nnd3s1 U7967 ( .DIN1(n7579), .DIN2(n7580), .DIN3(n7581), .Q(N278) );
  nnd2s1 U7968 ( .DIN1(n1598), .DIN2(n7582), .Q(n7581) );
  xor2s1 U7969 ( .DIN1(w0[28]), .DIN2(text_in_r[124]), .Q(n7582) );
  nnd2s1 U7970 ( .DIN1(n7583), .DIN2(n7584), .Q(n7580) );
  nnd2s1 U7971 ( .DIN1(n7585), .DIN2(n7586), .Q(n7583) );
  nnd2s1 U7972 ( .DIN1(n7587), .DIN2(n7588), .Q(n7586) );
  nnd2s1 U7973 ( .DIN1(n7589), .DIN2(n7590), .Q(n7585) );
  nnd2s1 U7974 ( .DIN1(n7591), .DIN2(n7592), .Q(n7579) );
  nnd2s1 U7975 ( .DIN1(n7593), .DIN2(n7594), .Q(n7592) );
  nnd2s1 U7976 ( .DIN1(n7589), .DIN2(n7588), .Q(n7594) );
  nnd2s1 U7977 ( .DIN1(n7590), .DIN2(n7587), .Q(n7593) );
  hi1s1 U7978 ( .DIN(n7588), .Q(n7590) );
  xor2s1 U7979 ( .DIN1(n7595), .DIN2(n7596), .Q(n7588) );
  xor2s1 U7980 ( .DIN1(n1540), .DIN2(n5081), .Q(n7595) );
  nnd3s1 U7981 ( .DIN1(n7597), .DIN2(n7598), .DIN3(n7599), .Q(N277) );
  nnd2s1 U7982 ( .DIN1(n1598), .DIN2(n7600), .Q(n7599) );
  xor2s1 U7983 ( .DIN1(w0[27]), .DIN2(text_in_r[123]), .Q(n7600) );
  nnd2s1 U7984 ( .DIN1(n7601), .DIN2(n7602), .Q(n7598) );
  nnd2s1 U7985 ( .DIN1(n7603), .DIN2(n7604), .Q(n7601) );
  nnd2s1 U7986 ( .DIN1(n7605), .DIN2(n7606), .Q(n7604) );
  nnd2s1 U7987 ( .DIN1(n7607), .DIN2(n7608), .Q(n7603) );
  nnd2s1 U7988 ( .DIN1(n7609), .DIN2(n7610), .Q(n7597) );
  nnd2s1 U7989 ( .DIN1(n7611), .DIN2(n7612), .Q(n7610) );
  nnd2s1 U7990 ( .DIN1(n7607), .DIN2(n7606), .Q(n7612) );
  nnd2s1 U7991 ( .DIN1(n7608), .DIN2(n7605), .Q(n7611) );
  hi1s1 U7992 ( .DIN(n7606), .Q(n7608) );
  xor2s1 U7993 ( .DIN1(n7613), .DIN2(n7591), .Q(n7606) );
  xor2s1 U7994 ( .DIN1(n5080), .DIN2(w0[27]), .Q(n7613) );
  nnd2s1 U7995 ( .DIN1(n7614), .DIN2(n7615), .Q(N276) );
  nnd2s1 U7996 ( .DIN1(n7616), .DIN2(n1617), .Q(n7615) );
  xor2s1 U7997 ( .DIN1(n7617), .DIN2(n7618), .Q(n7616) );
  xor2s1 U7998 ( .DIN1(n7619), .DIN2(n7620), .Q(n7618) );
  xor2s1 U7999 ( .DIN1(w0[26]), .DIN2(n7621), .Q(n7617) );
  nnd2s1 U8000 ( .DIN1(n7622), .DIN2(n1604), .Q(n7614) );
  xor2s1 U8001 ( .DIN1(w0[26]), .DIN2(text_in_r[122]), .Q(n7622) );
  nnd2s1 U8002 ( .DIN1(n7623), .DIN2(n7624), .Q(N275) );
  nnd2s1 U8003 ( .DIN1(n7625), .DIN2(n1617), .Q(n7624) );
  xor2s1 U8004 ( .DIN1(n7626), .DIN2(n7627), .Q(n7625) );
  xnr2s1 U8005 ( .DIN1(n7628), .DIN2(n7629), .Q(n7627) );
  xor2s1 U8006 ( .DIN1(n7630), .DIN2(n7591), .Q(n7626) );
  xor2s1 U8007 ( .DIN1(n5078), .DIN2(w0[25]), .Q(n7630) );
  nnd2s1 U8008 ( .DIN1(n7631), .DIN2(n1604), .Q(n7623) );
  xor2s1 U8009 ( .DIN1(w0[25]), .DIN2(text_in_r[121]), .Q(n7631) );
  nnd2s1 U8010 ( .DIN1(n7632), .DIN2(n7633), .Q(N274) );
  nnd2s1 U8011 ( .DIN1(n7634), .DIN2(n1618), .Q(n7633) );
  xor2s1 U8012 ( .DIN1(n7635), .DIN2(n7636), .Q(n7634) );
  xor2s1 U8013 ( .DIN1(n7591), .DIN2(n7637), .Q(n7636) );
  xor2s1 U8014 ( .DIN1(n1481), .DIN2(n5077), .Q(n7635) );
  nnd2s1 U8015 ( .DIN1(n7638), .DIN2(n1604), .Q(n7632) );
  xor2s1 U8016 ( .DIN1(w0[24]), .DIN2(text_in_r[120]), .Q(n7638) );
  nnd2s1 U8017 ( .DIN1(n7639), .DIN2(n7640), .Q(N265) );
  nnd2s1 U8018 ( .DIN1(n7641), .DIN2(n1618), .Q(n7640) );
  xor2s1 U8019 ( .DIN1(n7642), .DIN2(n7643), .Q(n7641) );
  xor2s1 U8020 ( .DIN1(n6115), .DIN2(n7644), .Q(n7643) );
  xor2s1 U8021 ( .DIN1(n5083), .DIN2(n7645), .Q(n7642) );
  xor2s1 U8022 ( .DIN1(n1463), .DIN2(n5059), .Q(n7645) );
  nnd2s1 U8023 ( .DIN1(n7646), .DIN2(n1604), .Q(n7639) );
  xor2s1 U8024 ( .DIN1(w0[23]), .DIN2(text_in_r[119]), .Q(n7646) );
  nnd3s1 U8025 ( .DIN1(n7647), .DIN2(n7648), .DIN3(n7649), .Q(N264) );
  nnd2s1 U8026 ( .DIN1(n1598), .DIN2(n7650), .Q(n7649) );
  xor2s1 U8027 ( .DIN1(w0[22]), .DIN2(text_in_r[118]), .Q(n7650) );
  nnd2s1 U8028 ( .DIN1(n7651), .DIN2(n7652), .Q(n7648) );
  nnd2s1 U8029 ( .DIN1(n7653), .DIN2(n7654), .Q(n7651) );
  nnd2s1 U8030 ( .DIN1(n7655), .DIN2(n7656), .Q(n7654) );
  nnd2s1 U8031 ( .DIN1(n7657), .DIN2(n7658), .Q(n7653) );
  nnd2s1 U8032 ( .DIN1(n7568), .DIN2(n7659), .Q(n7647) );
  nnd2s1 U8033 ( .DIN1(n7660), .DIN2(n7661), .Q(n7659) );
  nnd2s1 U8034 ( .DIN1(n7657), .DIN2(n7656), .Q(n7661) );
  nnd2s1 U8035 ( .DIN1(n7658), .DIN2(n7655), .Q(n7660) );
  hi1s1 U8036 ( .DIN(n7656), .Q(n7658) );
  xnr2s1 U8037 ( .DIN1(n5082), .DIN2(n7662), .Q(n7656) );
  xor2s1 U8038 ( .DIN1(w0[22]), .DIN2(n5058), .Q(n7662) );
  nnd3s1 U8039 ( .DIN1(n7663), .DIN2(n7664), .DIN3(n7665), .Q(N263) );
  nnd2s1 U8040 ( .DIN1(n1598), .DIN2(n7666), .Q(n7665) );
  xor2s1 U8041 ( .DIN1(w0[21]), .DIN2(text_in_r[117]), .Q(n7666) );
  nnd2s1 U8042 ( .DIN1(n7667), .DIN2(n7668), .Q(n7664) );
  nnd2s1 U8043 ( .DIN1(n7669), .DIN2(n7670), .Q(n7667) );
  nnd2s1 U8044 ( .DIN1(n7671), .DIN2(n7672), .Q(n7670) );
  nnd2s1 U8045 ( .DIN1(n7673), .DIN2(n7674), .Q(n7669) );
  nnd2s1 U8046 ( .DIN1(n7576), .DIN2(n7675), .Q(n7663) );
  nnd2s1 U8047 ( .DIN1(n7676), .DIN2(n7677), .Q(n7675) );
  nnd2s1 U8048 ( .DIN1(n7673), .DIN2(n7672), .Q(n7677) );
  nnd2s1 U8049 ( .DIN1(n7674), .DIN2(n7671), .Q(n7676) );
  hi1s1 U8050 ( .DIN(n7672), .Q(n7674) );
  xor2s1 U8051 ( .DIN1(n7678), .DIN2(n7679), .Q(n7672) );
  xor2s1 U8052 ( .DIN1(w0[21]), .DIN2(n5057), .Q(n7679) );
  nnd2s1 U8053 ( .DIN1(n7680), .DIN2(n7681), .Q(N262) );
  nnd2s1 U8054 ( .DIN1(n7682), .DIN2(n1618), .Q(n7681) );
  xor2s1 U8055 ( .DIN1(n7683), .DIN2(n7684), .Q(n7682) );
  xor2s1 U8056 ( .DIN1(n7685), .DIN2(n7686), .Q(n7684) );
  xnr2s1 U8057 ( .DIN1(n5706), .DIN2(n7596), .Q(n7686) );
  xor2s1 U8058 ( .DIN1(n5080), .DIN2(n7687), .Q(n7683) );
  xor2s1 U8059 ( .DIN1(n1464), .DIN2(n5056), .Q(n7687) );
  nnd2s1 U8060 ( .DIN1(n7688), .DIN2(n1604), .Q(n7680) );
  xor2s1 U8061 ( .DIN1(w0[20]), .DIN2(text_in_r[116]), .Q(n7688) );
  nnd2s1 U8062 ( .DIN1(n7689), .DIN2(n7690), .Q(N261) );
  nnd2s1 U8063 ( .DIN1(n7691), .DIN2(n1619), .Q(n7690) );
  xor2s1 U8064 ( .DIN1(n7692), .DIN2(n7693), .Q(n7691) );
  xor2s1 U8065 ( .DIN1(n7685), .DIN2(n7694), .Q(n7693) );
  xor2s1 U8066 ( .DIN1(n5705), .DIN2(n7602), .Q(n7694) );
  xor2s1 U8067 ( .DIN1(n7621), .DIN2(n7695), .Q(n7692) );
  xor2s1 U8068 ( .DIN1(n1500), .DIN2(n5055), .Q(n7695) );
  nnd2s1 U8069 ( .DIN1(n7696), .DIN2(n1604), .Q(n7689) );
  xor2s1 U8070 ( .DIN1(w0[19]), .DIN2(text_in_r[115]), .Q(n7696) );
  nnd2s1 U8071 ( .DIN1(n7697), .DIN2(n7698), .Q(N260) );
  nnd2s1 U8072 ( .DIN1(n7699), .DIN2(n1619), .Q(n7698) );
  xor2s1 U8073 ( .DIN1(n7700), .DIN2(n7701), .Q(n7699) );
  xor2s1 U8074 ( .DIN1(n5704), .DIN2(n7702), .Q(n7701) );
  xor2s1 U8075 ( .DIN1(n5078), .DIN2(n7703), .Q(n7700) );
  xor2s1 U8076 ( .DIN1(n1465), .DIN2(n5054), .Q(n7703) );
  nnd2s1 U8077 ( .DIN1(n7704), .DIN2(n1604), .Q(n7697) );
  xor2s1 U8078 ( .DIN1(w0[18]), .DIN2(text_in_r[114]), .Q(n7704) );
  nnd2s1 U8079 ( .DIN1(n7705), .DIN2(n7706), .Q(N259) );
  nnd2s1 U8080 ( .DIN1(n7707), .DIN2(n1619), .Q(n7706) );
  xor2s1 U8081 ( .DIN1(n7708), .DIN2(n7709), .Q(n7707) );
  xor2s1 U8082 ( .DIN1(n7685), .DIN2(n7710), .Q(n7709) );
  xor2s1 U8083 ( .DIN1(n5703), .DIN2(n7629), .Q(n7710) );
  xnr2s1 U8084 ( .DIN1(n5077), .DIN2(n7711), .Q(n7708) );
  xor2s1 U8085 ( .DIN1(n1501), .DIN2(n7712), .Q(n7711) );
  nnd2s1 U8086 ( .DIN1(n7713), .DIN2(n1604), .Q(n7705) );
  xor2s1 U8087 ( .DIN1(w0[17]), .DIN2(text_in_r[113]), .Q(n7713) );
  nnd2s1 U8088 ( .DIN1(n7714), .DIN2(n7715), .Q(N258) );
  nnd2s1 U8089 ( .DIN1(n7716), .DIN2(n1620), .Q(n7715) );
  xor2s1 U8090 ( .DIN1(n7717), .DIN2(n7718), .Q(n7716) );
  xor2s1 U8091 ( .DIN1(n7637), .DIN2(n7685), .Q(n7718) );
  xor2s1 U8092 ( .DIN1(n5084), .DIN2(n5060), .Q(n7685) );
  xor2s1 U8093 ( .DIN1(n1466), .DIN2(n5702), .Q(n7717) );
  nnd2s1 U8094 ( .DIN1(n7719), .DIN2(n1604), .Q(n7714) );
  xor2s1 U8095 ( .DIN1(w0[16]), .DIN2(text_in_r[112]), .Q(n7719) );
  nnd2s1 U8096 ( .DIN1(n7720), .DIN2(n7721), .Q(N249) );
  nnd2s1 U8097 ( .DIN1(n7722), .DIN2(n1620), .Q(n7721) );
  xor2s1 U8098 ( .DIN1(n7723), .DIN2(n7724), .Q(n7722) );
  xor2s1 U8099 ( .DIN1(n7568), .DIN2(n7591), .Q(n7724) );
  hi1s1 U8100 ( .DIN(n7652), .Q(n7568) );
  xor2s1 U8101 ( .DIN1(n5036), .DIN2(n7725), .Q(n7652) );
  hi1s1 U8102 ( .DIN(n5059), .Q(n7725) );
  xor2s1 U8103 ( .DIN1(n1467), .DIN2(n5037), .Q(n7723) );
  nnd2s1 U8104 ( .DIN1(n7726), .DIN2(n1604), .Q(n7720) );
  xor2s1 U8105 ( .DIN1(w0[15]), .DIN2(text_in_r[111]), .Q(n7726) );
  nnd2s1 U8106 ( .DIN1(n7727), .DIN2(n7728), .Q(N248) );
  nnd2s1 U8107 ( .DIN1(n7729), .DIN2(n1620), .Q(n7728) );
  xor2s1 U8108 ( .DIN1(n7730), .DIN2(n7731), .Q(n7729) );
  xor2s1 U8109 ( .DIN1(n1502), .DIN2(n5036), .Q(n7731) );
  xor2s1 U8110 ( .DIN1(n7668), .DIN2(n7560), .Q(n7730) );
  hi1s1 U8111 ( .DIN(n7576), .Q(n7668) );
  xnr2s1 U8112 ( .DIN1(n7732), .DIN2(n5058), .Q(n7576) );
  hi1s1 U8113 ( .DIN(n7733), .Q(n5058) );
  nnd2s1 U8114 ( .DIN1(n7734), .DIN2(n1604), .Q(n7727) );
  xor2s1 U8115 ( .DIN1(w0[14]), .DIN2(text_in_r[110]), .Q(n7734) );
  nnd2s1 U8116 ( .DIN1(n7735), .DIN2(n7736), .Q(N247) );
  nnd2s1 U8117 ( .DIN1(n7737), .DIN2(n1621), .Q(n7736) );
  xor2s1 U8118 ( .DIN1(n7738), .DIN2(n7739), .Q(n7737) );
  xor2s1 U8119 ( .DIN1(n7569), .DIN2(n7596), .Q(n7739) );
  xnr2s1 U8120 ( .DIN1(n7740), .DIN2(n5057), .Q(n7596) );
  hi1s1 U8121 ( .DIN(n7741), .Q(n5057) );
  xor2s1 U8122 ( .DIN1(n1468), .DIN2(n5035), .Q(n7738) );
  hi1s1 U8123 ( .DIN(n7732), .Q(n5035) );
  nnd2s1 U8124 ( .DIN1(n7742), .DIN2(n1604), .Q(n7735) );
  xor2s1 U8125 ( .DIN1(w0[13]), .DIN2(text_in_r[109]), .Q(n7742) );
  nnd2s1 U8126 ( .DIN1(n7743), .DIN2(n7744), .Q(N246) );
  nnd2s1 U8127 ( .DIN1(n7745), .DIN2(n1621), .Q(n7744) );
  xor2s1 U8128 ( .DIN1(n7746), .DIN2(n7747), .Q(n7745) );
  xor2s1 U8129 ( .DIN1(n7577), .DIN2(n7609), .Q(n7747) );
  hi1s1 U8130 ( .DIN(n7602), .Q(n7609) );
  xor2s1 U8131 ( .DIN1(n5033), .DIN2(n7748), .Q(n7602) );
  hi1s1 U8132 ( .DIN(n5056), .Q(n7748) );
  xor2s1 U8133 ( .DIN1(n7749), .DIN2(n7559), .Q(n7746) );
  xor2s1 U8134 ( .DIN1(n1469), .DIN2(n5034), .Q(n7749) );
  hi1s1 U8135 ( .DIN(n7740), .Q(n5034) );
  nnd2s1 U8136 ( .DIN1(n7750), .DIN2(n1603), .Q(n7743) );
  xor2s1 U8137 ( .DIN1(w0[12]), .DIN2(text_in_r[108]), .Q(n7750) );
  nnd3s1 U8138 ( .DIN1(n7751), .DIN2(n7752), .DIN3(n7753), .Q(N245) );
  nnd2s1 U8139 ( .DIN1(n1598), .DIN2(n7754), .Q(n7753) );
  xor2s1 U8140 ( .DIN1(w0[11]), .DIN2(text_in_r[107]), .Q(n7754) );
  nnd2s1 U8141 ( .DIN1(n7755), .DIN2(n7756), .Q(n7752) );
  nnd2s1 U8142 ( .DIN1(n7757), .DIN2(n7758), .Q(n7755) );
  nnd2s1 U8143 ( .DIN1(n7587), .DIN2(n7702), .Q(n7758) );
  nnd2s1 U8144 ( .DIN1(n7619), .DIN2(n7589), .Q(n7757) );
  nnd2s1 U8145 ( .DIN1(n7759), .DIN2(n7760), .Q(n7751) );
  nnd2s1 U8146 ( .DIN1(n7761), .DIN2(n7762), .Q(n7760) );
  nnd2s1 U8147 ( .DIN1(n7589), .DIN2(n7702), .Q(n7762) );
  and2s1 U8148 ( .DIN1(n7763), .DIN2(n1640), .Q(n7589) );
  nnd2s1 U8149 ( .DIN1(n7619), .DIN2(n7587), .Q(n7761) );
  nor2s1 U8150 ( .DIN1(n7763), .DIN2(n1595), .Q(n7587) );
  hi1s1 U8151 ( .DIN(n7702), .Q(n7619) );
  xor2s1 U8152 ( .DIN1(n5055), .DIN2(n7764), .Q(n7702) );
  hi1s1 U8153 ( .DIN(n7756), .Q(n7759) );
  xor2s1 U8154 ( .DIN1(n7765), .DIN2(n7559), .Q(n7756) );
  xor2s1 U8155 ( .DIN1(n5033), .DIN2(w0[11]), .Q(n7765) );
  nnd2s1 U8156 ( .DIN1(n7766), .DIN2(n7767), .Q(N244) );
  nnd2s1 U8157 ( .DIN1(n7768), .DIN2(n1621), .Q(n7767) );
  xor2s1 U8158 ( .DIN1(n7769), .DIN2(n7770), .Q(n7768) );
  xor2s1 U8159 ( .DIN1(n7771), .DIN2(n7629), .Q(n7770) );
  xnr2s1 U8160 ( .DIN1(n5054), .DIN2(n5031), .Q(n7629) );
  xor2s1 U8161 ( .DIN1(n1499), .DIN2(n7764), .Q(n7769) );
  hi1s1 U8162 ( .DIN(n5032), .Q(n7764) );
  nnd2s1 U8163 ( .DIN1(n7772), .DIN2(n1603), .Q(n7766) );
  xor2s1 U8164 ( .DIN1(w0[10]), .DIN2(text_in_r[106]), .Q(n7772) );
  nnd2s1 U8165 ( .DIN1(n7773), .DIN2(n7774), .Q(N243) );
  nnd2s1 U8166 ( .DIN1(n7775), .DIN2(n1622), .Q(n7774) );
  xor2s1 U8167 ( .DIN1(n7776), .DIN2(n7777), .Q(n7775) );
  xor2s1 U8168 ( .DIN1(n7559), .DIN2(n7778), .Q(n7777) );
  xor2s1 U8169 ( .DIN1(n1503), .DIN2(n5031), .Q(n7778) );
  xnr2s1 U8170 ( .DIN1(n7637), .DIN2(n7620), .Q(n7776) );
  xor2s1 U8171 ( .DIN1(n5053), .DIN2(n5030), .Q(n7637) );
  nnd2s1 U8172 ( .DIN1(n7779), .DIN2(n1603), .Q(n7773) );
  xor2s1 U8173 ( .DIN1(w0[9]), .DIN2(text_in_r[105]), .Q(n7779) );
  nnd2s1 U8174 ( .DIN1(n7780), .DIN2(n7781), .Q(N242) );
  nnd2s1 U8175 ( .DIN1(n7782), .DIN2(n1622), .Q(n7781) );
  xor2s1 U8176 ( .DIN1(n7783), .DIN2(n7784), .Q(n7782) );
  xor2s1 U8177 ( .DIN1(n7559), .DIN2(n7628), .Q(n7784) );
  hi1s1 U8178 ( .DIN(n7644), .Q(n7559) );
  xnr2s1 U8179 ( .DIN1(n5060), .DIN2(n5037), .Q(n7644) );
  xor2s1 U8180 ( .DIN1(n1470), .DIN2(n5030), .Q(n7783) );
  nnd2s1 U8181 ( .DIN1(n7785), .DIN2(n1603), .Q(n7780) );
  xor2s1 U8182 ( .DIN1(w0[8]), .DIN2(text_in_r[104]), .Q(n7785) );
  nnd3s1 U8183 ( .DIN1(n7786), .DIN2(n7787), .DIN3(n7788), .Q(N233) );
  nnd2s1 U8184 ( .DIN1(n1599), .DIN2(n7789), .Q(n7788) );
  xor2s1 U8185 ( .DIN1(w0[7]), .DIN2(text_in_r[103]), .Q(n7789) );
  nnd2s1 U8186 ( .DIN1(n7790), .DIN2(n7791), .Q(n7787) );
  nnd2s1 U8187 ( .DIN1(n7792), .DIN2(n7793), .Q(n7790) );
  nnd2s1 U8188 ( .DIN1(n7655), .DIN2(n7584), .Q(n7793) );
  nnd2s1 U8189 ( .DIN1(n7657), .DIN2(n7591), .Q(n7792) );
  nnd2s1 U8190 ( .DIN1(n7794), .DIN2(n7795), .Q(n7786) );
  nnd2s1 U8191 ( .DIN1(n7796), .DIN2(n7797), .Q(n7795) );
  nnd2s1 U8192 ( .DIN1(n7657), .DIN2(n7584), .Q(n7797) );
  nor2s1 U8193 ( .DIN1(n6114), .DIN2(n1596), .Q(n7657) );
  nnd2s1 U8194 ( .DIN1(n7655), .DIN2(n7591), .Q(n7796) );
  hi1s1 U8195 ( .DIN(n7584), .Q(n7591) );
  xor2s1 U8196 ( .DIN1(n6115), .DIN2(n5084), .Q(n7584) );
  hi1s1 U8197 ( .DIN(n7561), .Q(n5084) );
  or3s1 U8198 ( .DIN1(n7798), .DIN2(n7799), .DIN3(n7800), .Q(n7561) );
  nnd4s1 U8199 ( .DIN1(n7801), .DIN2(n7802), .DIN3(n7803), .DIN4(n7804), 
        .Q(n7800) );
  and4s1 U8200 ( .DIN1(n7805), .DIN2(n7806), .DIN3(n7807), .DIN4(n7808), 
        .Q(n7804) );
  nnd2s1 U8201 ( .DIN1(n7809), .DIN2(n7810), .Q(n7807) );
  nnd2s1 U8202 ( .DIN1(n7811), .DIN2(n7812), .Q(n7806) );
  nnd4s1 U8203 ( .DIN1(n7813), .DIN2(n7814), .DIN3(n7815), .DIN4(n7816), 
        .Q(n7799) );
  nnd2s1 U8204 ( .DIN1(n7817), .DIN2(n7818), .Q(n7816) );
  nnd2s1 U8205 ( .DIN1(n7819), .DIN2(n7820), .Q(n7815) );
  nnd2s1 U8206 ( .DIN1(n7821), .DIN2(n7822), .Q(n7814) );
  nnd4s1 U8207 ( .DIN1(n7823), .DIN2(n7824), .DIN3(n7825), .DIN4(n7826), 
        .Q(n7798) );
  nnd2s1 U8208 ( .DIN1(n7827), .DIN2(n7828), .Q(n7826) );
  nnd2s1 U8209 ( .DIN1(n7829), .DIN2(n7830), .Q(n7828) );
  nnd2s1 U8210 ( .DIN1(n7831), .DIN2(n7832), .Q(n7825) );
  nnd2s1 U8211 ( .DIN1(n7833), .DIN2(n7834), .Q(n7832) );
  nnd2s1 U8212 ( .DIN1(n7835), .DIN2(n7836), .Q(n7824) );
  nnd2s1 U8213 ( .DIN1(n7837), .DIN2(n7838), .Q(n7836) );
  nnd2s1 U8214 ( .DIN1(n7839), .DIN2(n7840), .Q(n7823) );
  and2s1 U8215 ( .DIN1(n6114), .DIN2(n1639), .Q(n7655) );
  hi1s1 U8216 ( .DIN(n7791), .Q(n7794) );
  xnr2s1 U8217 ( .DIN1(n5060), .DIN2(n7841), .Q(n7791) );
  xnr2s1 U8218 ( .DIN1(w0[7]), .DIN2(n5036), .Q(n7841) );
  or3s1 U8219 ( .DIN1(n7842), .DIN2(n7843), .DIN3(n7844), .Q(n5036) );
  nnd4s1 U8220 ( .DIN1(n7845), .DIN2(n7846), .DIN3(n7847), .DIN4(n7848), 
        .Q(n7844) );
  and3s1 U8221 ( .DIN1(n7849), .DIN2(n7850), .DIN3(n7851), .Q(n7848) );
  nnd2s1 U8222 ( .DIN1(n7852), .DIN2(n7853), .Q(n7845) );
  nnd3s1 U8223 ( .DIN1(n7854), .DIN2(n7855), .DIN3(n7856), .Q(n7843) );
  or2s1 U8224 ( .DIN1(n7857), .DIN2(n7858), .Q(n7856) );
  or2s1 U8225 ( .DIN1(n7859), .DIN2(n7860), .Q(n7855) );
  nnd2s1 U8226 ( .DIN1(n7861), .DIN2(n7862), .Q(n7854) );
  nnd3s1 U8227 ( .DIN1(n7863), .DIN2(n7864), .DIN3(n7865), .Q(n7842) );
  nnd2s1 U8228 ( .DIN1(n7866), .DIN2(n7867), .Q(n7865) );
  nnd2s1 U8229 ( .DIN1(n7868), .DIN2(n7869), .Q(n7867) );
  nnd2s1 U8230 ( .DIN1(n7870), .DIN2(n7871), .Q(n7864) );
  nnd2s1 U8231 ( .DIN1(n7872), .DIN2(n7873), .Q(n7871) );
  hi1s1 U8232 ( .DIN(n7874), .Q(n7873) );
  nnd2s1 U8233 ( .DIN1(n7875), .DIN2(n7876), .Q(n7863) );
  nnd2s1 U8234 ( .DIN1(n7877), .DIN2(n7878), .Q(n7876) );
  nor3s1 U8235 ( .DIN1(n7879), .DIN2(n7880), .DIN3(n7881), .Q(n5060) );
  nnd4s1 U8236 ( .DIN1(n7882), .DIN2(n7883), .DIN3(n7884), .DIN4(n7885), 
        .Q(n7881) );
  and4s1 U8237 ( .DIN1(n7886), .DIN2(n7887), .DIN3(n7888), .DIN4(n7889), 
        .Q(n7885) );
  nnd2s1 U8238 ( .DIN1(n7890), .DIN2(n7891), .Q(n7888) );
  nnd2s1 U8239 ( .DIN1(n7892), .DIN2(n7893), .Q(n7887) );
  nnd4s1 U8240 ( .DIN1(n7894), .DIN2(n7895), .DIN3(n7896), .DIN4(n7897), 
        .Q(n7880) );
  nnd2s1 U8241 ( .DIN1(n7898), .DIN2(n7899), .Q(n7897) );
  nnd2s1 U8242 ( .DIN1(n7900), .DIN2(n7901), .Q(n7896) );
  nnd2s1 U8243 ( .DIN1(n7902), .DIN2(n7903), .Q(n7895) );
  nnd4s1 U8244 ( .DIN1(n7904), .DIN2(n7905), .DIN3(n7906), .DIN4(n7907), 
        .Q(n7879) );
  nnd2s1 U8245 ( .DIN1(n7908), .DIN2(n7909), .Q(n7907) );
  nnd2s1 U8246 ( .DIN1(n7910), .DIN2(n7911), .Q(n7909) );
  nnd2s1 U8247 ( .DIN1(n7912), .DIN2(n7913), .Q(n7906) );
  nnd2s1 U8248 ( .DIN1(n7914), .DIN2(n7915), .Q(n7913) );
  nnd2s1 U8249 ( .DIN1(n7916), .DIN2(n7917), .Q(n7905) );
  nnd2s1 U8250 ( .DIN1(n7918), .DIN2(n7919), .Q(n7917) );
  nnd2s1 U8251 ( .DIN1(n7920), .DIN2(n7921), .Q(n7904) );
  nnd3s1 U8252 ( .DIN1(n7922), .DIN2(n7923), .DIN3(n7924), .Q(N232) );
  nnd2s1 U8253 ( .DIN1(n1599), .DIN2(n7925), .Q(n7924) );
  xor2s1 U8254 ( .DIN1(w0[6]), .DIN2(text_in_r[102]), .Q(n7925) );
  nnd2s1 U8255 ( .DIN1(n7926), .DIN2(n7927), .Q(n7923) );
  nnd2s1 U8256 ( .DIN1(n7928), .DIN2(n7929), .Q(n7926) );
  nnd2s1 U8257 ( .DIN1(n7671), .DIN2(n7930), .Q(n7929) );
  nnd2s1 U8258 ( .DIN1(n7560), .DIN2(n7673), .Q(n7928) );
  nnd2s1 U8259 ( .DIN1(n7931), .DIN2(n7932), .Q(n7922) );
  nnd2s1 U8260 ( .DIN1(n7933), .DIN2(n7934), .Q(n7932) );
  nnd2s1 U8261 ( .DIN1(n7673), .DIN2(n7930), .Q(n7934) );
  nor2s1 U8262 ( .DIN1(n7935), .DIN2(n1596), .Q(n7673) );
  nnd2s1 U8263 ( .DIN1(n7560), .DIN2(n7671), .Q(n7933) );
  nor2s1 U8264 ( .DIN1(n5707), .DIN2(n1596), .Q(n7671) );
  hi1s1 U8265 ( .DIN(n7935), .Q(n5707) );
  hi1s1 U8266 ( .DIN(n7930), .Q(n7560) );
  xor2s1 U8267 ( .DIN1(n6114), .DIN2(n7936), .Q(n7930) );
  hi1s1 U8268 ( .DIN(n5083), .Q(n7936) );
  or3s1 U8269 ( .DIN1(n7937), .DIN2(n7938), .DIN3(n7939), .Q(n5083) );
  nnd4s1 U8270 ( .DIN1(n7940), .DIN2(n7941), .DIN3(n7942), .DIN4(n7943), 
        .Q(n7939) );
  and3s1 U8271 ( .DIN1(n7944), .DIN2(n7945), .DIN3(n7946), .Q(n7943) );
  nnd2s1 U8272 ( .DIN1(n7947), .DIN2(n7819), .Q(n7941) );
  nnd2s1 U8273 ( .DIN1(n7810), .DIN2(n7948), .Q(n7940) );
  nnd3s1 U8274 ( .DIN1(n7949), .DIN2(n7950), .DIN3(n7951), .Q(n7938) );
  or2s1 U8275 ( .DIN1(n7952), .DIN2(n7953), .Q(n7951) );
  or2s1 U8276 ( .DIN1(n7834), .DIN2(n7954), .Q(n7950) );
  nnd2s1 U8277 ( .DIN1(n7835), .DIN2(n7955), .Q(n7949) );
  nnd3s1 U8278 ( .DIN1(n7956), .DIN2(n7957), .DIN3(n7958), .Q(n7937) );
  nnd2s1 U8279 ( .DIN1(n7959), .DIN2(n7960), .Q(n7958) );
  nnd2s1 U8280 ( .DIN1(n7961), .DIN2(n7962), .Q(n7960) );
  nnd2s1 U8281 ( .DIN1(n7963), .DIN2(n7964), .Q(n7957) );
  nnd2s1 U8282 ( .DIN1(n7965), .DIN2(n7966), .Q(n7964) );
  nnd2s1 U8283 ( .DIN1(n7811), .DIN2(n7967), .Q(n7956) );
  nnd2s1 U8284 ( .DIN1(n7968), .DIN2(n7969), .Q(n7967) );
  hi1s1 U8285 ( .DIN(n7970), .Q(n7969) );
  or3s1 U8286 ( .DIN1(n7971), .DIN2(n7972), .DIN3(n7973), .Q(n6114) );
  nnd4s1 U8287 ( .DIN1(n7974), .DIN2(n7975), .DIN3(n7976), .DIN4(n7977), 
        .Q(n7973) );
  and3s1 U8288 ( .DIN1(n7978), .DIN2(n7979), .DIN3(n7980), .Q(n7977) );
  nnd2s1 U8289 ( .DIN1(n7981), .DIN2(n7982), .Q(n7975) );
  nnd2s1 U8290 ( .DIN1(n7983), .DIN2(n7984), .Q(n7974) );
  nnd3s1 U8291 ( .DIN1(n7985), .DIN2(n7986), .DIN3(n7987), .Q(n7972) );
  or2s1 U8292 ( .DIN1(n7988), .DIN2(n7989), .Q(n7987) );
  or2s1 U8293 ( .DIN1(n7990), .DIN2(n7991), .Q(n7986) );
  nnd2s1 U8294 ( .DIN1(n7992), .DIN2(n7993), .Q(n7985) );
  nnd3s1 U8295 ( .DIN1(n7994), .DIN2(n7995), .DIN3(n7996), .Q(n7971) );
  nnd2s1 U8296 ( .DIN1(n7997), .DIN2(n7998), .Q(n7996) );
  nnd2s1 U8297 ( .DIN1(n7999), .DIN2(n8000), .Q(n7998) );
  nnd2s1 U8298 ( .DIN1(n8001), .DIN2(n8002), .Q(n7995) );
  nnd2s1 U8299 ( .DIN1(n8003), .DIN2(n8004), .Q(n8002) );
  nnd2s1 U8300 ( .DIN1(n8005), .DIN2(n8006), .Q(n7994) );
  nnd2s1 U8301 ( .DIN1(n8007), .DIN2(n8008), .Q(n8006) );
  hi1s1 U8302 ( .DIN(n8009), .Q(n8008) );
  hi1s1 U8303 ( .DIN(n7927), .Q(n7931) );
  xor2s1 U8304 ( .DIN1(n5059), .DIN2(n8010), .Q(n7927) );
  xor2s1 U8305 ( .DIN1(n1504), .DIN2(n7732), .Q(n8010) );
  or3s1 U8306 ( .DIN1(n8011), .DIN2(n8012), .DIN3(n8013), .Q(n7732) );
  nnd4s1 U8307 ( .DIN1(n8014), .DIN2(n8015), .DIN3(n7851), .DIN4(n8016), 
        .Q(n8013) );
  and4s1 U8308 ( .DIN1(n8017), .DIN2(n8018), .DIN3(n8019), .DIN4(n8020), 
        .Q(n8016) );
  nnd2s1 U8309 ( .DIN1(n7852), .DIN2(n8021), .Q(n8020) );
  nnd2s1 U8310 ( .DIN1(n7866), .DIN2(n8022), .Q(n8019) );
  nnd2s1 U8311 ( .DIN1(n8023), .DIN2(n7875), .Q(n8018) );
  nor2s1 U8312 ( .DIN1(n8024), .DIN2(n8025), .Q(n7851) );
  nnd4s1 U8313 ( .DIN1(n8026), .DIN2(n8027), .DIN3(n8028), .DIN4(n8029), 
        .Q(n8025) );
  nnd2s1 U8314 ( .DIN1(n8030), .DIN2(n8031), .Q(n8029) );
  nnd3s1 U8315 ( .DIN1(n8032), .DIN2(n7878), .DIN3(n8033), .Q(n8031) );
  nnd2s1 U8316 ( .DIN1(n8034), .DIN2(n8035), .Q(n8028) );
  nnd2s1 U8317 ( .DIN1(n8023), .DIN2(n8036), .Q(n8027) );
  nnd2s1 U8318 ( .DIN1(n8037), .DIN2(n8021), .Q(n8026) );
  nnd4s1 U8319 ( .DIN1(n8038), .DIN2(n8039), .DIN3(n8040), .DIN4(n8041), 
        .Q(n8024) );
  nnd2s1 U8320 ( .DIN1(n8042), .DIN2(n8043), .Q(n8041) );
  nnd2s1 U8321 ( .DIN1(n8044), .DIN2(n8045), .Q(n8043) );
  nnd2s1 U8322 ( .DIN1(n8022), .DIN2(n8046), .Q(n8040) );
  nnd2s1 U8323 ( .DIN1(n8047), .DIN2(n8048), .Q(n8046) );
  nnd2s1 U8324 ( .DIN1(n8049), .DIN2(n8050), .Q(n8039) );
  nnd2s1 U8325 ( .DIN1(n8051), .DIN2(n7869), .Q(n8050) );
  nnd2s1 U8326 ( .DIN1(n8052), .DIN2(n8053), .Q(n8038) );
  nnd2s1 U8327 ( .DIN1(n7878), .DIN2(n8054), .Q(n8053) );
  nnd4s1 U8328 ( .DIN1(n8055), .DIN2(n8056), .DIN3(n8057), .DIN4(n8058), 
        .Q(n8012) );
  or2s1 U8329 ( .DIN1(n8059), .DIN2(n8060), .Q(n8058) );
  nnd2s1 U8330 ( .DIN1(n8037), .DIN2(n8061), .Q(n8057) );
  nnd2s1 U8331 ( .DIN1(n8062), .DIN2(n8063), .Q(n8056) );
  nnd2s1 U8332 ( .DIN1(n8034), .DIN2(n8064), .Q(n8055) );
  nnd4s1 U8333 ( .DIN1(n8065), .DIN2(n8066), .DIN3(n8067), .DIN4(n8068), 
        .Q(n8011) );
  nnd2s1 U8334 ( .DIN1(n8069), .DIN2(n8070), .Q(n8068) );
  nnd2s1 U8335 ( .DIN1(n8032), .DIN2(n8071), .Q(n8070) );
  nnd2s1 U8336 ( .DIN1(n8072), .DIN2(n8073), .Q(n8067) );
  nnd2s1 U8337 ( .DIN1(n7868), .DIN2(n8074), .Q(n8073) );
  nnd2s1 U8338 ( .DIN1(n7861), .DIN2(n8075), .Q(n8066) );
  nnd2s1 U8339 ( .DIN1(n8076), .DIN2(n8077), .Q(n8075) );
  nnd2s1 U8340 ( .DIN1(n8078), .DIN2(n8079), .Q(n8065) );
  or3s1 U8341 ( .DIN1(n8080), .DIN2(n8081), .DIN3(n8082), .Q(n5059) );
  nnd4s1 U8342 ( .DIN1(n8083), .DIN2(n8084), .DIN3(n8085), .DIN4(n8086), 
        .Q(n8082) );
  and3s1 U8343 ( .DIN1(n8087), .DIN2(n8088), .DIN3(n8089), .Q(n8086) );
  nnd2s1 U8344 ( .DIN1(n8090), .DIN2(n7900), .Q(n8084) );
  nnd2s1 U8345 ( .DIN1(n7891), .DIN2(n8091), .Q(n8083) );
  nnd3s1 U8346 ( .DIN1(n8092), .DIN2(n8093), .DIN3(n8094), .Q(n8081) );
  or2s1 U8347 ( .DIN1(n8095), .DIN2(n8096), .Q(n8094) );
  or2s1 U8348 ( .DIN1(n7915), .DIN2(n8097), .Q(n8093) );
  nnd2s1 U8349 ( .DIN1(n7916), .DIN2(n8098), .Q(n8092) );
  nnd3s1 U8350 ( .DIN1(n8099), .DIN2(n8100), .DIN3(n8101), .Q(n8080) );
  nnd2s1 U8351 ( .DIN1(n8102), .DIN2(n8103), .Q(n8101) );
  nnd2s1 U8352 ( .DIN1(n8104), .DIN2(n8105), .Q(n8103) );
  nnd2s1 U8353 ( .DIN1(n8106), .DIN2(n8107), .Q(n8100) );
  nnd2s1 U8354 ( .DIN1(n8108), .DIN2(n8109), .Q(n8107) );
  nnd2s1 U8355 ( .DIN1(n7892), .DIN2(n8110), .Q(n8099) );
  nnd2s1 U8356 ( .DIN1(n8111), .DIN2(n8112), .Q(n8110) );
  hi1s1 U8357 ( .DIN(n8113), .Q(n8112) );
  nnd2s1 U8358 ( .DIN1(n8114), .DIN2(n8115), .Q(N231) );
  nnd2s1 U8359 ( .DIN1(n8116), .DIN2(n1622), .Q(n8115) );
  xor2s1 U8360 ( .DIN1(n8117), .DIN2(n8118), .Q(n8116) );
  xnr2s1 U8361 ( .DIN1(n5706), .DIN2(n7569), .Q(n8118) );
  xnr2s1 U8362 ( .DIN1(n7935), .DIN2(n5082), .Q(n7569) );
  nor3s1 U8363 ( .DIN1(n8119), .DIN2(n8120), .DIN3(n8121), .Q(n5082) );
  nnd4s1 U8364 ( .DIN1(n8122), .DIN2(n8123), .DIN3(n7946), .DIN4(n8124), 
        .Q(n8121) );
  and4s1 U8365 ( .DIN1(n8125), .DIN2(n8126), .DIN3(n8127), .DIN4(n7808), 
        .Q(n8124) );
  nnd2s1 U8366 ( .DIN1(n8128), .DIN2(n7963), .Q(n7808) );
  nnd2s1 U8367 ( .DIN1(n7959), .DIN2(n8129), .Q(n8127) );
  nnd2s1 U8368 ( .DIN1(n8130), .DIN2(n7812), .Q(n8126) );
  nor2s1 U8369 ( .DIN1(n8131), .DIN2(n8132), .Q(n7946) );
  nnd4s1 U8370 ( .DIN1(n8133), .DIN2(n8134), .DIN3(n8135), .DIN4(n8136), 
        .Q(n8132) );
  or2s1 U8371 ( .DIN1(n8137), .DIN2(n8138), .Q(n8136) );
  nnd2s1 U8372 ( .DIN1(n8130), .DIN2(n8139), .Q(n8135) );
  nnd2s1 U8373 ( .DIN1(n8128), .DIN2(n7810), .Q(n8134) );
  nnd2s1 U8374 ( .DIN1(n7822), .DIN2(n8140), .Q(n8133) );
  nnd4s1 U8375 ( .DIN1(n8141), .DIN2(n8142), .DIN3(n8143), .DIN4(n8144), 
        .Q(n8131) );
  nnd2s1 U8376 ( .DIN1(n7821), .DIN2(n8145), .Q(n8144) );
  nnd2s1 U8377 ( .DIN1(n7965), .DIN2(n8146), .Q(n8145) );
  nnd2s1 U8378 ( .DIN1(n8147), .DIN2(n8148), .Q(n8143) );
  nnd2s1 U8379 ( .DIN1(n7961), .DIN2(n8149), .Q(n8148) );
  nnd2s1 U8380 ( .DIN1(n8129), .DIN2(n8150), .Q(n8142) );
  nnd2s1 U8381 ( .DIN1(n8151), .DIN2(n8152), .Q(n8150) );
  nnd2s1 U8382 ( .DIN1(n7831), .DIN2(n8153), .Q(n8141) );
  nnd3s1 U8383 ( .DIN1(n8154), .DIN2(n7965), .DIN3(n8155), .Q(n8153) );
  nnd4s1 U8384 ( .DIN1(n8156), .DIN2(n8157), .DIN3(n8158), .DIN4(n8159), 
        .Q(n8120) );
  nnd2s1 U8385 ( .DIN1(n8160), .DIN2(n8161), .Q(n8159) );
  nnd2s1 U8386 ( .DIN1(n7822), .DIN2(n8162), .Q(n8158) );
  nnd2s1 U8387 ( .DIN1(n7809), .DIN2(n8163), .Q(n8157) );
  nnd2s1 U8388 ( .DIN1(n7947), .DIN2(n8140), .Q(n8156) );
  nnd4s1 U8389 ( .DIN1(n8164), .DIN2(n8165), .DIN3(n8166), .DIN4(n8167), 
        .Q(n8119) );
  nnd2s1 U8390 ( .DIN1(n7839), .DIN2(n8168), .Q(n8167) );
  nnd2s1 U8391 ( .DIN1(n7962), .DIN2(n8169), .Q(n8168) );
  nnd2s1 U8392 ( .DIN1(n8170), .DIN2(n8171), .Q(n8166) );
  nnd2s1 U8393 ( .DIN1(n7835), .DIN2(n8172), .Q(n8165) );
  nnd2s1 U8394 ( .DIN1(n8173), .DIN2(n7830), .Q(n8172) );
  nnd2s1 U8395 ( .DIN1(n7819), .DIN2(n8174), .Q(n8164) );
  or3s1 U8396 ( .DIN1(n8175), .DIN2(n8176), .DIN3(n8177), .Q(n7935) );
  nnd4s1 U8397 ( .DIN1(n8178), .DIN2(n8179), .DIN3(n7980), .DIN4(n8180), 
        .Q(n8177) );
  and4s1 U8398 ( .DIN1(n8181), .DIN2(n8182), .DIN3(n8183), .DIN4(n8184), 
        .Q(n8180) );
  nnd2s1 U8399 ( .DIN1(n7997), .DIN2(n8185), .Q(n8183) );
  nnd2s1 U8400 ( .DIN1(n8186), .DIN2(n8187), .Q(n8182) );
  nor2s1 U8401 ( .DIN1(n8188), .DIN2(n8189), .Q(n7980) );
  nnd4s1 U8402 ( .DIN1(n8190), .DIN2(n8191), .DIN3(n8192), .DIN4(n8193), 
        .Q(n8189) );
  or2s1 U8403 ( .DIN1(n8194), .DIN2(n8195), .Q(n8193) );
  nnd2s1 U8404 ( .DIN1(n8186), .DIN2(n8196), .Q(n8192) );
  nnd2s1 U8405 ( .DIN1(n8197), .DIN2(n7983), .Q(n8191) );
  nnd2s1 U8406 ( .DIN1(n8198), .DIN2(n8199), .Q(n8190) );
  nnd4s1 U8407 ( .DIN1(n8200), .DIN2(n8201), .DIN3(n8202), .DIN4(n8203), 
        .Q(n8188) );
  nnd2s1 U8408 ( .DIN1(n8204), .DIN2(n8205), .Q(n8203) );
  nnd2s1 U8409 ( .DIN1(n8003), .DIN2(n8206), .Q(n8205) );
  nnd2s1 U8410 ( .DIN1(n8207), .DIN2(n8208), .Q(n8202) );
  nnd2s1 U8411 ( .DIN1(n7999), .DIN2(n8209), .Q(n8208) );
  nnd2s1 U8412 ( .DIN1(n8185), .DIN2(n8210), .Q(n8201) );
  nnd2s1 U8413 ( .DIN1(n8211), .DIN2(n8212), .Q(n8210) );
  nnd2s1 U8414 ( .DIN1(n8213), .DIN2(n8214), .Q(n8200) );
  nnd3s1 U8415 ( .DIN1(n8215), .DIN2(n8003), .DIN3(n8216), .Q(n8214) );
  nnd4s1 U8416 ( .DIN1(n8217), .DIN2(n8218), .DIN3(n8219), .DIN4(n8220), 
        .Q(n8176) );
  nnd2s1 U8417 ( .DIN1(n8221), .DIN2(n8222), .Q(n8220) );
  nnd2s1 U8418 ( .DIN1(n8198), .DIN2(n8223), .Q(n8219) );
  nnd2s1 U8419 ( .DIN1(n8224), .DIN2(n8225), .Q(n8218) );
  nnd2s1 U8420 ( .DIN1(n7981), .DIN2(n8199), .Q(n8217) );
  nnd4s1 U8421 ( .DIN1(n8226), .DIN2(n8227), .DIN3(n8228), .DIN4(n8229), 
        .Q(n8175) );
  nnd2s1 U8422 ( .DIN1(n8230), .DIN2(n8231), .Q(n8229) );
  nnd2s1 U8423 ( .DIN1(n8000), .DIN2(n8232), .Q(n8231) );
  nnd2s1 U8424 ( .DIN1(n8233), .DIN2(n8234), .Q(n8228) );
  nnd2s1 U8425 ( .DIN1(n7992), .DIN2(n8235), .Q(n8227) );
  nnd2s1 U8426 ( .DIN1(n8236), .DIN2(n8237), .Q(n8235) );
  nnd2s1 U8427 ( .DIN1(n7982), .DIN2(n8238), .Q(n8226) );
  xor2s1 U8428 ( .DIN1(n7733), .DIN2(n8239), .Q(n8117) );
  xor2s1 U8429 ( .DIN1(n1471), .DIN2(n7740), .Q(n8239) );
  or3s1 U8430 ( .DIN1(n8240), .DIN2(n8241), .DIN3(n8242), .Q(n7740) );
  nnd4s1 U8431 ( .DIN1(n8243), .DIN2(n8244), .DIN3(n8245), .DIN4(n8246), 
        .Q(n8242) );
  and4s1 U8432 ( .DIN1(n8247), .DIN2(n8248), .DIN3(n8249), .DIN4(n8250), 
        .Q(n8246) );
  nnd2s1 U8433 ( .DIN1(n7852), .DIN2(n8251), .Q(n8250) );
  nnd2s1 U8434 ( .DIN1(n8252), .DIN2(n8253), .Q(n8251) );
  nnd2s1 U8435 ( .DIN1(n8254), .DIN2(n8255), .Q(n8249) );
  nnd2s1 U8436 ( .DIN1(n7868), .DIN2(n8054), .Q(n8255) );
  nnd2s1 U8437 ( .DIN1(n7875), .DIN2(n8256), .Q(n8248) );
  nnd2s1 U8438 ( .DIN1(n8257), .DIN2(n8258), .Q(n8247) );
  nnd2s1 U8439 ( .DIN1(n8259), .DIN2(n8260), .Q(n8258) );
  nnd2s1 U8440 ( .DIN1(n8034), .DIN2(n8261), .Q(n8245) );
  nnd2s1 U8441 ( .DIN1(n7853), .DIN2(n8079), .Q(n8244) );
  nnd2s1 U8442 ( .DIN1(n8022), .DIN2(n8061), .Q(n8243) );
  nnd3s1 U8443 ( .DIN1(n8014), .DIN2(n8262), .DIN3(n7849), .Q(n8241) );
  nor4s1 U8444 ( .DIN1(n8263), .DIN2(n8264), .DIN3(n8265), .DIN4(n8266), 
        .Q(n7849) );
  nnd4s1 U8445 ( .DIN1(n8267), .DIN2(n8268), .DIN3(n8269), .DIN4(n8270), 
        .Q(n8266) );
  nnd2s1 U8446 ( .DIN1(n8072), .DIN2(n8271), .Q(n8270) );
  nnd2s1 U8447 ( .DIN1(n7852), .DIN2(n8254), .Q(n8269) );
  nnd2s1 U8448 ( .DIN1(n8023), .DIN2(n7870), .Q(n8268) );
  nnd2s1 U8449 ( .DIN1(n8049), .DIN2(n8272), .Q(n8267) );
  nnd3s1 U8450 ( .DIN1(n8273), .DIN2(n8274), .DIN3(n8275), .Q(n8265) );
  nnd2s1 U8451 ( .DIN1(n8052), .DIN2(n8276), .Q(n8275) );
  nnd2s1 U8452 ( .DIN1(n8277), .DIN2(n8278), .Q(n8276) );
  nnd2s1 U8453 ( .DIN1(n8078), .DIN2(n8279), .Q(n8274) );
  nnd2s1 U8454 ( .DIN1(n8280), .DIN2(n8281), .Q(n8279) );
  nnd2s1 U8455 ( .DIN1(n8030), .DIN2(n8282), .Q(n8273) );
  nnd2s1 U8456 ( .DIN1(n8283), .DIN2(n8074), .Q(n8282) );
  nor2s1 U8457 ( .DIN1(n8051), .DIN2(n8284), .Q(n8264) );
  and2s1 U8458 ( .DIN1(n8036), .DIN2(n8285), .Q(n8263) );
  nnd3s1 U8459 ( .DIN1(n7878), .DIN2(n8286), .DIN3(n7868), .Q(n8285) );
  nor3s1 U8460 ( .DIN1(n8287), .DIN2(n8288), .DIN3(n8289), .Q(n8014) );
  nnd4s1 U8461 ( .DIN1(n8290), .DIN2(n8291), .DIN3(n7850), .DIN4(n8292), 
        .Q(n8289) );
  and3s1 U8462 ( .DIN1(n8293), .DIN2(n8294), .DIN3(n8295), .Q(n8292) );
  nnd2s1 U8463 ( .DIN1(n8023), .DIN2(n8021), .Q(n8294) );
  nnd2s1 U8464 ( .DIN1(n8072), .DIN2(n8022), .Q(n8293) );
  nor2s1 U8465 ( .DIN1(n8296), .DIN2(n8297), .Q(n7850) );
  nnd4s1 U8466 ( .DIN1(n8298), .DIN2(n8299), .DIN3(n8300), .DIN4(n8301), 
        .Q(n8297) );
  nnd2s1 U8467 ( .DIN1(n7866), .DIN2(n8302), .Q(n8301) );
  nnd2s1 U8468 ( .DIN1(n7861), .DIN2(n8303), .Q(n8300) );
  nnd2s1 U8469 ( .DIN1(n8254), .DIN2(n8261), .Q(n8299) );
  nnd2s1 U8470 ( .DIN1(n8030), .DIN2(n8042), .Q(n8298) );
  nnd4s1 U8471 ( .DIN1(n8304), .DIN2(n8305), .DIN3(n8306), .DIN4(n8307), 
        .Q(n8296) );
  nnd2s1 U8472 ( .DIN1(n8062), .DIN2(n8308), .Q(n8307) );
  nnd2s1 U8473 ( .DIN1(n8252), .DIN2(n8260), .Q(n8308) );
  nnd2s1 U8474 ( .DIN1(n7852), .DIN2(n8303), .Q(n8306) );
  nnd2s1 U8475 ( .DIN1(n8052), .DIN2(n8309), .Q(n8305) );
  nnd2s1 U8476 ( .DIN1(n7877), .DIN2(n8051), .Q(n8309) );
  nnd2s1 U8477 ( .DIN1(n8310), .DIN2(n8311), .Q(n8304) );
  nnd3s1 U8478 ( .DIN1(n8059), .DIN2(n8253), .DIN3(n8312), .Q(n8311) );
  nnd3s1 U8479 ( .DIN1(n8313), .DIN2(n8314), .DIN3(n8315), .Q(n8288) );
  nnd2s1 U8480 ( .DIN1(n8316), .DIN2(n8037), .Q(n8315) );
  nnd2s1 U8481 ( .DIN1(n8062), .DIN2(n8317), .Q(n8314) );
  nnd3s1 U8482 ( .DIN1(n8318), .DIN2(n8048), .DIN3(n7860), .Q(n8317) );
  nor2s1 U8483 ( .DIN1(n7870), .DIN2(n8069), .Q(n7860) );
  nnd2s1 U8484 ( .DIN1(n8310), .DIN2(n7870), .Q(n8313) );
  nnd3s1 U8485 ( .DIN1(n8319), .DIN2(n8320), .DIN3(n8321), .Q(n8287) );
  nnd2s1 U8486 ( .DIN1(n7866), .DIN2(n8322), .Q(n8321) );
  nnd2s1 U8487 ( .DIN1(n8323), .DIN2(n7859), .Q(n8322) );
  nnd2s1 U8488 ( .DIN1(n8078), .DIN2(n8324), .Q(n8320) );
  nnd2s1 U8489 ( .DIN1(n8074), .DIN2(n8278), .Q(n8324) );
  nnd2s1 U8490 ( .DIN1(n7853), .DIN2(n8325), .Q(n8319) );
  nnd2s1 U8491 ( .DIN1(n8051), .DIN2(n8278), .Q(n8325) );
  nnd3s1 U8492 ( .DIN1(n8326), .DIN2(n8327), .DIN3(n8328), .Q(n8240) );
  or3s1 U8493 ( .DIN1(n8329), .DIN2(n8330), .DIN3(n8331), .Q(n7733) );
  nnd4s1 U8494 ( .DIN1(n8332), .DIN2(n8333), .DIN3(n8089), .DIN4(n8334), 
        .Q(n8331) );
  and4s1 U8495 ( .DIN1(n8335), .DIN2(n8336), .DIN3(n8337), .DIN4(n7889), 
        .Q(n8334) );
  nnd2s1 U8496 ( .DIN1(n8338), .DIN2(n8106), .Q(n7889) );
  nnd2s1 U8497 ( .DIN1(n8102), .DIN2(n8339), .Q(n8337) );
  nnd2s1 U8498 ( .DIN1(n8340), .DIN2(n7893), .Q(n8336) );
  nor2s1 U8499 ( .DIN1(n8341), .DIN2(n8342), .Q(n8089) );
  nnd4s1 U8500 ( .DIN1(n8343), .DIN2(n8344), .DIN3(n8345), .DIN4(n8346), 
        .Q(n8342) );
  or2s1 U8501 ( .DIN1(n8347), .DIN2(n8348), .Q(n8346) );
  nnd2s1 U8502 ( .DIN1(n8340), .DIN2(n8349), .Q(n8345) );
  nnd2s1 U8503 ( .DIN1(n8338), .DIN2(n7891), .Q(n8344) );
  nnd2s1 U8504 ( .DIN1(n7903), .DIN2(n8350), .Q(n8343) );
  nnd4s1 U8505 ( .DIN1(n8351), .DIN2(n8352), .DIN3(n8353), .DIN4(n8354), 
        .Q(n8341) );
  nnd2s1 U8506 ( .DIN1(n7902), .DIN2(n8355), .Q(n8354) );
  nnd2s1 U8507 ( .DIN1(n8108), .DIN2(n8356), .Q(n8355) );
  nnd2s1 U8508 ( .DIN1(n8357), .DIN2(n8358), .Q(n8353) );
  nnd2s1 U8509 ( .DIN1(n8104), .DIN2(n8359), .Q(n8358) );
  nnd2s1 U8510 ( .DIN1(n8339), .DIN2(n8360), .Q(n8352) );
  nnd2s1 U8511 ( .DIN1(n8361), .DIN2(n8362), .Q(n8360) );
  nnd2s1 U8512 ( .DIN1(n7912), .DIN2(n8363), .Q(n8351) );
  nnd3s1 U8513 ( .DIN1(n8364), .DIN2(n8108), .DIN3(n8365), .Q(n8363) );
  nnd4s1 U8514 ( .DIN1(n8366), .DIN2(n8367), .DIN3(n8368), .DIN4(n8369), 
        .Q(n8330) );
  nnd2s1 U8515 ( .DIN1(n8370), .DIN2(n8371), .Q(n8369) );
  nnd2s1 U8516 ( .DIN1(n7903), .DIN2(n8372), .Q(n8368) );
  nnd2s1 U8517 ( .DIN1(n7890), .DIN2(n8373), .Q(n8367) );
  nnd2s1 U8518 ( .DIN1(n8090), .DIN2(n8350), .Q(n8366) );
  nnd4s1 U8519 ( .DIN1(n8374), .DIN2(n8375), .DIN3(n8376), .DIN4(n8377), 
        .Q(n8329) );
  nnd2s1 U8520 ( .DIN1(n7920), .DIN2(n8378), .Q(n8377) );
  nnd2s1 U8521 ( .DIN1(n8105), .DIN2(n8379), .Q(n8378) );
  nnd2s1 U8522 ( .DIN1(n8380), .DIN2(n8381), .Q(n8376) );
  nnd2s1 U8523 ( .DIN1(n7916), .DIN2(n8382), .Q(n8375) );
  nnd2s1 U8524 ( .DIN1(n8383), .DIN2(n7911), .Q(n8382) );
  nnd2s1 U8525 ( .DIN1(n7900), .DIN2(n8384), .Q(n8374) );
  nnd2s1 U8526 ( .DIN1(n8385), .DIN2(n1603), .Q(n8114) );
  xor2s1 U8527 ( .DIN1(w0[5]), .DIN2(text_in_r[101]), .Q(n8385) );
  nnd2s1 U8528 ( .DIN1(n8386), .DIN2(n8387), .Q(N230) );
  nnd2s1 U8529 ( .DIN1(n8388), .DIN2(n1623), .Q(n8387) );
  xor2s1 U8530 ( .DIN1(n8389), .DIN2(n8390), .Q(n8388) );
  xor2s1 U8531 ( .DIN1(n8391), .DIN2(n8392), .Q(n8390) );
  xnr2s1 U8532 ( .DIN1(n5705), .DIN2(n7577), .Q(n8392) );
  xnr2s1 U8533 ( .DIN1(n5706), .DIN2(n5081), .Q(n7577) );
  hi1s1 U8534 ( .DIN(n7678), .Q(n5081) );
  or3s1 U8535 ( .DIN1(n8393), .DIN2(n8394), .DIN3(n8395), .Q(n7678) );
  nnd4s1 U8536 ( .DIN1(n8122), .DIN2(n8396), .DIN3(n7944), .DIN4(n8397), 
        .Q(n8395) );
  and3s1 U8537 ( .DIN1(n8398), .DIN2(n8399), .DIN3(n8400), .Q(n8397) );
  nor4s1 U8538 ( .DIN1(n8401), .DIN2(n8402), .DIN3(n8403), .DIN4(n8404), 
        .Q(n7944) );
  nnd4s1 U8539 ( .DIN1(n8405), .DIN2(n8406), .DIN3(n8407), .DIN4(n8408), 
        .Q(n8404) );
  nnd2s1 U8540 ( .DIN1(n7947), .DIN2(n7817), .Q(n8408) );
  nnd2s1 U8541 ( .DIN1(n8130), .DIN2(n8409), .Q(n8406) );
  nnd2s1 U8542 ( .DIN1(n8147), .DIN2(n7818), .Q(n8405) );
  nnd3s1 U8543 ( .DIN1(n8410), .DIN2(n8411), .DIN3(n8412), .Q(n8403) );
  nnd2s1 U8544 ( .DIN1(n8160), .DIN2(n8413), .Q(n8412) );
  nnd2s1 U8545 ( .DIN1(n8414), .DIN2(n7833), .Q(n8413) );
  nnd2s1 U8546 ( .DIN1(n7831), .DIN2(n8415), .Q(n8411) );
  nnd2s1 U8547 ( .DIN1(n8416), .DIN2(n8169), .Q(n8415) );
  nnd2s1 U8548 ( .DIN1(n8128), .DIN2(n8417), .Q(n8410) );
  nnd2s1 U8549 ( .DIN1(n8418), .DIN2(n7830), .Q(n8417) );
  nor2s1 U8550 ( .DIN1(n8419), .DIN2(n8420), .Q(n8402) );
  and2s1 U8551 ( .DIN1(n7810), .DIN2(n8421), .Q(n8401) );
  nnd3s1 U8552 ( .DIN1(n8422), .DIN2(n7965), .DIN3(n7962), .Q(n8421) );
  nor3s1 U8553 ( .DIN1(n8423), .DIN2(n8424), .DIN3(n8425), .Q(n8122) );
  nnd4s1 U8554 ( .DIN1(n8426), .DIN2(n8427), .DIN3(n7945), .DIN4(n8428), 
        .Q(n8425) );
  and3s1 U8555 ( .DIN1(n8429), .DIN2(n8430), .DIN3(n8431), .Q(n8428) );
  nnd2s1 U8556 ( .DIN1(n8128), .DIN2(n8140), .Q(n8431) );
  nnd2s1 U8557 ( .DIN1(n8432), .DIN2(n7811), .Q(n8430) );
  nnd2s1 U8558 ( .DIN1(n8433), .DIN2(n7822), .Q(n8429) );
  nor2s1 U8559 ( .DIN1(n8434), .DIN2(n8435), .Q(n7945) );
  nnd4s1 U8560 ( .DIN1(n8436), .DIN2(n8437), .DIN3(n8438), .DIN4(n8439), 
        .Q(n8435) );
  nnd2s1 U8561 ( .DIN1(n7959), .DIN2(n8440), .Q(n8439) );
  nnd2s1 U8562 ( .DIN1(n7835), .DIN2(n8441), .Q(n8438) );
  nnd2s1 U8563 ( .DIN1(n7817), .DIN2(n8442), .Q(n8437) );
  nnd2s1 U8564 ( .DIN1(n7831), .DIN2(n7948), .Q(n8436) );
  nnd4s1 U8565 ( .DIN1(n8443), .DIN2(n8444), .DIN3(n8445), .DIN4(n8446), 
        .Q(n8434) );
  nnd2s1 U8566 ( .DIN1(n7947), .DIN2(n8441), .Q(n8446) );
  nnd2s1 U8567 ( .DIN1(n7821), .DIN2(n8447), .Q(n8445) );
  nnd2s1 U8568 ( .DIN1(n7966), .DIN2(n8149), .Q(n8447) );
  nnd2s1 U8569 ( .DIN1(n7809), .DIN2(n8448), .Q(n8444) );
  nnd2s1 U8570 ( .DIN1(n8449), .DIN2(n8450), .Q(n8448) );
  nnd2s1 U8571 ( .DIN1(n8432), .DIN2(n8451), .Q(n8443) );
  nnd3s1 U8572 ( .DIN1(n8452), .DIN2(n8453), .DIN3(n7838), .Q(n8451) );
  nnd3s1 U8573 ( .DIN1(n8454), .DIN2(n8455), .DIN3(n7813), .Q(n8424) );
  nnd2s1 U8574 ( .DIN1(n8147), .DIN2(n8139), .Q(n7813) );
  nnd2s1 U8575 ( .DIN1(n7809), .DIN2(n8456), .Q(n8455) );
  nnd3s1 U8576 ( .DIN1(n8457), .DIN2(n8152), .DIN3(n7954), .Q(n8456) );
  nor2s1 U8577 ( .DIN1(n8170), .DIN2(n7811), .Q(n7954) );
  nnd2s1 U8578 ( .DIN1(n8129), .DIN2(n7839), .Q(n8454) );
  nnd3s1 U8579 ( .DIN1(n8458), .DIN2(n8459), .DIN3(n8460), .Q(n8423) );
  nnd2s1 U8580 ( .DIN1(n8160), .DIN2(n8461), .Q(n8460) );
  nnd2s1 U8581 ( .DIN1(n8137), .DIN2(n8169), .Q(n8461) );
  nnd2s1 U8582 ( .DIN1(n7819), .DIN2(n8462), .Q(n8459) );
  nnd2s1 U8583 ( .DIN1(n8149), .DIN2(n8137), .Q(n8462) );
  nnd2s1 U8584 ( .DIN1(n7959), .DIN2(n8463), .Q(n8458) );
  nnd2s1 U8585 ( .DIN1(n8416), .DIN2(n7966), .Q(n8463) );
  nnd3s1 U8586 ( .DIN1(n8464), .DIN2(n8465), .DIN3(n8466), .Q(n8394) );
  nnd2s1 U8587 ( .DIN1(n8130), .DIN2(n8442), .Q(n8466) );
  nnd2s1 U8588 ( .DIN1(n7819), .DIN2(n8161), .Q(n8465) );
  nnd2s1 U8589 ( .DIN1(n8129), .DIN2(n8162), .Q(n8464) );
  nnd4s1 U8590 ( .DIN1(n8467), .DIN2(n8468), .DIN3(n8469), .DIN4(n8470), 
        .Q(n8393) );
  nnd2s1 U8591 ( .DIN1(n7817), .DIN2(n8471), .Q(n8470) );
  nnd2s1 U8592 ( .DIN1(n8146), .DIN2(n7962), .Q(n8471) );
  nnd2s1 U8593 ( .DIN1(n7947), .DIN2(n8472), .Q(n8469) );
  nnd2s1 U8594 ( .DIN1(n8453), .DIN2(n8449), .Q(n8472) );
  nnd2s1 U8595 ( .DIN1(n7963), .DIN2(n8473), .Q(n8468) );
  nnd2s1 U8596 ( .DIN1(n7827), .DIN2(n8474), .Q(n8467) );
  nnd2s1 U8597 ( .DIN1(n8475), .DIN2(n8450), .Q(n8474) );
  or3s1 U8598 ( .DIN1(n8476), .DIN2(n8477), .DIN3(n8478), .Q(n5706) );
  nnd4s1 U8599 ( .DIN1(n8178), .DIN2(n8479), .DIN3(n7978), .DIN4(n8480), 
        .Q(n8478) );
  and3s1 U8600 ( .DIN1(n8481), .DIN2(n8482), .DIN3(n8483), .Q(n8480) );
  nor4s1 U8601 ( .DIN1(n8484), .DIN2(n8485), .DIN3(n8486), .DIN4(n8487), 
        .Q(n7978) );
  nnd4s1 U8602 ( .DIN1(n8488), .DIN2(n8489), .DIN3(n8490), .DIN4(n8491), 
        .Q(n8487) );
  nnd2s1 U8603 ( .DIN1(n7981), .DIN2(n8492), .Q(n8491) );
  nnd2s1 U8604 ( .DIN1(n8186), .DIN2(n8493), .Q(n8489) );
  nnd2s1 U8605 ( .DIN1(n8207), .DIN2(n8494), .Q(n8488) );
  nnd3s1 U8606 ( .DIN1(n8495), .DIN2(n8496), .DIN3(n8497), .Q(n8486) );
  nnd2s1 U8607 ( .DIN1(n8221), .DIN2(n8498), .Q(n8497) );
  nnd2s1 U8608 ( .DIN1(n8499), .DIN2(n8500), .Q(n8498) );
  nnd2s1 U8609 ( .DIN1(n8213), .DIN2(n8501), .Q(n8496) );
  nnd2s1 U8610 ( .DIN1(n8502), .DIN2(n8232), .Q(n8501) );
  nnd2s1 U8611 ( .DIN1(n8197), .DIN2(n8503), .Q(n8495) );
  nnd2s1 U8612 ( .DIN1(n8504), .DIN2(n8237), .Q(n8503) );
  nor2s1 U8613 ( .DIN1(n8505), .DIN2(n8506), .Q(n8485) );
  and2s1 U8614 ( .DIN1(n7983), .DIN2(n8507), .Q(n8484) );
  nnd3s1 U8615 ( .DIN1(n8508), .DIN2(n8003), .DIN3(n8000), .Q(n8507) );
  nor3s1 U8616 ( .DIN1(n8509), .DIN2(n8510), .DIN3(n8511), .Q(n8178) );
  nnd4s1 U8617 ( .DIN1(n8512), .DIN2(n8513), .DIN3(n7979), .DIN4(n8514), 
        .Q(n8511) );
  and3s1 U8618 ( .DIN1(n8515), .DIN2(n8516), .DIN3(n8517), .Q(n8514) );
  nnd2s1 U8619 ( .DIN1(n8197), .DIN2(n8199), .Q(n8517) );
  nnd2s1 U8620 ( .DIN1(n8518), .DIN2(n8005), .Q(n8516) );
  nnd2s1 U8621 ( .DIN1(n8519), .DIN2(n8198), .Q(n8515) );
  nor2s1 U8622 ( .DIN1(n8520), .DIN2(n8521), .Q(n7979) );
  nnd4s1 U8623 ( .DIN1(n8522), .DIN2(n8523), .DIN3(n8524), .DIN4(n8525), 
        .Q(n8521) );
  nnd2s1 U8624 ( .DIN1(n7997), .DIN2(n8526), .Q(n8525) );
  nnd2s1 U8625 ( .DIN1(n7992), .DIN2(n8527), .Q(n8524) );
  nnd2s1 U8626 ( .DIN1(n8492), .DIN2(n8528), .Q(n8523) );
  nnd2s1 U8627 ( .DIN1(n8213), .DIN2(n7984), .Q(n8522) );
  nnd4s1 U8628 ( .DIN1(n8529), .DIN2(n8530), .DIN3(n8531), .DIN4(n8532), 
        .Q(n8520) );
  nnd2s1 U8629 ( .DIN1(n7981), .DIN2(n8527), .Q(n8532) );
  nnd2s1 U8630 ( .DIN1(n8204), .DIN2(n8533), .Q(n8531) );
  nnd2s1 U8631 ( .DIN1(n8004), .DIN2(n8209), .Q(n8533) );
  nnd2s1 U8632 ( .DIN1(n8224), .DIN2(n8534), .Q(n8530) );
  nnd2s1 U8633 ( .DIN1(n8535), .DIN2(n8536), .Q(n8534) );
  nnd2s1 U8634 ( .DIN1(n8518), .DIN2(n8537), .Q(n8529) );
  nnd3s1 U8635 ( .DIN1(n8538), .DIN2(n8539), .DIN3(n8540), .Q(n8537) );
  nnd3s1 U8636 ( .DIN1(n8541), .DIN2(n8542), .DIN3(n8543), .Q(n8510) );
  nnd2s1 U8637 ( .DIN1(n8224), .DIN2(n8544), .Q(n8542) );
  nnd3s1 U8638 ( .DIN1(n8545), .DIN2(n8212), .DIN3(n7991), .Q(n8544) );
  nor2s1 U8639 ( .DIN1(n8233), .DIN2(n8005), .Q(n7991) );
  nnd2s1 U8640 ( .DIN1(n8185), .DIN2(n8230), .Q(n8541) );
  nnd3s1 U8641 ( .DIN1(n8546), .DIN2(n8547), .DIN3(n8548), .Q(n8509) );
  nnd2s1 U8642 ( .DIN1(n8221), .DIN2(n8549), .Q(n8548) );
  nnd2s1 U8643 ( .DIN1(n8194), .DIN2(n8232), .Q(n8549) );
  nnd2s1 U8644 ( .DIN1(n7982), .DIN2(n8550), .Q(n8547) );
  nnd2s1 U8645 ( .DIN1(n8209), .DIN2(n8194), .Q(n8550) );
  nnd2s1 U8646 ( .DIN1(n7997), .DIN2(n8551), .Q(n8546) );
  nnd2s1 U8647 ( .DIN1(n8502), .DIN2(n8004), .Q(n8551) );
  nnd3s1 U8648 ( .DIN1(n8552), .DIN2(n8553), .DIN3(n8554), .Q(n8477) );
  nnd2s1 U8649 ( .DIN1(n8186), .DIN2(n8528), .Q(n8554) );
  nnd2s1 U8650 ( .DIN1(n7982), .DIN2(n8222), .Q(n8553) );
  nnd2s1 U8651 ( .DIN1(n8185), .DIN2(n8223), .Q(n8552) );
  nnd4s1 U8652 ( .DIN1(n8555), .DIN2(n8556), .DIN3(n8557), .DIN4(n8558), 
        .Q(n8476) );
  nnd2s1 U8653 ( .DIN1(n8492), .DIN2(n8559), .Q(n8558) );
  nnd2s1 U8654 ( .DIN1(n8206), .DIN2(n8000), .Q(n8559) );
  nnd2s1 U8655 ( .DIN1(n7981), .DIN2(n8560), .Q(n8557) );
  nnd2s1 U8656 ( .DIN1(n8539), .DIN2(n8535), .Q(n8560) );
  nnd2s1 U8657 ( .DIN1(n8001), .DIN2(n8561), .Q(n8556) );
  nnd2s1 U8658 ( .DIN1(n8562), .DIN2(n8563), .Q(n8555) );
  nnd2s1 U8659 ( .DIN1(n8564), .DIN2(n8536), .Q(n8563) );
  xor2s1 U8660 ( .DIN1(n7741), .DIN2(n8565), .Q(n8389) );
  xor2s1 U8661 ( .DIN1(n1472), .DIN2(n5033), .Q(n8565) );
  or3s1 U8662 ( .DIN1(n8566), .DIN2(n8567), .DIN3(n8568), .Q(n5033) );
  nnd4s1 U8663 ( .DIN1(n8569), .DIN2(n8570), .DIN3(n7847), .DIN4(n8571), 
        .Q(n8568) );
  and3s1 U8664 ( .DIN1(n8015), .DIN2(n8290), .DIN3(n8262), .Q(n8571) );
  nor4s1 U8665 ( .DIN1(n8572), .DIN2(n8573), .DIN3(n8574), .DIN4(n8575), 
        .Q(n8262) );
  nnd4s1 U8666 ( .DIN1(n8576), .DIN2(n8577), .DIN3(n8578), .DIN4(n8579), 
        .Q(n8575) );
  nor2s1 U8667 ( .DIN1(n8580), .DIN2(n8581), .Q(n8579) );
  nor2s1 U8668 ( .DIN1(n8284), .DIN2(n8074), .Q(n8581) );
  nor2s1 U8669 ( .DIN1(n8060), .DIN2(n8253), .Q(n8580) );
  or2s1 U8670 ( .DIN1(n8277), .DIN2(n8582), .Q(n8578) );
  nnd2s1 U8671 ( .DIN1(n8316), .DIN2(n8583), .Q(n8577) );
  nnd3s1 U8672 ( .DIN1(n8278), .DIN2(n7859), .DIN3(n7869), .Q(n8583) );
  nnd2s1 U8673 ( .DIN1(n8584), .DIN2(n8585), .Q(n8576) );
  nnd3s1 U8674 ( .DIN1(n8586), .DIN2(n8044), .DIN3(n8059), .Q(n8585) );
  nnd3s1 U8675 ( .DIN1(n8587), .DIN2(n8588), .DIN3(n8589), .Q(n8574) );
  nnd2s1 U8676 ( .DIN1(n8064), .DIN2(n8021), .Q(n8589) );
  nnd2s1 U8677 ( .DIN1(n8078), .DIN2(n8035), .Q(n8588) );
  nnd2s1 U8678 ( .DIN1(n8254), .DIN2(n8042), .Q(n8587) );
  nor2s1 U8679 ( .DIN1(n8590), .DIN2(n7857), .Q(n8573) );
  nor2s1 U8680 ( .DIN1(n8252), .DIN2(n8591), .Q(n8572) );
  nor4s1 U8681 ( .DIN1(n8592), .DIN2(n8593), .DIN3(n8594), .DIN4(n8595), 
        .Q(n8290) );
  nnd4s1 U8682 ( .DIN1(n8596), .DIN2(n8597), .DIN3(n8598), .DIN4(n8599), 
        .Q(n8595) );
  nnd2s1 U8683 ( .DIN1(n8036), .DIN2(n8272), .Q(n8599) );
  nor2s1 U8684 ( .DIN1(n8600), .DIN2(n8601), .Q(n8598) );
  nor2s1 U8685 ( .DIN1(n8586), .DIN2(n8277), .Q(n8601) );
  nor2s1 U8686 ( .DIN1(n8054), .DIN2(n8284), .Q(n8600) );
  nnd2s1 U8687 ( .DIN1(n8072), .DIN2(n8042), .Q(n8597) );
  nnd2s1 U8688 ( .DIN1(n7853), .DIN2(n8022), .Q(n8596) );
  nnd3s1 U8689 ( .DIN1(n8602), .DIN2(n8603), .DIN3(n8604), .Q(n8594) );
  nnd2s1 U8690 ( .DIN1(n7852), .DIN2(n8605), .Q(n8604) );
  nnd2s1 U8691 ( .DIN1(n8259), .DIN2(n8044), .Q(n8605) );
  nnd2s1 U8692 ( .DIN1(n8021), .DIN2(n8606), .Q(n8603) );
  nnd2s1 U8693 ( .DIN1(n8607), .DIN2(n8278), .Q(n8606) );
  nnd2s1 U8694 ( .DIN1(n8064), .DIN2(n8608), .Q(n8602) );
  nnd2s1 U8695 ( .DIN1(n8318), .DIN2(n8077), .Q(n8608) );
  nor2s1 U8696 ( .DIN1(n8609), .DIN2(n8076), .Q(n8593) );
  nor2s1 U8697 ( .DIN1(n8271), .DIN2(n8257), .Q(n8609) );
  nor2s1 U8698 ( .DIN1(n8610), .DIN2(n7868), .Q(n8592) );
  nor2s1 U8699 ( .DIN1(n8316), .DIN2(n8069), .Q(n8610) );
  nor4s1 U8700 ( .DIN1(n8611), .DIN2(n8612), .DIN3(n8613), .DIN4(n8614), 
        .Q(n8015) );
  nnd4s1 U8701 ( .DIN1(n8615), .DIN2(n8616), .DIN3(n8617), .DIN4(n8618), 
        .Q(n8614) );
  nor2s1 U8702 ( .DIN1(n8619), .DIN2(n8620), .Q(n8617) );
  nor2s1 U8703 ( .DIN1(n8260), .DIN2(n7878), .Q(n8620) );
  nor2s1 U8704 ( .DIN1(n8032), .DIN2(n8284), .Q(n8619) );
  nnd2s1 U8705 ( .DIN1(n8254), .DIN2(n8272), .Q(n8616) );
  nnd2s1 U8706 ( .DIN1(n8023), .DIN2(n8049), .Q(n8615) );
  nnd3s1 U8707 ( .DIN1(n8621), .DIN2(n8622), .DIN3(n8623), .Q(n8613) );
  nnd2s1 U8708 ( .DIN1(n7853), .DIN2(n8624), .Q(n8623) );
  nnd2s1 U8709 ( .DIN1(n7861), .DIN2(n8625), .Q(n8622) );
  nnd2s1 U8710 ( .DIN1(n8044), .DIN2(n8260), .Q(n8625) );
  nnd2s1 U8711 ( .DIN1(n8316), .DIN2(n8626), .Q(n8621) );
  nnd3s1 U8712 ( .DIN1(n8286), .DIN2(n8277), .DIN3(n8627), .Q(n8626) );
  nor2s1 U8713 ( .DIN1(n8045), .DIN2(n7877), .Q(n8612) );
  nor2s1 U8714 ( .DIN1(n7872), .DIN2(n8076), .Q(n8611) );
  nor3s1 U8715 ( .DIN1(n8628), .DIN2(n8629), .DIN3(n8630), .Q(n7847) );
  nnd4s1 U8716 ( .DIN1(n8291), .DIN2(n8017), .DIN3(n8328), .DIN4(n8631), 
        .Q(n8630) );
  and3s1 U8717 ( .DIN1(n8632), .DIN2(n8633), .DIN3(n8634), .Q(n8631) );
  nnd2s1 U8718 ( .DIN1(n7853), .DIN2(n8257), .Q(n8634) );
  nnd2s1 U8719 ( .DIN1(n8034), .DIN2(n8272), .Q(n8633) );
  nnd2s1 U8720 ( .DIN1(n8062), .DIN2(n7875), .Q(n8632) );
  nor4s1 U8721 ( .DIN1(n8635), .DIN2(n8636), .DIN3(n8637), .DIN4(n8638), 
        .Q(n8328) );
  nnd4s1 U8722 ( .DIN1(n8639), .DIN2(n8640), .DIN3(n8641), .DIN4(n8642), 
        .Q(n8638) );
  nnd2s1 U8723 ( .DIN1(n7875), .DIN2(n8643), .Q(n8642) );
  nor2s1 U8724 ( .DIN1(n8644), .DIN2(n8645), .Q(n8641) );
  nor2s1 U8725 ( .DIN1(n8646), .DIN2(n8286), .Q(n8645) );
  nor2s1 U8726 ( .DIN1(n8034), .DIN2(n8254), .Q(n8646) );
  nor2s1 U8727 ( .DIN1(n8647), .DIN2(n8077), .Q(n8644) );
  nor2s1 U8728 ( .DIN1(n8062), .DIN2(n7874), .Q(n8647) );
  nnd2s1 U8729 ( .DIN1(n8257), .DIN2(n8648), .Q(n8640) );
  nnd3s1 U8730 ( .DIN1(n8045), .DIN2(n8252), .DIN3(n8312), .Q(n8648) );
  nnd2s1 U8731 ( .DIN1(n8069), .DIN2(n8649), .Q(n8639) );
  nnd3s1 U8732 ( .DIN1(n8650), .DIN2(n8651), .DIN3(n8652), .Q(n8637) );
  nnd2s1 U8733 ( .DIN1(n8316), .DIN2(n8271), .Q(n8652) );
  nnd2s1 U8734 ( .DIN1(n8064), .DIN2(n8078), .Q(n8650) );
  nor2s1 U8735 ( .DIN1(n8259), .DIN2(n8277), .Q(n8636) );
  nor2s1 U8736 ( .DIN1(n8076), .DIN2(n8074), .Q(n8635) );
  nor4s1 U8737 ( .DIN1(n8653), .DIN2(n8654), .DIN3(n8655), .DIN4(n8656), 
        .Q(n8017) );
  nnd4s1 U8738 ( .DIN1(n8657), .DIN2(n8658), .DIN3(n8659), .DIN4(n8660), 
        .Q(n8656) );
  nnd2s1 U8739 ( .DIN1(n8257), .DIN2(n8078), .Q(n8660) );
  nnd2s1 U8740 ( .DIN1(n8069), .DIN2(n8584), .Q(n8659) );
  nnd2s1 U8741 ( .DIN1(n8072), .DIN2(n8272), .Q(n8658) );
  nnd2s1 U8742 ( .DIN1(n7875), .DIN2(n8035), .Q(n8657) );
  nnd3s1 U8743 ( .DIN1(n8661), .DIN2(n8662), .DIN3(n8663), .Q(n8655) );
  nnd2s1 U8744 ( .DIN1(n7870), .DIN2(n8664), .Q(n8663) );
  nnd2s1 U8745 ( .DIN1(n8323), .DIN2(n8051), .Q(n8664) );
  nor2s1 U8746 ( .DIN1(n8064), .DIN2(n8271), .Q(n8323) );
  nnd2s1 U8747 ( .DIN1(n8063), .DIN2(n8665), .Q(n8662) );
  nnd2s1 U8748 ( .DIN1(n8607), .DIN2(n8051), .Q(n8665) );
  nor2s1 U8749 ( .DIN1(n8271), .DIN2(n8649), .Q(n8607) );
  nnd2s1 U8750 ( .DIN1(n8310), .DIN2(n8666), .Q(n8661) );
  nnd2s1 U8751 ( .DIN1(n8259), .DIN2(n8284), .Q(n8666) );
  nor2s1 U8752 ( .DIN1(n8284), .DIN2(n8277), .Q(n8654) );
  nor2s1 U8753 ( .DIN1(n8033), .DIN2(n8260), .Q(n8653) );
  hi1s1 U8754 ( .DIN(n8667), .Q(n8033) );
  nor2s1 U8755 ( .DIN1(n8668), .DIN2(n8669), .Q(n8291) );
  nnd4s1 U8756 ( .DIN1(n8670), .DIN2(n8671), .DIN3(n8672), .DIN4(n8673), 
        .Q(n8669) );
  nnd2s1 U8757 ( .DIN1(n8272), .DIN2(n8674), .Q(n8673) );
  nnd3s1 U8758 ( .DIN1(n8586), .DIN2(n8260), .DIN3(n8045), .Q(n8674) );
  nnd2s1 U8759 ( .DIN1(n8254), .DIN2(n8022), .Q(n8670) );
  nnd4s1 U8760 ( .DIN1(n8675), .DIN2(n8676), .DIN3(n8677), .DIN4(n8678), 
        .Q(n8668) );
  nnd2s1 U8761 ( .DIN1(n8036), .DIN2(n8679), .Q(n8678) );
  nnd2s1 U8762 ( .DIN1(n8310), .DIN2(n8680), .Q(n8677) );
  nnd2s1 U8763 ( .DIN1(n7858), .DIN2(n8252), .Q(n8680) );
  nnd2s1 U8764 ( .DIN1(n8072), .DIN2(n8681), .Q(n8676) );
  nnd2s1 U8765 ( .DIN1(n8682), .DIN2(n7877), .Q(n8681) );
  nnd2s1 U8766 ( .DIN1(n7861), .DIN2(n8683), .Q(n8675) );
  nnd2s1 U8767 ( .DIN1(n8253), .DIN2(n8045), .Q(n8683) );
  nnd3s1 U8768 ( .DIN1(n8684), .DIN2(n8685), .DIN3(n8686), .Q(n8629) );
  nnd2s1 U8769 ( .DIN1(n8030), .DIN2(n8649), .Q(n8686) );
  nnd2s1 U8770 ( .DIN1(n8271), .DIN2(n8687), .Q(n8685) );
  nnd3s1 U8771 ( .DIN1(n8312), .DIN2(n8586), .DIN3(n8688), .Q(n8687) );
  or2s1 U8772 ( .DIN1(n8051), .DIN2(n8689), .Q(n8684) );
  nnd3s1 U8773 ( .DIN1(n8690), .DIN2(n8691), .DIN3(n8692), .Q(n8628) );
  nnd2s1 U8774 ( .DIN1(n7861), .DIN2(n8693), .Q(n8692) );
  nnd2s1 U8775 ( .DIN1(n8059), .DIN2(n8318), .Q(n8693) );
  nnd2s1 U8776 ( .DIN1(n8069), .DIN2(n8694), .Q(n8691) );
  nnd2s1 U8777 ( .DIN1(n8281), .DIN2(n8278), .Q(n8694) );
  nnd2s1 U8778 ( .DIN1(n8049), .DIN2(n8695), .Q(n8690) );
  nnd2s1 U8779 ( .DIN1(n8060), .DIN2(n8286), .Q(n8695) );
  nor2s1 U8780 ( .DIN1(n8037), .DIN2(n8064), .Q(n8060) );
  nnd2s1 U8781 ( .DIN1(n8023), .DIN2(n8030), .Q(n8570) );
  nnd3s1 U8782 ( .DIN1(n8696), .DIN2(n8697), .DIN3(n8698), .Q(n8567) );
  nnd2s1 U8783 ( .DIN1(n7875), .DIN2(n8042), .Q(n8698) );
  nnd2s1 U8784 ( .DIN1(n8699), .DIN2(n8700), .Q(n8697) );
  nnd2s1 U8785 ( .DIN1(n8649), .DIN2(n8072), .Q(n8696) );
  nnd4s1 U8786 ( .DIN1(n8701), .DIN2(n8702), .DIN3(n8703), .DIN4(n8704), 
        .Q(n8566) );
  nnd2s1 U8787 ( .DIN1(n8063), .DIN2(n8705), .Q(n8704) );
  nnd2s1 U8788 ( .DIN1(n7872), .DIN2(n8074), .Q(n8705) );
  nor2s1 U8789 ( .DIN1(n8035), .DIN2(n8022), .Q(n7872) );
  nnd2s1 U8790 ( .DIN1(n8064), .DIN2(n8706), .Q(n8703) );
  nnd2s1 U8791 ( .DIN1(n8312), .DIN2(n8048), .Q(n8706) );
  nnd2s1 U8792 ( .DIN1(n8035), .DIN2(n8707), .Q(n8702) );
  nnd2s1 U8793 ( .DIN1(n8047), .DIN2(n8059), .Q(n8707) );
  nnd2s1 U8794 ( .DIN1(n8257), .DIN2(n8303), .Q(n8701) );
  or3s1 U8795 ( .DIN1(n8708), .DIN2(n8709), .DIN3(n8710), .Q(n7741) );
  nnd4s1 U8796 ( .DIN1(n8332), .DIN2(n8711), .DIN3(n8087), .DIN4(n8712), 
        .Q(n8710) );
  and3s1 U8797 ( .DIN1(n8713), .DIN2(n8714), .DIN3(n8715), .Q(n8712) );
  nor4s1 U8798 ( .DIN1(n8716), .DIN2(n8717), .DIN3(n8718), .DIN4(n8719), 
        .Q(n8087) );
  nnd4s1 U8799 ( .DIN1(n8720), .DIN2(n8721), .DIN3(n8722), .DIN4(n8723), 
        .Q(n8719) );
  nnd2s1 U8800 ( .DIN1(n8090), .DIN2(n7898), .Q(n8723) );
  nnd2s1 U8801 ( .DIN1(n8340), .DIN2(n8724), .Q(n8721) );
  nnd2s1 U8802 ( .DIN1(n8357), .DIN2(n7899), .Q(n8720) );
  nnd3s1 U8803 ( .DIN1(n8725), .DIN2(n8726), .DIN3(n8727), .Q(n8718) );
  nnd2s1 U8804 ( .DIN1(n8370), .DIN2(n8728), .Q(n8727) );
  nnd2s1 U8805 ( .DIN1(n8729), .DIN2(n7914), .Q(n8728) );
  nnd2s1 U8806 ( .DIN1(n7912), .DIN2(n8730), .Q(n8726) );
  nnd2s1 U8807 ( .DIN1(n8731), .DIN2(n8379), .Q(n8730) );
  nnd2s1 U8808 ( .DIN1(n8338), .DIN2(n8732), .Q(n8725) );
  nnd2s1 U8809 ( .DIN1(n8733), .DIN2(n7911), .Q(n8732) );
  nor2s1 U8810 ( .DIN1(n8734), .DIN2(n8735), .Q(n8717) );
  and2s1 U8811 ( .DIN1(n7891), .DIN2(n8736), .Q(n8716) );
  nnd3s1 U8812 ( .DIN1(n8737), .DIN2(n8108), .DIN3(n8105), .Q(n8736) );
  nor3s1 U8813 ( .DIN1(n8738), .DIN2(n8739), .DIN3(n8740), .Q(n8332) );
  nnd4s1 U8814 ( .DIN1(n8741), .DIN2(n8742), .DIN3(n8088), .DIN4(n8743), 
        .Q(n8740) );
  and3s1 U8815 ( .DIN1(n8744), .DIN2(n8745), .DIN3(n8746), .Q(n8743) );
  nnd2s1 U8816 ( .DIN1(n8338), .DIN2(n8350), .Q(n8746) );
  nnd2s1 U8817 ( .DIN1(n8747), .DIN2(n7892), .Q(n8745) );
  nnd2s1 U8818 ( .DIN1(n8748), .DIN2(n7903), .Q(n8744) );
  nor2s1 U8819 ( .DIN1(n8749), .DIN2(n8750), .Q(n8088) );
  nnd4s1 U8820 ( .DIN1(n8751), .DIN2(n8752), .DIN3(n8753), .DIN4(n8754), 
        .Q(n8750) );
  nnd2s1 U8821 ( .DIN1(n8102), .DIN2(n8755), .Q(n8754) );
  nnd2s1 U8822 ( .DIN1(n7916), .DIN2(n8756), .Q(n8753) );
  nnd2s1 U8823 ( .DIN1(n7898), .DIN2(n8757), .Q(n8752) );
  nnd2s1 U8824 ( .DIN1(n7912), .DIN2(n8091), .Q(n8751) );
  nnd4s1 U8825 ( .DIN1(n8758), .DIN2(n8759), .DIN3(n8760), .DIN4(n8761), 
        .Q(n8749) );
  nnd2s1 U8826 ( .DIN1(n8090), .DIN2(n8756), .Q(n8761) );
  nnd2s1 U8827 ( .DIN1(n7902), .DIN2(n8762), .Q(n8760) );
  nnd2s1 U8828 ( .DIN1(n8109), .DIN2(n8359), .Q(n8762) );
  nnd2s1 U8829 ( .DIN1(n7890), .DIN2(n8763), .Q(n8759) );
  nnd2s1 U8830 ( .DIN1(n8764), .DIN2(n8765), .Q(n8763) );
  nnd2s1 U8831 ( .DIN1(n8747), .DIN2(n8766), .Q(n8758) );
  nnd3s1 U8832 ( .DIN1(n8767), .DIN2(n8768), .DIN3(n7919), .Q(n8766) );
  nnd3s1 U8833 ( .DIN1(n8769), .DIN2(n8770), .DIN3(n7894), .Q(n8739) );
  nnd2s1 U8834 ( .DIN1(n8357), .DIN2(n8349), .Q(n7894) );
  nnd2s1 U8835 ( .DIN1(n7890), .DIN2(n8771), .Q(n8770) );
  nnd3s1 U8836 ( .DIN1(n8772), .DIN2(n8362), .DIN3(n8097), .Q(n8771) );
  nor2s1 U8837 ( .DIN1(n8380), .DIN2(n7892), .Q(n8097) );
  nnd2s1 U8838 ( .DIN1(n8339), .DIN2(n7920), .Q(n8769) );
  nnd3s1 U8839 ( .DIN1(n8773), .DIN2(n8774), .DIN3(n8775), .Q(n8738) );
  nnd2s1 U8840 ( .DIN1(n8370), .DIN2(n8776), .Q(n8775) );
  nnd2s1 U8841 ( .DIN1(n8347), .DIN2(n8379), .Q(n8776) );
  nnd2s1 U8842 ( .DIN1(n7900), .DIN2(n8777), .Q(n8774) );
  nnd2s1 U8843 ( .DIN1(n8359), .DIN2(n8347), .Q(n8777) );
  nnd2s1 U8844 ( .DIN1(n8102), .DIN2(n8778), .Q(n8773) );
  nnd2s1 U8845 ( .DIN1(n8731), .DIN2(n8109), .Q(n8778) );
  nnd3s1 U8846 ( .DIN1(n8779), .DIN2(n8780), .DIN3(n8781), .Q(n8709) );
  nnd2s1 U8847 ( .DIN1(n8340), .DIN2(n8757), .Q(n8781) );
  nnd2s1 U8848 ( .DIN1(n7900), .DIN2(n8371), .Q(n8780) );
  nnd2s1 U8849 ( .DIN1(n8339), .DIN2(n8372), .Q(n8779) );
  nnd4s1 U8850 ( .DIN1(n8782), .DIN2(n8783), .DIN3(n8784), .DIN4(n8785), 
        .Q(n8708) );
  nnd2s1 U8851 ( .DIN1(n7898), .DIN2(n8786), .Q(n8785) );
  nnd2s1 U8852 ( .DIN1(n8356), .DIN2(n8105), .Q(n8786) );
  nnd2s1 U8853 ( .DIN1(n8090), .DIN2(n8787), .Q(n8784) );
  nnd2s1 U8854 ( .DIN1(n8768), .DIN2(n8764), .Q(n8787) );
  nnd2s1 U8855 ( .DIN1(n8106), .DIN2(n8788), .Q(n8783) );
  nnd2s1 U8856 ( .DIN1(n7908), .DIN2(n8789), .Q(n8782) );
  nnd2s1 U8857 ( .DIN1(n8790), .DIN2(n8765), .Q(n8789) );
  nnd2s1 U8858 ( .DIN1(n8791), .DIN2(n1603), .Q(n8386) );
  xor2s1 U8859 ( .DIN1(w0[4]), .DIN2(text_in_r[100]), .Q(n8791) );
  and4s1 U8860 ( .DIN1(n1360), .DIN2(n1409), .DIN3(n1526), .DIN4(n8792), 
        .Q(N23) );
  nor2s1 U8861 ( .DIN1(ld), .DIN2(n1449), .Q(n8792) );
  nnd2s1 U8862 ( .DIN1(n8793), .DIN2(n8794), .Q(N229) );
  nnd2s1 U8863 ( .DIN1(n8795), .DIN2(n1623), .Q(n8794) );
  xor2s1 U8864 ( .DIN1(n8796), .DIN2(n8797), .Q(n8795) );
  xor2s1 U8865 ( .DIN1(n8798), .DIN2(n8799), .Q(n8797) );
  xor2s1 U8866 ( .DIN1(n5704), .DIN2(n7763), .Q(n8799) );
  xnr2s1 U8867 ( .DIN1(n5705), .DIN2(n8800), .Q(n7763) );
  hi1s1 U8868 ( .DIN(n5080), .Q(n8800) );
  or3s1 U8869 ( .DIN1(n8801), .DIN2(n8802), .DIN3(n8803), .Q(n5080) );
  nnd4s1 U8870 ( .DIN1(n8804), .DIN2(n8805), .DIN3(n7942), .DIN4(n8806), 
        .Q(n8803) );
  and3s1 U8871 ( .DIN1(n8123), .DIN2(n8426), .DIN3(n8396), .Q(n8806) );
  nor4s1 U8872 ( .DIN1(n8807), .DIN2(n8808), .DIN3(n8809), .DIN4(n8810), 
        .Q(n8396) );
  nnd4s1 U8873 ( .DIN1(n8811), .DIN2(n8812), .DIN3(n8813), .DIN4(n8814), 
        .Q(n8810) );
  nnd2s1 U8874 ( .DIN1(n7822), .DIN2(n7963), .Q(n8814) );
  nor2s1 U8875 ( .DIN1(n8815), .DIN2(n8816), .Q(n8813) );
  nor2s1 U8876 ( .DIN1(n7962), .DIN2(n8817), .Q(n8816) );
  nor2s1 U8877 ( .DIN1(n8818), .DIN2(n8169), .Q(n8815) );
  nnd2s1 U8878 ( .DIN1(n7812), .DIN2(n8140), .Q(n8812) );
  nnd2s1 U8879 ( .DIN1(n8147), .DIN2(n7835), .Q(n8811) );
  nnd3s1 U8880 ( .DIN1(n8819), .DIN2(n8820), .DIN3(n8821), .Q(n8809) );
  nnd2s1 U8881 ( .DIN1(n8170), .DIN2(n8174), .Q(n8821) );
  nnd2s1 U8882 ( .DIN1(n7820), .DIN2(n8822), .Q(n8820) );
  nnd3s1 U8883 ( .DIN1(n8418), .DIN2(n8817), .DIN3(n8452), .Q(n8822) );
  nnd2s1 U8884 ( .DIN1(n8433), .DIN2(n8823), .Q(n8819) );
  nnd3s1 U8885 ( .DIN1(n8137), .DIN2(n7834), .DIN3(n7961), .Q(n8823) );
  nor2s1 U8886 ( .DIN1(n8137), .DIN2(n7838), .Q(n8808) );
  nor2s1 U8887 ( .DIN1(n8824), .DIN2(n8825), .Q(n8807) );
  nor4s1 U8888 ( .DIN1(n8826), .DIN2(n8827), .DIN3(n8828), .DIN4(n8829), 
        .Q(n8426) );
  nnd4s1 U8889 ( .DIN1(n8830), .DIN2(n8831), .DIN3(n8832), .DIN4(n8833), 
        .Q(n8829) );
  nor2s1 U8890 ( .DIN1(n8834), .DIN2(n8835), .Q(n8833) );
  nor2s1 U8891 ( .DIN1(n8817), .DIN2(n8825), .Q(n8835) );
  nor2s1 U8892 ( .DIN1(n8173), .DIN2(n7834), .Q(n8834) );
  nnd2s1 U8893 ( .DIN1(n7948), .DIN2(n7839), .Q(n8831) );
  nnd2s1 U8894 ( .DIN1(n8129), .DIN2(n7819), .Q(n8830) );
  nnd3s1 U8895 ( .DIN1(n8836), .DIN2(n8837), .DIN3(n8838), .Q(n8828) );
  nnd2s1 U8896 ( .DIN1(n8139), .DIN2(n8839), .Q(n8838) );
  nnd2s1 U8897 ( .DIN1(n8453), .DIN2(n8152), .Q(n8839) );
  nnd2s1 U8898 ( .DIN1(n7947), .DIN2(n8840), .Q(n8837) );
  nnd2s1 U8899 ( .DIN1(n8475), .DIN2(n8418), .Q(n8840) );
  nnd2s1 U8900 ( .DIN1(n7821), .DIN2(n8171), .Q(n8836) );
  nnd2s1 U8901 ( .DIN1(n8154), .DIN2(n8419), .Q(n8171) );
  nor2s1 U8902 ( .DIN1(n8841), .DIN2(n7966), .Q(n8827) );
  nor2s1 U8903 ( .DIN1(n7810), .DIN2(n7831), .Q(n8841) );
  nor2s1 U8904 ( .DIN1(n8842), .DIN2(n8450), .Q(n8826) );
  and2s1 U8905 ( .DIN1(n8137), .DIN2(n8843), .Q(n8842) );
  nor4s1 U8906 ( .DIN1(n8844), .DIN2(n8845), .DIN3(n8846), .DIN4(n8847), 
        .Q(n8123) );
  nnd4s1 U8907 ( .DIN1(n8848), .DIN2(n8849), .DIN3(n8850), .DIN4(n8851), 
        .Q(n8847) );
  nnd2s1 U8908 ( .DIN1(n8432), .DIN2(n8140), .Q(n8851) );
  nor2s1 U8909 ( .DIN1(n8852), .DIN2(n8853), .Q(n8850) );
  nor2s1 U8910 ( .DIN1(n8854), .DIN2(n7966), .Q(n8852) );
  nnd2s1 U8911 ( .DIN1(n8128), .DIN2(n8147), .Q(n8849) );
  nnd2s1 U8912 ( .DIN1(n8130), .DIN2(n7827), .Q(n8848) );
  nnd3s1 U8913 ( .DIN1(n8855), .DIN2(n8856), .DIN3(n8857), .Q(n8846) );
  nnd2s1 U8914 ( .DIN1(n7819), .DIN2(n8858), .Q(n8857) );
  nnd2s1 U8915 ( .DIN1(n7835), .DIN2(n8859), .Q(n8856) );
  nnd2s1 U8916 ( .DIN1(n8450), .DIN2(n8418), .Q(n8859) );
  nnd2s1 U8917 ( .DIN1(n8433), .DIN2(n8860), .Q(n8855) );
  nnd3s1 U8918 ( .DIN1(n8422), .DIN2(n8825), .DIN3(n8861), .Q(n8860) );
  nor2s1 U8919 ( .DIN1(n7834), .DIN2(n7838), .Q(n8845) );
  nor2s1 U8920 ( .DIN1(n7968), .DIN2(n7830), .Q(n8844) );
  nor3s1 U8921 ( .DIN1(n8862), .DIN2(n8863), .DIN3(n8864), .Q(n7942) );
  nnd4s1 U8922 ( .DIN1(n8427), .DIN2(n8125), .DIN3(n8400), .DIN4(n8865), 
        .Q(n8864) );
  and3s1 U8923 ( .DIN1(n8866), .DIN2(n8867), .DIN3(n8868), .Q(n8865) );
  nnd2s1 U8924 ( .DIN1(n8130), .DIN2(n7818), .Q(n8868) );
  nnd2s1 U8925 ( .DIN1(n7809), .DIN2(n7963), .Q(n8866) );
  nor4s1 U8926 ( .DIN1(n8869), .DIN2(n8870), .DIN3(n8871), .DIN4(n8872), 
        .Q(n8400) );
  nnd4s1 U8927 ( .DIN1(n8873), .DIN2(n8874), .DIN3(n8875), .DIN4(n8876), 
        .Q(n8872) );
  nnd2s1 U8928 ( .DIN1(n8130), .DIN2(n8877), .Q(n8876) );
  nnd2s1 U8929 ( .DIN1(n8878), .DIN2(n8422), .Q(n8877) );
  nor2s1 U8930 ( .DIN1(n8879), .DIN2(n8880), .Q(n8875) );
  nor2s1 U8931 ( .DIN1(n8881), .DIN2(n8173), .Q(n8880) );
  nor2s1 U8932 ( .DIN1(n7809), .DIN2(n7970), .Q(n8881) );
  nor2s1 U8933 ( .DIN1(n8882), .DIN2(n7837), .Q(n8879) );
  nor2s1 U8934 ( .DIN1(n8883), .DIN2(n8129), .Q(n8882) );
  nnd2s1 U8935 ( .DIN1(n7827), .DIN2(n8884), .Q(n8874) );
  nnd3s1 U8936 ( .DIN1(n8854), .DIN2(n8449), .DIN3(n7838), .Q(n8884) );
  nnd2s1 U8937 ( .DIN1(n8433), .DIN2(n8883), .Q(n8873) );
  nnd3s1 U8938 ( .DIN1(n8885), .DIN2(n8886), .DIN3(n8887), .Q(n8871) );
  nnd2s1 U8939 ( .DIN1(n8170), .DIN2(n8888), .Q(n8887) );
  nnd2s1 U8940 ( .DIN1(n7817), .DIN2(n7820), .Q(n8886) );
  nnd2s1 U8941 ( .DIN1(n7947), .DIN2(n7821), .Q(n8885) );
  nor2s1 U8942 ( .DIN1(n8817), .DIN2(n7966), .Q(n8870) );
  nor2s1 U8943 ( .DIN1(n8475), .DIN2(n8825), .Q(n8869) );
  nor4s1 U8944 ( .DIN1(n8889), .DIN2(n8890), .DIN3(n8891), .DIN4(n8892), 
        .Q(n8125) );
  nnd4s1 U8945 ( .DIN1(n8893), .DIN2(n8894), .DIN3(n8895), .DIN4(n8896), 
        .Q(n8892) );
  nnd2s1 U8946 ( .DIN1(n7818), .DIN2(n7839), .Q(n8896) );
  nnd2s1 U8947 ( .DIN1(n7963), .DIN2(n8139), .Q(n8895) );
  nnd2s1 U8948 ( .DIN1(n8160), .DIN2(n7827), .Q(n8894) );
  nnd2s1 U8949 ( .DIN1(n8128), .DIN2(n8130), .Q(n8893) );
  nnd3s1 U8950 ( .DIN1(n8897), .DIN2(n8898), .DIN3(n8899), .Q(n8891) );
  nnd2s1 U8951 ( .DIN1(n7811), .DIN2(n8900), .Q(n8899) );
  nnd3s1 U8952 ( .DIN1(n8149), .DIN2(n8419), .DIN3(n7966), .Q(n8900) );
  nnd2s1 U8953 ( .DIN1(n8163), .DIN2(n8901), .Q(n8898) );
  nnd2s1 U8954 ( .DIN1(n8843), .DIN2(n8149), .Q(n8901) );
  nor2s1 U8955 ( .DIN1(n8888), .DIN2(n8883), .Q(n8843) );
  nnd2s1 U8956 ( .DIN1(n8432), .DIN2(n8902), .Q(n8897) );
  nnd2s1 U8957 ( .DIN1(n8818), .DIN2(n8475), .Q(n8902) );
  nor2s1 U8958 ( .DIN1(n8422), .DIN2(n8453), .Q(n8890) );
  nor2s1 U8959 ( .DIN1(n8155), .DIN2(n8450), .Q(n8889) );
  hi1s1 U8960 ( .DIN(n7840), .Q(n8155) );
  nor2s1 U8961 ( .DIN1(n8903), .DIN2(n8904), .Q(n8427) );
  nnd4s1 U8962 ( .DIN1(n8905), .DIN2(n8906), .DIN3(n8907), .DIN4(n8908), 
        .Q(n8904) );
  nnd2s1 U8963 ( .DIN1(n7818), .DIN2(n8909), .Q(n8908) );
  nnd3s1 U8964 ( .DIN1(n8450), .DIN2(n8817), .DIN3(n8854), .Q(n8909) );
  nnd2s1 U8965 ( .DIN1(n7817), .DIN2(n8129), .Q(n8906) );
  nnd4s1 U8966 ( .DIN1(n8910), .DIN2(n8911), .DIN3(n8912), .DIN4(n8913), 
        .Q(n8903) );
  nnd2s1 U8967 ( .DIN1(n7839), .DIN2(n8914), .Q(n8913) );
  nnd2s1 U8968 ( .DIN1(n8915), .DIN2(n7966), .Q(n8914) );
  nnd2s1 U8969 ( .DIN1(n7810), .DIN2(n8916), .Q(n8912) );
  nnd2s1 U8970 ( .DIN1(n7835), .DIN2(n8917), .Q(n8911) );
  nnd2s1 U8971 ( .DIN1(n8453), .DIN2(n8854), .Q(n8917) );
  nnd2s1 U8972 ( .DIN1(n8432), .DIN2(n8918), .Q(n8910) );
  nnd2s1 U8973 ( .DIN1(n7953), .DIN2(n8449), .Q(n8918) );
  nnd3s1 U8974 ( .DIN1(n8919), .DIN2(n8920), .DIN3(n8921), .Q(n8863) );
  nnd2s1 U8975 ( .DIN1(n7819), .DIN2(n7827), .Q(n8921) );
  nnd2s1 U8976 ( .DIN1(n8883), .DIN2(n8922), .Q(n8920) );
  nnd3s1 U8977 ( .DIN1(n7838), .DIN2(n8817), .DIN3(n8923), .Q(n8922) );
  or2s1 U8978 ( .DIN1(n8149), .DIN2(n8924), .Q(n8919) );
  nnd3s1 U8979 ( .DIN1(n8925), .DIN2(n8926), .DIN3(n8927), .Q(n8862) );
  nnd2s1 U8980 ( .DIN1(n7835), .DIN2(n8928), .Q(n8927) );
  nnd2s1 U8981 ( .DIN1(n8457), .DIN2(n8452), .Q(n8928) );
  nnd2s1 U8982 ( .DIN1(n8147), .DIN2(n8929), .Q(n8926) );
  or2s1 U8983 ( .DIN1(n8174), .DIN2(n7820), .Q(n8929) );
  nnd2s1 U8984 ( .DIN1(n7966), .DIN2(n7952), .Q(n8174) );
  nnd2s1 U8985 ( .DIN1(n8170), .DIN2(n8930), .Q(n8925) );
  nnd2s1 U8986 ( .DIN1(n7833), .DIN2(n8137), .Q(n8930) );
  nnd2s1 U8987 ( .DIN1(n7963), .DIN2(n7948), .Q(n8805) );
  nnd2s1 U8988 ( .DIN1(n8128), .DIN2(n7831), .Q(n8804) );
  nnd3s1 U8989 ( .DIN1(n8931), .DIN2(n8932), .DIN3(n8933), .Q(n8802) );
  nnd2s1 U8990 ( .DIN1(n8888), .DIN2(n7839), .Q(n8933) );
  nnd2s1 U8991 ( .DIN1(n8409), .DIN2(n8934), .Q(n8932) );
  nnd4s1 U8992 ( .DIN1(n8935), .DIN2(n8936), .DIN3(n8937), .DIN4(n8938), 
        .Q(n8801) );
  nnd2s1 U8993 ( .DIN1(n8163), .DIN2(n8939), .Q(n8938) );
  nnd2s1 U8994 ( .DIN1(n7968), .DIN2(n8169), .Q(n8939) );
  nor2s1 U8995 ( .DIN1(n8129), .DIN2(n8139), .Q(n7968) );
  nnd2s1 U8996 ( .DIN1(n8139), .DIN2(n8940), .Q(n8937) );
  nnd2s1 U8997 ( .DIN1(n8151), .DIN2(n8452), .Q(n8940) );
  nnd2s1 U8998 ( .DIN1(n7812), .DIN2(n8941), .Q(n8936) );
  nnd2s1 U8999 ( .DIN1(n8152), .DIN2(n7838), .Q(n8941) );
  nnd2s1 U9000 ( .DIN1(n7827), .DIN2(n8441), .Q(n8935) );
  or3s1 U9001 ( .DIN1(n8942), .DIN2(n8943), .DIN3(n8944), .Q(n5705) );
  nnd4s1 U9002 ( .DIN1(n8945), .DIN2(n8946), .DIN3(n7976), .DIN4(n8947), 
        .Q(n8944) );
  and3s1 U9003 ( .DIN1(n8179), .DIN2(n8512), .DIN3(n8479), .Q(n8947) );
  nor4s1 U9004 ( .DIN1(n8948), .DIN2(n8949), .DIN3(n8950), .DIN4(n8951), 
        .Q(n8479) );
  nnd4s1 U9005 ( .DIN1(n8952), .DIN2(n8953), .DIN3(n8954), .DIN4(n8955), 
        .Q(n8951) );
  nnd2s1 U9006 ( .DIN1(n8198), .DIN2(n8001), .Q(n8955) );
  nor2s1 U9007 ( .DIN1(n8956), .DIN2(n8957), .Q(n8954) );
  nor2s1 U9008 ( .DIN1(n8000), .DIN2(n8958), .Q(n8957) );
  nor2s1 U9009 ( .DIN1(n8959), .DIN2(n8232), .Q(n8956) );
  nnd2s1 U9010 ( .DIN1(n8187), .DIN2(n8199), .Q(n8953) );
  nnd2s1 U9011 ( .DIN1(n8207), .DIN2(n7992), .Q(n8952) );
  nnd3s1 U9012 ( .DIN1(n8960), .DIN2(n8961), .DIN3(n8962), .Q(n8950) );
  nnd2s1 U9013 ( .DIN1(n8233), .DIN2(n8238), .Q(n8962) );
  nnd2s1 U9014 ( .DIN1(n8963), .DIN2(n8964), .Q(n8961) );
  nnd3s1 U9015 ( .DIN1(n8504), .DIN2(n8958), .DIN3(n8538), .Q(n8964) );
  nnd2s1 U9016 ( .DIN1(n8519), .DIN2(n8965), .Q(n8960) );
  nnd3s1 U9017 ( .DIN1(n8194), .DIN2(n7990), .DIN3(n7999), .Q(n8965) );
  nor2s1 U9018 ( .DIN1(n8194), .DIN2(n8540), .Q(n8949) );
  nor2s1 U9019 ( .DIN1(n8966), .DIN2(n8967), .Q(n8948) );
  nor4s1 U9020 ( .DIN1(n8968), .DIN2(n8969), .DIN3(n8970), .DIN4(n8971), 
        .Q(n8512) );
  nnd4s1 U9021 ( .DIN1(n8972), .DIN2(n8973), .DIN3(n8974), .DIN4(n8975), 
        .Q(n8971) );
  nor2s1 U9022 ( .DIN1(n8976), .DIN2(n8977), .Q(n8975) );
  nor2s1 U9023 ( .DIN1(n8958), .DIN2(n8967), .Q(n8977) );
  nor2s1 U9024 ( .DIN1(n8236), .DIN2(n7990), .Q(n8976) );
  nnd2s1 U9025 ( .DIN1(n7984), .DIN2(n8230), .Q(n8973) );
  nnd2s1 U9026 ( .DIN1(n8185), .DIN2(n7982), .Q(n8972) );
  nnd3s1 U9027 ( .DIN1(n8978), .DIN2(n8979), .DIN3(n8980), .Q(n8970) );
  nnd2s1 U9028 ( .DIN1(n8196), .DIN2(n8981), .Q(n8980) );
  nnd2s1 U9029 ( .DIN1(n8539), .DIN2(n8212), .Q(n8981) );
  nnd2s1 U9030 ( .DIN1(n7981), .DIN2(n8982), .Q(n8979) );
  nnd2s1 U9031 ( .DIN1(n8564), .DIN2(n8504), .Q(n8982) );
  nnd2s1 U9032 ( .DIN1(n8204), .DIN2(n8234), .Q(n8978) );
  nnd2s1 U9033 ( .DIN1(n8215), .DIN2(n8505), .Q(n8234) );
  nor2s1 U9034 ( .DIN1(n8983), .DIN2(n8004), .Q(n8969) );
  nor2s1 U9035 ( .DIN1(n7983), .DIN2(n8213), .Q(n8983) );
  nor2s1 U9036 ( .DIN1(n8984), .DIN2(n8536), .Q(n8968) );
  and2s1 U9037 ( .DIN1(n8194), .DIN2(n8985), .Q(n8984) );
  nor4s1 U9038 ( .DIN1(n8986), .DIN2(n8987), .DIN3(n8988), .DIN4(n8989), 
        .Q(n8179) );
  nnd4s1 U9039 ( .DIN1(n8990), .DIN2(n8991), .DIN3(n8992), .DIN4(n8993), 
        .Q(n8989) );
  nnd2s1 U9040 ( .DIN1(n8518), .DIN2(n8199), .Q(n8993) );
  nor2s1 U9041 ( .DIN1(n8994), .DIN2(n8995), .Q(n8992) );
  nor2s1 U9042 ( .DIN1(n8996), .DIN2(n8004), .Q(n8994) );
  nnd2s1 U9043 ( .DIN1(n8197), .DIN2(n8207), .Q(n8991) );
  nnd2s1 U9044 ( .DIN1(n8186), .DIN2(n8562), .Q(n8990) );
  nnd3s1 U9045 ( .DIN1(n8997), .DIN2(n8998), .DIN3(n8999), .Q(n8988) );
  nnd2s1 U9046 ( .DIN1(n7982), .DIN2(n9000), .Q(n8999) );
  nnd2s1 U9047 ( .DIN1(n7992), .DIN2(n9001), .Q(n8998) );
  nnd2s1 U9048 ( .DIN1(n8536), .DIN2(n8504), .Q(n9001) );
  nnd2s1 U9049 ( .DIN1(n8519), .DIN2(n9002), .Q(n8997) );
  nnd3s1 U9050 ( .DIN1(n8508), .DIN2(n8967), .DIN3(n9003), .Q(n9002) );
  nor2s1 U9051 ( .DIN1(n7990), .DIN2(n8540), .Q(n8987) );
  nor2s1 U9052 ( .DIN1(n8007), .DIN2(n8237), .Q(n8986) );
  nor3s1 U9053 ( .DIN1(n9004), .DIN2(n9005), .DIN3(n9006), .Q(n7976) );
  nnd4s1 U9054 ( .DIN1(n8513), .DIN2(n8181), .DIN3(n8483), .DIN4(n9007), 
        .Q(n9006) );
  and3s1 U9055 ( .DIN1(n9008), .DIN2(n9009), .DIN3(n9010), .Q(n9007) );
  nnd2s1 U9056 ( .DIN1(n8186), .DIN2(n8494), .Q(n9010) );
  nnd2s1 U9057 ( .DIN1(n8224), .DIN2(n8001), .Q(n9008) );
  nor4s1 U9058 ( .DIN1(n9011), .DIN2(n9012), .DIN3(n9013), .DIN4(n9014), 
        .Q(n8483) );
  nnd4s1 U9059 ( .DIN1(n9015), .DIN2(n9016), .DIN3(n9017), .DIN4(n9018), 
        .Q(n9014) );
  nnd2s1 U9060 ( .DIN1(n8186), .DIN2(n9019), .Q(n9018) );
  nnd2s1 U9061 ( .DIN1(n9020), .DIN2(n8508), .Q(n9019) );
  nor2s1 U9062 ( .DIN1(n9021), .DIN2(n9022), .Q(n9017) );
  nor2s1 U9063 ( .DIN1(n9023), .DIN2(n8236), .Q(n9022) );
  nor2s1 U9064 ( .DIN1(n8224), .DIN2(n8009), .Q(n9023) );
  nor2s1 U9065 ( .DIN1(n9024), .DIN2(n9025), .Q(n9021) );
  nor2s1 U9066 ( .DIN1(n9026), .DIN2(n8185), .Q(n9024) );
  nnd2s1 U9067 ( .DIN1(n8562), .DIN2(n9027), .Q(n9016) );
  nnd3s1 U9068 ( .DIN1(n8996), .DIN2(n8535), .DIN3(n8540), .Q(n9027) );
  nnd2s1 U9069 ( .DIN1(n8519), .DIN2(n9026), .Q(n9015) );
  nnd3s1 U9070 ( .DIN1(n9028), .DIN2(n9029), .DIN3(n9030), .Q(n9013) );
  nnd2s1 U9071 ( .DIN1(n8233), .DIN2(n9031), .Q(n9030) );
  nnd2s1 U9072 ( .DIN1(n8492), .DIN2(n8963), .Q(n9029) );
  nnd2s1 U9073 ( .DIN1(n7981), .DIN2(n8204), .Q(n9028) );
  nor2s1 U9074 ( .DIN1(n8958), .DIN2(n8004), .Q(n9012) );
  nor2s1 U9075 ( .DIN1(n8564), .DIN2(n8967), .Q(n9011) );
  nor4s1 U9076 ( .DIN1(n9032), .DIN2(n9033), .DIN3(n9034), .DIN4(n9035), 
        .Q(n8181) );
  nnd4s1 U9077 ( .DIN1(n9036), .DIN2(n9037), .DIN3(n9038), .DIN4(n9039), 
        .Q(n9035) );
  nnd2s1 U9078 ( .DIN1(n8494), .DIN2(n8230), .Q(n9039) );
  nnd2s1 U9079 ( .DIN1(n8001), .DIN2(n8196), .Q(n9038) );
  nnd2s1 U9080 ( .DIN1(n8221), .DIN2(n8562), .Q(n9037) );
  nnd2s1 U9081 ( .DIN1(n8197), .DIN2(n8186), .Q(n9036) );
  nnd3s1 U9082 ( .DIN1(n9040), .DIN2(n9041), .DIN3(n9042), .Q(n9034) );
  nnd2s1 U9083 ( .DIN1(n8005), .DIN2(n9043), .Q(n9042) );
  nnd3s1 U9084 ( .DIN1(n8209), .DIN2(n8505), .DIN3(n8004), .Q(n9043) );
  nnd2s1 U9085 ( .DIN1(n8225), .DIN2(n9044), .Q(n9041) );
  nnd2s1 U9086 ( .DIN1(n8985), .DIN2(n8209), .Q(n9044) );
  nor2s1 U9087 ( .DIN1(n9031), .DIN2(n9026), .Q(n8985) );
  nnd2s1 U9088 ( .DIN1(n8518), .DIN2(n9045), .Q(n9040) );
  nnd2s1 U9089 ( .DIN1(n8959), .DIN2(n8564), .Q(n9045) );
  nor2s1 U9090 ( .DIN1(n8508), .DIN2(n8539), .Q(n9033) );
  nor2s1 U9091 ( .DIN1(n8216), .DIN2(n8536), .Q(n9032) );
  hi1s1 U9092 ( .DIN(n9046), .Q(n8216) );
  nor2s1 U9093 ( .DIN1(n9047), .DIN2(n9048), .Q(n8513) );
  nnd4s1 U9094 ( .DIN1(n9049), .DIN2(n9050), .DIN3(n9051), .DIN4(n9052), 
        .Q(n9048) );
  nnd2s1 U9095 ( .DIN1(n8494), .DIN2(n9053), .Q(n9052) );
  nnd3s1 U9096 ( .DIN1(n8536), .DIN2(n8958), .DIN3(n8996), .Q(n9053) );
  nnd2s1 U9097 ( .DIN1(n8492), .DIN2(n8185), .Q(n9050) );
  nnd4s1 U9098 ( .DIN1(n9054), .DIN2(n9055), .DIN3(n9056), .DIN4(n9057), 
        .Q(n9047) );
  nnd2s1 U9099 ( .DIN1(n8230), .DIN2(n9058), .Q(n9057) );
  nnd2s1 U9100 ( .DIN1(n9059), .DIN2(n8004), .Q(n9058) );
  nnd2s1 U9101 ( .DIN1(n7983), .DIN2(n9060), .Q(n9056) );
  nnd2s1 U9102 ( .DIN1(n7992), .DIN2(n9061), .Q(n9055) );
  nnd2s1 U9103 ( .DIN1(n8539), .DIN2(n8996), .Q(n9061) );
  nnd2s1 U9104 ( .DIN1(n8518), .DIN2(n9062), .Q(n9054) );
  nnd2s1 U9105 ( .DIN1(n7989), .DIN2(n8535), .Q(n9062) );
  nnd3s1 U9106 ( .DIN1(n9063), .DIN2(n9064), .DIN3(n9065), .Q(n9005) );
  nnd2s1 U9107 ( .DIN1(n7982), .DIN2(n8562), .Q(n9065) );
  nnd2s1 U9108 ( .DIN1(n9026), .DIN2(n9066), .Q(n9064) );
  nnd3s1 U9109 ( .DIN1(n8540), .DIN2(n8958), .DIN3(n9067), .Q(n9066) );
  or2s1 U9110 ( .DIN1(n8209), .DIN2(n9068), .Q(n9063) );
  nnd3s1 U9111 ( .DIN1(n9069), .DIN2(n9070), .DIN3(n9071), .Q(n9004) );
  nnd2s1 U9112 ( .DIN1(n7992), .DIN2(n9072), .Q(n9071) );
  nnd2s1 U9113 ( .DIN1(n8545), .DIN2(n8538), .Q(n9072) );
  nnd2s1 U9114 ( .DIN1(n8207), .DIN2(n9073), .Q(n9070) );
  or2s1 U9115 ( .DIN1(n8238), .DIN2(n8963), .Q(n9073) );
  nnd2s1 U9116 ( .DIN1(n8004), .DIN2(n7988), .Q(n8238) );
  nnd2s1 U9117 ( .DIN1(n8233), .DIN2(n9074), .Q(n9069) );
  nnd2s1 U9118 ( .DIN1(n8500), .DIN2(n8194), .Q(n9074) );
  nnd2s1 U9119 ( .DIN1(n8001), .DIN2(n7984), .Q(n8946) );
  nnd2s1 U9120 ( .DIN1(n8197), .DIN2(n8213), .Q(n8945) );
  nnd3s1 U9121 ( .DIN1(n9075), .DIN2(n9076), .DIN3(n9077), .Q(n8943) );
  nnd2s1 U9122 ( .DIN1(n9031), .DIN2(n8230), .Q(n9077) );
  nnd2s1 U9123 ( .DIN1(n8493), .DIN2(n9078), .Q(n9076) );
  nnd4s1 U9124 ( .DIN1(n9079), .DIN2(n9080), .DIN3(n9081), .DIN4(n9082), 
        .Q(n8942) );
  nnd2s1 U9125 ( .DIN1(n8225), .DIN2(n9083), .Q(n9082) );
  nnd2s1 U9126 ( .DIN1(n8007), .DIN2(n8232), .Q(n9083) );
  nor2s1 U9127 ( .DIN1(n8185), .DIN2(n8196), .Q(n8007) );
  nnd2s1 U9128 ( .DIN1(n8196), .DIN2(n9084), .Q(n9081) );
  nnd2s1 U9129 ( .DIN1(n8211), .DIN2(n8538), .Q(n9084) );
  nnd2s1 U9130 ( .DIN1(n8187), .DIN2(n9085), .Q(n9080) );
  nnd2s1 U9131 ( .DIN1(n8212), .DIN2(n8540), .Q(n9085) );
  nnd2s1 U9132 ( .DIN1(n8562), .DIN2(n8527), .Q(n9079) );
  xor2s1 U9133 ( .DIN1(n5056), .DIN2(n9086), .Q(n8796) );
  xor2s1 U9134 ( .DIN1(n1505), .DIN2(n5032), .Q(n9086) );
  or3s1 U9135 ( .DIN1(n9087), .DIN2(n9088), .DIN3(n9089), .Q(n5032) );
  nnd4s1 U9136 ( .DIN1(n9090), .DIN2(n9091), .DIN3(n9092), .DIN4(n9093), 
        .Q(n9089) );
  and3s1 U9137 ( .DIN1(n9094), .DIN2(n9095), .DIN3(n9096), .Q(n9093) );
  nnd2s1 U9138 ( .DIN1(n8030), .DIN2(n8037), .Q(n9095) );
  nnd2s1 U9139 ( .DIN1(n8023), .DIN2(n7853), .Q(n9094) );
  nnd3s1 U9140 ( .DIN1(n9097), .DIN2(n9098), .DIN3(n9099), .Q(n9088) );
  nnd2s1 U9141 ( .DIN1(n8257), .DIN2(n8021), .Q(n9099) );
  or2s1 U9142 ( .DIN1(n8281), .DIN2(n9100), .Q(n9098) );
  nnd2s1 U9143 ( .DIN1(n8310), .DIN2(n8072), .Q(n9097) );
  nnd4s1 U9144 ( .DIN1(n9101), .DIN2(n9102), .DIN3(n9103), .DIN4(n9104), 
        .Q(n9087) );
  nnd2s1 U9145 ( .DIN1(n8649), .DIN2(n9105), .Q(n9104) );
  nnd2s1 U9146 ( .DIN1(n8689), .DIN2(n8252), .Q(n9105) );
  nnd2s1 U9147 ( .DIN1(n8036), .DIN2(n9106), .Q(n9103) );
  nnd2s1 U9148 ( .DIN1(n8283), .DIN2(n7868), .Q(n9106) );
  nor2s1 U9149 ( .DIN1(n8272), .DIN2(n8271), .Q(n8283) );
  nnd2s1 U9150 ( .DIN1(n8064), .DIN2(n9107), .Q(n9102) );
  nnd2s1 U9151 ( .DIN1(n8076), .DIN2(n8253), .Q(n9107) );
  nnd2s1 U9152 ( .DIN1(n7870), .DIN2(n9108), .Q(n9101) );
  or3s1 U9153 ( .DIN1(n9109), .DIN2(n9110), .DIN3(n9111), .Q(n5056) );
  nnd4s1 U9154 ( .DIN1(n9112), .DIN2(n9113), .DIN3(n8085), .DIN4(n9114), 
        .Q(n9111) );
  and3s1 U9155 ( .DIN1(n8333), .DIN2(n8741), .DIN3(n8711), .Q(n9114) );
  nor4s1 U9156 ( .DIN1(n9115), .DIN2(n9116), .DIN3(n9117), .DIN4(n9118), 
        .Q(n8711) );
  nnd4s1 U9157 ( .DIN1(n9119), .DIN2(n9120), .DIN3(n9121), .DIN4(n9122), 
        .Q(n9118) );
  nnd2s1 U9158 ( .DIN1(n7903), .DIN2(n8106), .Q(n9122) );
  nor2s1 U9159 ( .DIN1(n9123), .DIN2(n9124), .Q(n9121) );
  nor2s1 U9160 ( .DIN1(n8105), .DIN2(n9125), .Q(n9124) );
  nor2s1 U9161 ( .DIN1(n9126), .DIN2(n8379), .Q(n9123) );
  nnd2s1 U9162 ( .DIN1(n7893), .DIN2(n8350), .Q(n9120) );
  nnd2s1 U9163 ( .DIN1(n8357), .DIN2(n7916), .Q(n9119) );
  nnd3s1 U9164 ( .DIN1(n9127), .DIN2(n9128), .DIN3(n9129), .Q(n9117) );
  nnd2s1 U9165 ( .DIN1(n8380), .DIN2(n8384), .Q(n9129) );
  nnd2s1 U9166 ( .DIN1(n7901), .DIN2(n9130), .Q(n9128) );
  nnd3s1 U9167 ( .DIN1(n8733), .DIN2(n9125), .DIN3(n8767), .Q(n9130) );
  nnd2s1 U9168 ( .DIN1(n8748), .DIN2(n9131), .Q(n9127) );
  nnd3s1 U9169 ( .DIN1(n8347), .DIN2(n7915), .DIN3(n8104), .Q(n9131) );
  nor2s1 U9170 ( .DIN1(n8347), .DIN2(n7919), .Q(n9116) );
  nor2s1 U9171 ( .DIN1(n9132), .DIN2(n9133), .Q(n9115) );
  nor4s1 U9172 ( .DIN1(n9134), .DIN2(n9135), .DIN3(n9136), .DIN4(n9137), 
        .Q(n8741) );
  nnd4s1 U9173 ( .DIN1(n9138), .DIN2(n9139), .DIN3(n9140), .DIN4(n9141), 
        .Q(n9137) );
  nor2s1 U9174 ( .DIN1(n9142), .DIN2(n9143), .Q(n9141) );
  nor2s1 U9175 ( .DIN1(n9125), .DIN2(n9133), .Q(n9143) );
  nor2s1 U9176 ( .DIN1(n8383), .DIN2(n7915), .Q(n9142) );
  nnd2s1 U9177 ( .DIN1(n8091), .DIN2(n7920), .Q(n9139) );
  nnd2s1 U9178 ( .DIN1(n8339), .DIN2(n7900), .Q(n9138) );
  nnd3s1 U9179 ( .DIN1(n9144), .DIN2(n9145), .DIN3(n9146), .Q(n9136) );
  nnd2s1 U9180 ( .DIN1(n8349), .DIN2(n9147), .Q(n9146) );
  nnd2s1 U9181 ( .DIN1(n8768), .DIN2(n8362), .Q(n9147) );
  nnd2s1 U9182 ( .DIN1(n8090), .DIN2(n9148), .Q(n9145) );
  nnd2s1 U9183 ( .DIN1(n8790), .DIN2(n8733), .Q(n9148) );
  nnd2s1 U9184 ( .DIN1(n7902), .DIN2(n8381), .Q(n9144) );
  nnd2s1 U9185 ( .DIN1(n8364), .DIN2(n8734), .Q(n8381) );
  nor2s1 U9186 ( .DIN1(n9149), .DIN2(n8109), .Q(n9135) );
  nor2s1 U9187 ( .DIN1(n7891), .DIN2(n7912), .Q(n9149) );
  nor2s1 U9188 ( .DIN1(n9150), .DIN2(n8765), .Q(n9134) );
  and2s1 U9189 ( .DIN1(n8347), .DIN2(n9151), .Q(n9150) );
  nor4s1 U9190 ( .DIN1(n9152), .DIN2(n9153), .DIN3(n9154), .DIN4(n9155), 
        .Q(n8333) );
  nnd4s1 U9191 ( .DIN1(n9156), .DIN2(n9157), .DIN3(n9158), .DIN4(n9159), 
        .Q(n9155) );
  nnd2s1 U9192 ( .DIN1(n8747), .DIN2(n8350), .Q(n9159) );
  nor2s1 U9193 ( .DIN1(n9160), .DIN2(n9161), .Q(n9158) );
  nor2s1 U9194 ( .DIN1(n9162), .DIN2(n8109), .Q(n9160) );
  nnd2s1 U9195 ( .DIN1(n8338), .DIN2(n8357), .Q(n9157) );
  nnd2s1 U9196 ( .DIN1(n8340), .DIN2(n7908), .Q(n9156) );
  nnd3s1 U9197 ( .DIN1(n9163), .DIN2(n9164), .DIN3(n9165), .Q(n9154) );
  nnd2s1 U9198 ( .DIN1(n7900), .DIN2(n9166), .Q(n9165) );
  nnd2s1 U9199 ( .DIN1(n7916), .DIN2(n9167), .Q(n9164) );
  nnd2s1 U9200 ( .DIN1(n8765), .DIN2(n8733), .Q(n9167) );
  nnd2s1 U9201 ( .DIN1(n8748), .DIN2(n9168), .Q(n9163) );
  nnd3s1 U9202 ( .DIN1(n8737), .DIN2(n9133), .DIN3(n9169), .Q(n9168) );
  nor2s1 U9203 ( .DIN1(n7915), .DIN2(n7919), .Q(n9153) );
  nor2s1 U9204 ( .DIN1(n8111), .DIN2(n7911), .Q(n9152) );
  nor3s1 U9205 ( .DIN1(n9170), .DIN2(n9171), .DIN3(n9172), .Q(n8085) );
  nnd4s1 U9206 ( .DIN1(n8742), .DIN2(n8335), .DIN3(n8715), .DIN4(n9173), 
        .Q(n9172) );
  and3s1 U9207 ( .DIN1(n9174), .DIN2(n9175), .DIN3(n9176), .Q(n9173) );
  nnd2s1 U9208 ( .DIN1(n8340), .DIN2(n7899), .Q(n9176) );
  nnd2s1 U9209 ( .DIN1(n7890), .DIN2(n8106), .Q(n9174) );
  nor4s1 U9210 ( .DIN1(n9177), .DIN2(n9178), .DIN3(n9179), .DIN4(n9180), 
        .Q(n8715) );
  nnd4s1 U9211 ( .DIN1(n9181), .DIN2(n9182), .DIN3(n9183), .DIN4(n9184), 
        .Q(n9180) );
  nnd2s1 U9212 ( .DIN1(n8340), .DIN2(n9185), .Q(n9184) );
  nnd2s1 U9213 ( .DIN1(n9186), .DIN2(n8737), .Q(n9185) );
  nor2s1 U9214 ( .DIN1(n9187), .DIN2(n9188), .Q(n9183) );
  nor2s1 U9215 ( .DIN1(n9189), .DIN2(n8383), .Q(n9188) );
  nor2s1 U9216 ( .DIN1(n7890), .DIN2(n8113), .Q(n9189) );
  nor2s1 U9217 ( .DIN1(n9190), .DIN2(n7918), .Q(n9187) );
  nor2s1 U9218 ( .DIN1(n9191), .DIN2(n8339), .Q(n9190) );
  nnd2s1 U9219 ( .DIN1(n7908), .DIN2(n9192), .Q(n9182) );
  nnd3s1 U9220 ( .DIN1(n9162), .DIN2(n8764), .DIN3(n7919), .Q(n9192) );
  nnd2s1 U9221 ( .DIN1(n8748), .DIN2(n9191), .Q(n9181) );
  nnd3s1 U9222 ( .DIN1(n9193), .DIN2(n9194), .DIN3(n9195), .Q(n9179) );
  nnd2s1 U9223 ( .DIN1(n8380), .DIN2(n9196), .Q(n9195) );
  nnd2s1 U9224 ( .DIN1(n7898), .DIN2(n7901), .Q(n9194) );
  nnd2s1 U9225 ( .DIN1(n8090), .DIN2(n7902), .Q(n9193) );
  nor2s1 U9226 ( .DIN1(n9125), .DIN2(n8109), .Q(n9178) );
  nor2s1 U9227 ( .DIN1(n8790), .DIN2(n9133), .Q(n9177) );
  nor4s1 U9228 ( .DIN1(n9197), .DIN2(n9198), .DIN3(n9199), .DIN4(n9200), 
        .Q(n8335) );
  nnd4s1 U9229 ( .DIN1(n9201), .DIN2(n9202), .DIN3(n9203), .DIN4(n9204), 
        .Q(n9200) );
  nnd2s1 U9230 ( .DIN1(n7899), .DIN2(n7920), .Q(n9204) );
  nnd2s1 U9231 ( .DIN1(n8106), .DIN2(n8349), .Q(n9203) );
  nnd2s1 U9232 ( .DIN1(n8370), .DIN2(n7908), .Q(n9202) );
  nnd2s1 U9233 ( .DIN1(n8338), .DIN2(n8340), .Q(n9201) );
  nnd3s1 U9234 ( .DIN1(n9205), .DIN2(n9206), .DIN3(n9207), .Q(n9199) );
  nnd2s1 U9235 ( .DIN1(n7892), .DIN2(n9208), .Q(n9207) );
  nnd3s1 U9236 ( .DIN1(n8359), .DIN2(n8734), .DIN3(n8109), .Q(n9208) );
  nnd2s1 U9237 ( .DIN1(n8373), .DIN2(n9209), .Q(n9206) );
  nnd2s1 U9238 ( .DIN1(n9151), .DIN2(n8359), .Q(n9209) );
  nor2s1 U9239 ( .DIN1(n9196), .DIN2(n9191), .Q(n9151) );
  nnd2s1 U9240 ( .DIN1(n8747), .DIN2(n9210), .Q(n9205) );
  nnd2s1 U9241 ( .DIN1(n9126), .DIN2(n8790), .Q(n9210) );
  nor2s1 U9242 ( .DIN1(n8737), .DIN2(n8768), .Q(n9198) );
  nor2s1 U9243 ( .DIN1(n8365), .DIN2(n8765), .Q(n9197) );
  hi1s1 U9244 ( .DIN(n7921), .Q(n8365) );
  nor2s1 U9245 ( .DIN1(n9211), .DIN2(n9212), .Q(n8742) );
  nnd4s1 U9246 ( .DIN1(n9213), .DIN2(n9214), .DIN3(n9215), .DIN4(n9216), 
        .Q(n9212) );
  nnd2s1 U9247 ( .DIN1(n7899), .DIN2(n9217), .Q(n9216) );
  nnd3s1 U9248 ( .DIN1(n8765), .DIN2(n9125), .DIN3(n9162), .Q(n9217) );
  nnd2s1 U9249 ( .DIN1(n7898), .DIN2(n8339), .Q(n9214) );
  nnd4s1 U9250 ( .DIN1(n9218), .DIN2(n9219), .DIN3(n9220), .DIN4(n9221), 
        .Q(n9211) );
  nnd2s1 U9251 ( .DIN1(n7920), .DIN2(n9222), .Q(n9221) );
  nnd2s1 U9252 ( .DIN1(n9223), .DIN2(n8109), .Q(n9222) );
  nnd2s1 U9253 ( .DIN1(n7891), .DIN2(n9224), .Q(n9220) );
  nnd2s1 U9254 ( .DIN1(n7916), .DIN2(n9225), .Q(n9219) );
  nnd2s1 U9255 ( .DIN1(n8768), .DIN2(n9162), .Q(n9225) );
  nnd2s1 U9256 ( .DIN1(n8747), .DIN2(n9226), .Q(n9218) );
  nnd2s1 U9257 ( .DIN1(n8096), .DIN2(n8764), .Q(n9226) );
  nnd3s1 U9258 ( .DIN1(n9227), .DIN2(n9228), .DIN3(n9229), .Q(n9171) );
  nnd2s1 U9259 ( .DIN1(n7900), .DIN2(n7908), .Q(n9229) );
  nnd2s1 U9260 ( .DIN1(n9191), .DIN2(n9230), .Q(n9228) );
  nnd3s1 U9261 ( .DIN1(n7919), .DIN2(n9125), .DIN3(n9231), .Q(n9230) );
  or2s1 U9262 ( .DIN1(n8359), .DIN2(n9232), .Q(n9227) );
  nnd3s1 U9263 ( .DIN1(n9233), .DIN2(n9234), .DIN3(n9235), .Q(n9170) );
  nnd2s1 U9264 ( .DIN1(n7916), .DIN2(n9236), .Q(n9235) );
  nnd2s1 U9265 ( .DIN1(n8772), .DIN2(n8767), .Q(n9236) );
  nnd2s1 U9266 ( .DIN1(n8357), .DIN2(n9237), .Q(n9234) );
  or2s1 U9267 ( .DIN1(n8384), .DIN2(n7901), .Q(n9237) );
  nnd2s1 U9268 ( .DIN1(n8109), .DIN2(n8095), .Q(n8384) );
  nnd2s1 U9269 ( .DIN1(n8380), .DIN2(n9238), .Q(n9233) );
  nnd2s1 U9270 ( .DIN1(n7914), .DIN2(n8347), .Q(n9238) );
  nnd2s1 U9271 ( .DIN1(n8106), .DIN2(n8091), .Q(n9113) );
  nnd2s1 U9272 ( .DIN1(n8338), .DIN2(n7912), .Q(n9112) );
  nnd3s1 U9273 ( .DIN1(n9239), .DIN2(n9240), .DIN3(n9241), .Q(n9110) );
  nnd2s1 U9274 ( .DIN1(n9196), .DIN2(n7920), .Q(n9241) );
  nnd2s1 U9275 ( .DIN1(n8724), .DIN2(n9242), .Q(n9240) );
  nnd4s1 U9276 ( .DIN1(n9243), .DIN2(n9244), .DIN3(n9245), .DIN4(n9246), 
        .Q(n9109) );
  nnd2s1 U9277 ( .DIN1(n8373), .DIN2(n9247), .Q(n9246) );
  nnd2s1 U9278 ( .DIN1(n8111), .DIN2(n8379), .Q(n9247) );
  nor2s1 U9279 ( .DIN1(n8339), .DIN2(n8349), .Q(n8111) );
  nnd2s1 U9280 ( .DIN1(n8349), .DIN2(n9248), .Q(n9245) );
  nnd2s1 U9281 ( .DIN1(n8361), .DIN2(n8767), .Q(n9248) );
  nnd2s1 U9282 ( .DIN1(n7893), .DIN2(n9249), .Q(n9244) );
  nnd2s1 U9283 ( .DIN1(n8362), .DIN2(n7919), .Q(n9249) );
  nnd2s1 U9284 ( .DIN1(n7908), .DIN2(n8756), .Q(n9243) );
  nnd2s1 U9285 ( .DIN1(n9250), .DIN2(n1603), .Q(n8793) );
  xor2s1 U9286 ( .DIN1(w0[3]), .DIN2(text_in_r[99]), .Q(n9250) );
  nnd3s1 U9287 ( .DIN1(n9251), .DIN2(n9252), .DIN3(n9253), .Q(N228) );
  nnd2s1 U9288 ( .DIN1(n1597), .DIN2(n9254), .Q(n9253) );
  xor2s1 U9289 ( .DIN1(w0[2]), .DIN2(text_in_r[98]), .Q(n9254) );
  nnd2s1 U9290 ( .DIN1(n9255), .DIN2(n5703), .Q(n9252) );
  nnd2s1 U9291 ( .DIN1(n9256), .DIN2(n9257), .Q(n9255) );
  nnd2s1 U9292 ( .DIN1(n7605), .DIN2(n9258), .Q(n9257) );
  nnd2s1 U9293 ( .DIN1(n9259), .DIN2(n7607), .Q(n9256) );
  nnd2s1 U9294 ( .DIN1(n9260), .DIN2(n9261), .Q(n9251) );
  nnd2s1 U9295 ( .DIN1(n9262), .DIN2(n9263), .Q(n9261) );
  nnd2s1 U9296 ( .DIN1(n7607), .DIN2(n9258), .Q(n9263) );
  nor2s1 U9297 ( .DIN1(n7771), .DIN2(n1596), .Q(n7607) );
  nnd2s1 U9298 ( .DIN1(n9259), .DIN2(n7605), .Q(n9262) );
  nor2s1 U9299 ( .DIN1(n9264), .DIN2(n1594), .Q(n7605) );
  hi1s1 U9300 ( .DIN(n7771), .Q(n9264) );
  xor2s1 U9301 ( .DIN1(n5704), .DIN2(n5079), .Q(n7771) );
  hi1s1 U9302 ( .DIN(n7621), .Q(n5079) );
  or3s1 U9303 ( .DIN1(n9265), .DIN2(n9266), .DIN3(n9267), .Q(n7621) );
  nnd4s1 U9304 ( .DIN1(n9268), .DIN2(n9269), .DIN3(n7803), .DIN4(n9270), 
        .Q(n9267) );
  and3s1 U9305 ( .DIN1(n9271), .DIN2(n9272), .DIN3(n9273), .Q(n9270) );
  nnd2s1 U9306 ( .DIN1(n7831), .DIN2(n7822), .Q(n9272) );
  nnd2s1 U9307 ( .DIN1(n7827), .DIN2(n8140), .Q(n9271) );
  nor3s1 U9308 ( .DIN1(n9274), .DIN2(n9275), .DIN3(n9276), .Q(n7803) );
  nnd4s1 U9309 ( .DIN1(n9277), .DIN2(n9278), .DIN3(n9279), .DIN4(n9280), 
        .Q(n9276) );
  and3s1 U9310 ( .DIN1(n9281), .DIN2(n9282), .DIN3(n9283), .Q(n9280) );
  nnd2s1 U9311 ( .DIN1(n7959), .DIN2(n7812), .Q(n9283) );
  nnd2s1 U9312 ( .DIN1(n8128), .DIN2(n7817), .Q(n9282) );
  nnd2s1 U9313 ( .DIN1(n7831), .DIN2(n8139), .Q(n9281) );
  nnd3s1 U9314 ( .DIN1(n9284), .DIN2(n9285), .DIN3(n8907), .Q(n9275) );
  nnd2s1 U9315 ( .DIN1(n8130), .DIN2(n8883), .Q(n8907) );
  or2s1 U9316 ( .DIN1(n7837), .DIN2(n8915), .Q(n9285) );
  nor2s1 U9317 ( .DIN1(n7809), .DIN2(n7820), .Q(n8915) );
  nnd2s1 U9318 ( .DIN1(n8163), .DIN2(n7970), .Q(n9284) );
  nnd2s1 U9319 ( .DIN1(n8154), .DIN2(n7961), .Q(n7970) );
  nnd4s1 U9320 ( .DIN1(n9286), .DIN2(n9287), .DIN3(n9288), .DIN4(n9289), 
        .Q(n9274) );
  nnd2s1 U9321 ( .DIN1(n8409), .DIN2(n9290), .Q(n9289) );
  nnd2s1 U9322 ( .DIN1(n7811), .DIN2(n9291), .Q(n9288) );
  nnd2s1 U9323 ( .DIN1(n7961), .DIN2(n8169), .Q(n9291) );
  nnd2s1 U9324 ( .DIN1(n8129), .DIN2(n9292), .Q(n9287) );
  nnd2s1 U9325 ( .DIN1(n8152), .DIN2(n7830), .Q(n9292) );
  nnd2s1 U9326 ( .DIN1(n7835), .DIN2(n9293), .Q(n9286) );
  nnd2s1 U9327 ( .DIN1(n8923), .DIN2(n8817), .Q(n9293) );
  hi1s1 U9328 ( .DIN(n8162), .Q(n8923) );
  nnd2s1 U9329 ( .DIN1(n8449), .DIN2(n8173), .Q(n8162) );
  nnd3s1 U9330 ( .DIN1(n9294), .DIN2(n9295), .DIN3(n9296), .Q(n9266) );
  nnd2s1 U9331 ( .DIN1(n8128), .DIN2(n7819), .Q(n9296) );
  or2s1 U9332 ( .DIN1(n7833), .DIN2(n7829), .Q(n9295) );
  nor2s1 U9333 ( .DIN1(n7959), .DIN2(n7963), .Q(n7829) );
  nnd2s1 U9334 ( .DIN1(n8432), .DIN2(n7839), .Q(n9294) );
  nnd4s1 U9335 ( .DIN1(n9297), .DIN2(n9298), .DIN3(n9299), .DIN4(n9300), 
        .Q(n9265) );
  nnd2s1 U9336 ( .DIN1(n8888), .DIN2(n9301), .Q(n9300) );
  nnd2s1 U9337 ( .DIN1(n8924), .DIN2(n8449), .Q(n9301) );
  nnd2s1 U9338 ( .DIN1(n7810), .DIN2(n9302), .Q(n9299) );
  nnd2s1 U9339 ( .DIN1(n8416), .DIN2(n7962), .Q(n9302) );
  nor2s1 U9340 ( .DIN1(n7818), .DIN2(n8883), .Q(n8416) );
  nnd2s1 U9341 ( .DIN1(n7811), .DIN2(n9303), .Q(n9298) );
  nnd2s1 U9342 ( .DIN1(n7812), .DIN2(n9290), .Q(n9297) );
  nnd2s1 U9343 ( .DIN1(n8453), .DIN2(n7830), .Q(n9290) );
  or3s1 U9344 ( .DIN1(n9304), .DIN2(n9305), .DIN3(n9306), .Q(n5704) );
  nnd4s1 U9345 ( .DIN1(n9307), .DIN2(n9308), .DIN3(n9309), .DIN4(n9310), 
        .Q(n9306) );
  and3s1 U9346 ( .DIN1(n9311), .DIN2(n9312), .DIN3(n9313), .Q(n9310) );
  nnd2s1 U9347 ( .DIN1(n8213), .DIN2(n8198), .Q(n9312) );
  nnd2s1 U9348 ( .DIN1(n8562), .DIN2(n8199), .Q(n9311) );
  nnd3s1 U9349 ( .DIN1(n9314), .DIN2(n9315), .DIN3(n9316), .Q(n9305) );
  nnd2s1 U9350 ( .DIN1(n8197), .DIN2(n7982), .Q(n9316) );
  or2s1 U9351 ( .DIN1(n8500), .DIN2(n9317), .Q(n9315) );
  nnd2s1 U9352 ( .DIN1(n8518), .DIN2(n8230), .Q(n9314) );
  nnd4s1 U9353 ( .DIN1(n9318), .DIN2(n9319), .DIN3(n9320), .DIN4(n9321), 
        .Q(n9304) );
  nnd2s1 U9354 ( .DIN1(n9031), .DIN2(n9322), .Q(n9321) );
  nnd2s1 U9355 ( .DIN1(n9068), .DIN2(n8535), .Q(n9322) );
  nnd2s1 U9356 ( .DIN1(n7983), .DIN2(n9323), .Q(n9320) );
  nnd2s1 U9357 ( .DIN1(n8502), .DIN2(n8000), .Q(n9323) );
  nor2s1 U9358 ( .DIN1(n8494), .DIN2(n9026), .Q(n8502) );
  nnd2s1 U9359 ( .DIN1(n8005), .DIN2(n9324), .Q(n9319) );
  nnd2s1 U9360 ( .DIN1(n8187), .DIN2(n9325), .Q(n9318) );
  hi1s1 U9361 ( .DIN(n9258), .Q(n9259) );
  xor2s1 U9362 ( .DIN1(n5055), .DIN2(n9326), .Q(n9258) );
  xnr2s1 U9363 ( .DIN1(w0[2]), .DIN2(n5031), .Q(n9326) );
  or3s1 U9364 ( .DIN1(n9327), .DIN2(n9328), .DIN3(n9329), .Q(n5031) );
  nnd4s1 U9365 ( .DIN1(n8326), .DIN2(n9330), .DIN3(n9331), .DIN4(n9332), 
        .Q(n9329) );
  and4s1 U9366 ( .DIN1(n9333), .DIN2(n9334), .DIN3(n9335), .DIN4(n9336), 
        .Q(n9332) );
  nnd2s1 U9367 ( .DIN1(n7866), .DIN2(n9337), .Q(n9336) );
  nnd2s1 U9368 ( .DIN1(n8277), .DIN2(n7868), .Q(n9337) );
  nnd2s1 U9369 ( .DIN1(n8257), .DIN2(n9338), .Q(n9335) );
  nnd2s1 U9370 ( .DIN1(n8253), .DIN2(n8284), .Q(n9338) );
  nnd2s1 U9371 ( .DIN1(n8022), .DIN2(n9339), .Q(n9334) );
  nnd3s1 U9372 ( .DIN1(n8059), .DIN2(n8260), .DIN3(n7858), .Q(n9339) );
  nnd2s1 U9373 ( .DIN1(n7870), .DIN2(n9340), .Q(n9333) );
  nnd2s1 U9374 ( .DIN1(n8049), .DIN2(n8271), .Q(n9331) );
  nnd2s1 U9375 ( .DIN1(n8023), .DIN2(n8063), .Q(n9330) );
  nnd2s1 U9376 ( .DIN1(n8037), .DIN2(n8078), .Q(n8326) );
  nnd3s1 U9377 ( .DIN1(n9341), .DIN2(n9342), .DIN3(n9090), .Q(n9328) );
  nor4s1 U9378 ( .DIN1(n9343), .DIN2(n9344), .DIN3(n9345), .DIN4(n9346), 
        .Q(n9090) );
  nnd4s1 U9379 ( .DIN1(n9347), .DIN2(n9348), .DIN3(n8672), .DIN4(n9349), 
        .Q(n9346) );
  nnd2s1 U9380 ( .DIN1(n8078), .DIN2(n8667), .Q(n9349) );
  nnd2s1 U9381 ( .DIN1(n8052), .DIN2(n8649), .Q(n8672) );
  nnd2s1 U9382 ( .DIN1(n8064), .DIN2(n8063), .Q(n9348) );
  nnd2s1 U9383 ( .DIN1(n7866), .DIN2(n8699), .Q(n9347) );
  nnd3s1 U9384 ( .DIN1(n9350), .DIN2(n9351), .DIN3(n9352), .Q(n9345) );
  nnd2s1 U9385 ( .DIN1(n8254), .DIN2(n9353), .Q(n9352) );
  nnd2s1 U9386 ( .DIN1(n7868), .DIN2(n7878), .Q(n9353) );
  nnd2s1 U9387 ( .DIN1(n8034), .DIN2(n9354), .Q(n9351) );
  nnd2s1 U9388 ( .DIN1(n8277), .DIN2(n8281), .Q(n9354) );
  nnd2s1 U9389 ( .DIN1(n8042), .DIN2(n9355), .Q(n9350) );
  nnd2s1 U9390 ( .DIN1(n7858), .DIN2(n8590), .Q(n9355) );
  nor2s1 U9391 ( .DIN1(n8072), .DIN2(n8063), .Q(n7858) );
  nor2s1 U9392 ( .DIN1(n8582), .DIN2(n8054), .Q(n9344) );
  nor2s1 U9393 ( .DIN1(n8069), .DIN2(n8063), .Q(n8582) );
  nor2s1 U9394 ( .DIN1(n9356), .DIN2(n8032), .Q(n9343) );
  nor2s1 U9395 ( .DIN1(n8036), .DIN2(n7870), .Q(n9356) );
  nnd4s1 U9396 ( .DIN1(n9357), .DIN2(n9358), .DIN3(n9359), .DIN4(n9360), 
        .Q(n9327) );
  nnd2s1 U9397 ( .DIN1(n8699), .DIN2(n8036), .Q(n9360) );
  nnd2s1 U9398 ( .DIN1(n8316), .DIN2(n7861), .Q(n9359) );
  nnd2s1 U9399 ( .DIN1(n8052), .DIN2(n8272), .Q(n9358) );
  or3s1 U9400 ( .DIN1(n9361), .DIN2(n9362), .DIN3(n9363), .Q(n5055) );
  nnd4s1 U9401 ( .DIN1(n9364), .DIN2(n9365), .DIN3(n7884), .DIN4(n9366), 
        .Q(n9363) );
  and3s1 U9402 ( .DIN1(n9367), .DIN2(n9368), .DIN3(n9369), .Q(n9366) );
  nnd2s1 U9403 ( .DIN1(n7912), .DIN2(n7903), .Q(n9368) );
  nnd2s1 U9404 ( .DIN1(n7908), .DIN2(n8350), .Q(n9367) );
  nor3s1 U9405 ( .DIN1(n9370), .DIN2(n9371), .DIN3(n9372), .Q(n7884) );
  nnd4s1 U9406 ( .DIN1(n9373), .DIN2(n9374), .DIN3(n9375), .DIN4(n9376), 
        .Q(n9372) );
  and3s1 U9407 ( .DIN1(n9377), .DIN2(n9378), .DIN3(n9379), .Q(n9376) );
  nnd2s1 U9408 ( .DIN1(n8102), .DIN2(n7893), .Q(n9379) );
  nnd2s1 U9409 ( .DIN1(n8338), .DIN2(n7898), .Q(n9378) );
  nnd2s1 U9410 ( .DIN1(n7912), .DIN2(n8349), .Q(n9377) );
  nnd3s1 U9411 ( .DIN1(n9380), .DIN2(n9381), .DIN3(n9215), .Q(n9371) );
  nnd2s1 U9412 ( .DIN1(n8340), .DIN2(n9191), .Q(n9215) );
  or2s1 U9413 ( .DIN1(n7918), .DIN2(n9223), .Q(n9381) );
  nor2s1 U9414 ( .DIN1(n7890), .DIN2(n7901), .Q(n9223) );
  nnd2s1 U9415 ( .DIN1(n8373), .DIN2(n8113), .Q(n9380) );
  nnd2s1 U9416 ( .DIN1(n8364), .DIN2(n8104), .Q(n8113) );
  nnd4s1 U9417 ( .DIN1(n9382), .DIN2(n9383), .DIN3(n9384), .DIN4(n9385), 
        .Q(n9370) );
  nnd2s1 U9418 ( .DIN1(n8724), .DIN2(n9386), .Q(n9385) );
  nnd2s1 U9419 ( .DIN1(n7892), .DIN2(n9387), .Q(n9384) );
  nnd2s1 U9420 ( .DIN1(n8104), .DIN2(n8379), .Q(n9387) );
  nnd2s1 U9421 ( .DIN1(n8339), .DIN2(n9388), .Q(n9383) );
  nnd2s1 U9422 ( .DIN1(n8362), .DIN2(n7911), .Q(n9388) );
  nnd2s1 U9423 ( .DIN1(n7916), .DIN2(n9389), .Q(n9382) );
  nnd2s1 U9424 ( .DIN1(n9231), .DIN2(n9125), .Q(n9389) );
  hi1s1 U9425 ( .DIN(n8372), .Q(n9231) );
  nnd2s1 U9426 ( .DIN1(n8764), .DIN2(n8383), .Q(n8372) );
  nnd3s1 U9427 ( .DIN1(n9390), .DIN2(n9391), .DIN3(n9392), .Q(n9362) );
  nnd2s1 U9428 ( .DIN1(n8338), .DIN2(n7900), .Q(n9392) );
  or2s1 U9429 ( .DIN1(n7914), .DIN2(n7910), .Q(n9391) );
  nor2s1 U9430 ( .DIN1(n8102), .DIN2(n8106), .Q(n7910) );
  nnd2s1 U9431 ( .DIN1(n8747), .DIN2(n7920), .Q(n9390) );
  nnd4s1 U9432 ( .DIN1(n9393), .DIN2(n9394), .DIN3(n9395), .DIN4(n9396), 
        .Q(n9361) );
  nnd2s1 U9433 ( .DIN1(n9196), .DIN2(n9397), .Q(n9396) );
  nnd2s1 U9434 ( .DIN1(n9232), .DIN2(n8764), .Q(n9397) );
  nnd2s1 U9435 ( .DIN1(n7891), .DIN2(n9398), .Q(n9395) );
  nnd2s1 U9436 ( .DIN1(n8731), .DIN2(n8105), .Q(n9398) );
  nor2s1 U9437 ( .DIN1(n7899), .DIN2(n9191), .Q(n8731) );
  nnd2s1 U9438 ( .DIN1(n7892), .DIN2(n9399), .Q(n9394) );
  nnd2s1 U9439 ( .DIN1(n7893), .DIN2(n9386), .Q(n9393) );
  nnd2s1 U9440 ( .DIN1(n8768), .DIN2(n7911), .Q(n9386) );
  hi1s1 U9441 ( .DIN(n5703), .Q(n9260) );
  nnd2s1 U9442 ( .DIN1(n9400), .DIN2(n9401), .Q(N227) );
  nnd2s1 U9443 ( .DIN1(n9402), .DIN2(n1623), .Q(n9401) );
  xor2s1 U9444 ( .DIN1(n9403), .DIN2(n9404), .Q(n9402) );
  xor2s1 U9445 ( .DIN1(n8798), .DIN2(n9405), .Q(n9404) );
  xor2s1 U9446 ( .DIN1(n9406), .DIN2(n7620), .Q(n9405) );
  xor2s1 U9447 ( .DIN1(n5703), .DIN2(n5078), .Q(n7620) );
  or3s1 U9448 ( .DIN1(n9407), .DIN2(n9408), .DIN3(n9409), .Q(n5078) );
  nnd4s1 U9449 ( .DIN1(n9410), .DIN2(n8398), .DIN3(n9411), .DIN4(n9412), 
        .Q(n9409) );
  and3s1 U9450 ( .DIN1(n7801), .DIN2(n9279), .DIN3(n9268), .Q(n9412) );
  nor4s1 U9451 ( .DIN1(n9413), .DIN2(n9414), .DIN3(n9415), .DIN4(n9416), 
        .Q(n9268) );
  nnd4s1 U9452 ( .DIN1(n9417), .DIN2(n8905), .DIN3(n9418), .DIN4(n9419), 
        .Q(n9416) );
  nnd2s1 U9453 ( .DIN1(n8160), .DIN2(n7840), .Q(n9419) );
  nnd2s1 U9454 ( .DIN1(n7812), .DIN2(n8163), .Q(n9418) );
  nnd2s1 U9455 ( .DIN1(n7821), .DIN2(n8888), .Q(n8905) );
  nnd2s1 U9456 ( .DIN1(n7959), .DIN2(n8409), .Q(n9417) );
  nnd3s1 U9457 ( .DIN1(n9420), .DIN2(n9421), .DIN3(n9422), .Q(n9415) );
  nnd2s1 U9458 ( .DIN1(n7827), .DIN2(n9423), .Q(n9422) );
  nnd2s1 U9459 ( .DIN1(n7817), .DIN2(n9424), .Q(n9421) );
  nnd2s1 U9460 ( .DIN1(n7965), .DIN2(n7962), .Q(n9424) );
  nnd2s1 U9461 ( .DIN1(n7948), .DIN2(n9425), .Q(n9420) );
  nnd2s1 U9462 ( .DIN1(n7953), .DIN2(n7837), .Q(n9425) );
  nor2s1 U9463 ( .DIN1(n8824), .DIN2(n8146), .Q(n9414) );
  nor2s1 U9464 ( .DIN1(n8170), .DIN2(n8163), .Q(n8824) );
  nor2s1 U9465 ( .DIN1(n9426), .DIN2(n8818), .Q(n9413) );
  nor2s1 U9466 ( .DIN1(n8129), .DIN2(n8128), .Q(n9426) );
  nor2s1 U9467 ( .DIN1(n9427), .DIN2(n9428), .Q(n9279) );
  nnd4s1 U9468 ( .DIN1(n9429), .DIN2(n9430), .DIN3(n8931), .DIN4(n9431), 
        .Q(n9428) );
  nnd2s1 U9469 ( .DIN1(n7948), .DIN2(n7955), .Q(n9431) );
  nnd2s1 U9470 ( .DIN1(n8475), .DIN2(n7838), .Q(n7955) );
  nnd2s1 U9471 ( .DIN1(n7959), .DIN2(n7820), .Q(n8931) );
  nnd2s1 U9472 ( .DIN1(n8433), .DIN2(n8409), .Q(n9430) );
  nnd2s1 U9473 ( .DIN1(n7812), .DIN2(n7963), .Q(n9429) );
  nnd4s1 U9474 ( .DIN1(n9432), .DIN2(n9433), .DIN3(n9434), .DIN4(n9435), 
        .Q(n9427) );
  nnd2s1 U9475 ( .DIN1(n7821), .DIN2(n9436), .Q(n9435) );
  nnd2s1 U9476 ( .DIN1(n8825), .DIN2(n8419), .Q(n9436) );
  nnd2s1 U9477 ( .DIN1(n8160), .DIN2(n9437), .Q(n9434) );
  nnd2s1 U9478 ( .DIN1(n8154), .DIN2(n8169), .Q(n9437) );
  nnd2s1 U9479 ( .DIN1(n8130), .DIN2(n9438), .Q(n9433) );
  nnd3s1 U9480 ( .DIN1(n7966), .DIN2(n7962), .DIN3(n7952), .Q(n9438) );
  nnd2s1 U9481 ( .DIN1(n8147), .DIN2(n9439), .Q(n9432) );
  nnd4s1 U9482 ( .DIN1(n8137), .DIN2(n8154), .DIN3(n8422), .DIN4(n7965), 
        .Q(n9439) );
  nor2s1 U9483 ( .DIN1(n9440), .DIN2(n9441), .Q(n7801) );
  nnd4s1 U9484 ( .DIN1(n9442), .DIN2(n9443), .DIN3(n9444), .DIN4(n9445), 
        .Q(n9441) );
  nnd2s1 U9485 ( .DIN1(n7822), .DIN2(n8441), .Q(n9445) );
  nnd2s1 U9486 ( .DIN1(n8152), .DIN2(n7837), .Q(n8441) );
  nnd2s1 U9487 ( .DIN1(n7818), .DIN2(n7819), .Q(n9444) );
  nnd2s1 U9488 ( .DIN1(n7811), .DIN2(n8129), .Q(n9443) );
  nnd2s1 U9489 ( .DIN1(n8170), .DIN2(n8432), .Q(n9442) );
  nnd4s1 U9490 ( .DIN1(n9446), .DIN2(n9447), .DIN3(n9448), .DIN4(n9449), 
        .Q(n9440) );
  nnd2s1 U9491 ( .DIN1(n7947), .DIN2(n9450), .Q(n9449) );
  or2s1 U9492 ( .DIN1(n8934), .DIN2(n7821), .Q(n9450) );
  nnd2s1 U9493 ( .DIN1(n8140), .DIN2(n9451), .Q(n9448) );
  nnd2s1 U9494 ( .DIN1(n7952), .DIN2(n8149), .Q(n9451) );
  nnd2s1 U9495 ( .DIN1(n7812), .DIN2(n9452), .Q(n9447) );
  nnd2s1 U9496 ( .DIN1(n8457), .DIN2(n7838), .Q(n9452) );
  nnd2s1 U9497 ( .DIN1(n7835), .DIN2(n9453), .Q(n9446) );
  nnd3s1 U9498 ( .DIN1(n8457), .DIN2(n8453), .DIN3(n9454), .Q(n9453) );
  nnd2s1 U9499 ( .DIN1(n7822), .DIN2(n8160), .Q(n8398) );
  nnd2s1 U9500 ( .DIN1(n8433), .DIN2(n7835), .Q(n9410) );
  nnd3s1 U9501 ( .DIN1(n9455), .DIN2(n9456), .DIN3(n9457), .Q(n9408) );
  nnd2s1 U9502 ( .DIN1(n7959), .DIN2(n8139), .Q(n9457) );
  nnd2s1 U9503 ( .DIN1(n7821), .DIN2(n7818), .Q(n9456) );
  nnd2s1 U9504 ( .DIN1(n8409), .DIN2(n7810), .Q(n9455) );
  nnd4s1 U9505 ( .DIN1(n9458), .DIN2(n9459), .DIN3(n9460), .DIN4(n9461), 
        .Q(n9407) );
  nnd2s1 U9506 ( .DIN1(n8883), .DIN2(n9462), .Q(n9461) );
  nnd2s1 U9507 ( .DIN1(n8449), .DIN2(n8418), .Q(n9462) );
  nnd2s1 U9508 ( .DIN1(n7827), .DIN2(n9463), .Q(n9460) );
  nnd2s1 U9509 ( .DIN1(n8818), .DIN2(n8453), .Q(n9463) );
  nnd2s1 U9510 ( .DIN1(n8128), .DIN2(n9464), .Q(n9459) );
  nnd2s1 U9511 ( .DIN1(n8138), .DIN2(n8475), .Q(n9464) );
  nor2s1 U9512 ( .DIN1(n7811), .DIN2(n8163), .Q(n8138) );
  nnd2s1 U9513 ( .DIN1(n8129), .DIN2(n9465), .Q(n9458) );
  nnd3s1 U9514 ( .DIN1(n8452), .DIN2(n8450), .DIN3(n7953), .Q(n9465) );
  nor2s1 U9515 ( .DIN1(n7839), .DIN2(n8163), .Q(n7953) );
  or3s1 U9516 ( .DIN1(n9466), .DIN2(n9467), .DIN3(n9468), .Q(n5703) );
  nnd4s1 U9517 ( .DIN1(n9469), .DIN2(n8481), .DIN3(n9470), .DIN4(n9471), 
        .Q(n9468) );
  and3s1 U9518 ( .DIN1(n9472), .DIN2(n9473), .DIN3(n9307), .Q(n9471) );
  nor4s1 U9519 ( .DIN1(n9474), .DIN2(n9475), .DIN3(n9476), .DIN4(n9477), 
        .Q(n9307) );
  nnd4s1 U9520 ( .DIN1(n9478), .DIN2(n9049), .DIN3(n9479), .DIN4(n9480), 
        .Q(n9477) );
  nnd2s1 U9521 ( .DIN1(n8221), .DIN2(n9046), .Q(n9480) );
  nnd2s1 U9522 ( .DIN1(n8187), .DIN2(n8225), .Q(n9479) );
  nnd2s1 U9523 ( .DIN1(n8204), .DIN2(n9031), .Q(n9049) );
  nnd2s1 U9524 ( .DIN1(n7997), .DIN2(n8493), .Q(n9478) );
  nnd3s1 U9525 ( .DIN1(n9481), .DIN2(n9482), .DIN3(n9483), .Q(n9476) );
  nnd2s1 U9526 ( .DIN1(n8562), .DIN2(n9484), .Q(n9483) );
  nnd2s1 U9527 ( .DIN1(n8492), .DIN2(n9485), .Q(n9482) );
  nnd2s1 U9528 ( .DIN1(n8003), .DIN2(n8000), .Q(n9485) );
  nnd2s1 U9529 ( .DIN1(n7984), .DIN2(n9486), .Q(n9481) );
  nnd2s1 U9530 ( .DIN1(n7989), .DIN2(n9025), .Q(n9486) );
  nor2s1 U9531 ( .DIN1(n8966), .DIN2(n8206), .Q(n9475) );
  nor2s1 U9532 ( .DIN1(n8233), .DIN2(n8225), .Q(n8966) );
  nor2s1 U9533 ( .DIN1(n9487), .DIN2(n8959), .Q(n9474) );
  nor2s1 U9534 ( .DIN1(n8185), .DIN2(n8197), .Q(n9487) );
  nnd2s1 U9535 ( .DIN1(n8198), .DIN2(n8221), .Q(n8481) );
  nnd2s1 U9536 ( .DIN1(n8519), .DIN2(n7992), .Q(n9469) );
  nnd3s1 U9537 ( .DIN1(n9488), .DIN2(n9489), .DIN3(n9490), .Q(n9467) );
  nnd2s1 U9538 ( .DIN1(n7997), .DIN2(n8196), .Q(n9490) );
  nnd2s1 U9539 ( .DIN1(n8204), .DIN2(n8494), .Q(n9489) );
  nnd2s1 U9540 ( .DIN1(n8493), .DIN2(n7983), .Q(n9488) );
  nnd4s1 U9541 ( .DIN1(n9491), .DIN2(n9492), .DIN3(n9493), .DIN4(n9494), 
        .Q(n9466) );
  nnd2s1 U9542 ( .DIN1(n9026), .DIN2(n9495), .Q(n9494) );
  nnd2s1 U9543 ( .DIN1(n8535), .DIN2(n8504), .Q(n9495) );
  nnd2s1 U9544 ( .DIN1(n8562), .DIN2(n9496), .Q(n9493) );
  nnd2s1 U9545 ( .DIN1(n8959), .DIN2(n8539), .Q(n9496) );
  nnd2s1 U9546 ( .DIN1(n8197), .DIN2(n9497), .Q(n9492) );
  nnd2s1 U9547 ( .DIN1(n8195), .DIN2(n8564), .Q(n9497) );
  nor2s1 U9548 ( .DIN1(n8005), .DIN2(n8225), .Q(n8195) );
  nnd2s1 U9549 ( .DIN1(n8185), .DIN2(n9498), .Q(n9491) );
  nnd3s1 U9550 ( .DIN1(n8538), .DIN2(n8536), .DIN3(n7989), .Q(n9498) );
  nor2s1 U9551 ( .DIN1(n8230), .DIN2(n8225), .Q(n7989) );
  xor2s1 U9552 ( .DIN1(n5054), .DIN2(n9499), .Q(n9403) );
  xor2s1 U9553 ( .DIN1(w0[1]), .DIN2(n5030), .Q(n9499) );
  nor4s1 U9554 ( .DIN1(n9500), .DIN2(n9501), .DIN3(n9502), .DIN4(n9503), 
        .Q(n5030) );
  nnd4s1 U9555 ( .DIN1(n8651), .DIN2(n8327), .DIN3(n9504), .DIN4(n9505), 
        .Q(n9503) );
  nnd2s1 U9556 ( .DIN1(n8022), .DIN2(n8700), .Q(n9505) );
  nnd2s1 U9557 ( .DIN1(n8069), .DIN2(n8667), .Q(n9504) );
  nnd2s1 U9558 ( .DIN1(n8063), .DIN2(n8584), .Q(n8327) );
  nnd2s1 U9559 ( .DIN1(n8034), .DIN2(n7861), .Q(n8651) );
  nnd4s1 U9560 ( .DIN1(n9506), .DIN2(n9507), .DIN3(n9508), .DIN4(n9509), 
        .Q(n9502) );
  nnd2s1 U9561 ( .DIN1(n7870), .DIN2(n9510), .Q(n9509) );
  nnd2s1 U9562 ( .DIN1(n7868), .DIN2(n8278), .Q(n9510) );
  nnd2s1 U9563 ( .DIN1(n8023), .DIN2(n9511), .Q(n9508) );
  nnd2s1 U9564 ( .DIN1(n8252), .DIN2(n8318), .Q(n9511) );
  nnd2s1 U9565 ( .DIN1(n8316), .DIN2(n8079), .Q(n9507) );
  nnd2s1 U9566 ( .DIN1(n8054), .DIN2(n7869), .Q(n8079) );
  or2s1 U9567 ( .DIN1(n8074), .DIN2(n8047), .Q(n9506) );
  nor2s1 U9568 ( .DIN1(n8030), .DIN2(n8021), .Q(n8047) );
  nnd3s1 U9569 ( .DIN1(n9091), .DIN2(n9512), .DIN3(n9513), .Q(n9501) );
  nor4s1 U9570 ( .DIN1(n9514), .DIN2(n9515), .DIN3(n9516), .DIN4(n9517), 
        .Q(n9091) );
  nnd4s1 U9571 ( .DIN1(n9518), .DIN2(n9519), .DIN3(n9520), .DIN4(n9521), 
        .Q(n9517) );
  nor2s1 U9572 ( .DIN1(n9522), .DIN2(n9523), .Q(n9521) );
  nor2s1 U9573 ( .DIN1(n8059), .DIN2(n7877), .Q(n9523) );
  nor2s1 U9574 ( .DIN1(n8051), .DIN2(n8252), .Q(n9522) );
  nnd2s1 U9575 ( .DIN1(n8062), .DIN2(n8254), .Q(n9520) );
  or2s1 U9576 ( .DIN1(n8045), .DIN2(n8280), .Q(n9519) );
  nor2s1 U9577 ( .DIN1(n7861), .DIN2(n8699), .Q(n8280) );
  nnd2s1 U9578 ( .DIN1(n8649), .DIN2(n8021), .Q(n9518) );
  nnd3s1 U9579 ( .DIN1(n9524), .DIN2(n9525), .DIN3(n9526), .Q(n9516) );
  nnd2s1 U9580 ( .DIN1(n8272), .DIN2(n9527), .Q(n9526) );
  nnd2s1 U9581 ( .DIN1(n8044), .DIN2(n8284), .Q(n9527) );
  nnd2s1 U9582 ( .DIN1(n8036), .DIN2(n8256), .Q(n9525) );
  nnd2s1 U9583 ( .DIN1(n8286), .DIN2(n7869), .Q(n8256) );
  nnd2s1 U9584 ( .DIN1(n8042), .DIN2(n9528), .Q(n9524) );
  nnd2s1 U9585 ( .DIN1(n8048), .DIN2(n8586), .Q(n9528) );
  nor2s1 U9586 ( .DIN1(n9529), .DIN2(n7857), .Q(n9515) );
  nor2s1 U9587 ( .DIN1(n8254), .DIN2(n7866), .Q(n9529) );
  nor2s1 U9588 ( .DIN1(n9530), .DIN2(n7868), .Q(n9514) );
  nor2s1 U9589 ( .DIN1(n8063), .DIN2(n8052), .Q(n9530) );
  nnd4s1 U9590 ( .DIN1(n9357), .DIN2(n9531), .DIN3(n9532), .DIN4(n9533), 
        .Q(n9500) );
  nnd2s1 U9591 ( .DIN1(n8062), .DIN2(n8049), .Q(n9533) );
  nnd2s1 U9592 ( .DIN1(n8310), .DIN2(n8078), .Q(n9532) );
  nnd2s1 U9593 ( .DIN1(n8271), .DIN2(n8021), .Q(n9531) );
  nor3s1 U9594 ( .DIN1(n9534), .DIN2(n9535), .DIN3(n9536), .Q(n9357) );
  nnd4s1 U9595 ( .DIN1(n9537), .DIN2(n9538), .DIN3(n9096), .DIN4(n9539), 
        .Q(n9536) );
  and3s1 U9596 ( .DIN1(n9540), .DIN2(n9541), .DIN3(n9542), .Q(n9539) );
  nnd2s1 U9597 ( .DIN1(n7866), .DIN2(n8272), .Q(n9542) );
  nnd2s1 U9598 ( .DIN1(n8316), .DIN2(n8257), .Q(n9541) );
  nnd2s1 U9599 ( .DIN1(n8064), .DIN2(n8049), .Q(n9540) );
  nor2s1 U9600 ( .DIN1(n9543), .DIN2(n9544), .Q(n9096) );
  nnd4s1 U9601 ( .DIN1(n9545), .DIN2(n9546), .DIN3(n9547), .DIN4(n9548), 
        .Q(n9544) );
  nnd2s1 U9602 ( .DIN1(n7866), .DIN2(n9549), .Q(n9548) );
  nnd2s1 U9603 ( .DIN1(n8591), .DIN2(n7878), .Q(n9549) );
  nnd2s1 U9604 ( .DIN1(n8021), .DIN2(n9550), .Q(n9547) );
  nnd3s1 U9605 ( .DIN1(n7859), .DIN2(n7868), .DIN3(n7877), .Q(n9550) );
  nnd2s1 U9606 ( .DIN1(n8034), .DIN2(n8062), .Q(n9546) );
  nnd2s1 U9607 ( .DIN1(n8023), .DIN2(n8316), .Q(n9545) );
  nnd4s1 U9608 ( .DIN1(n9551), .DIN2(n9552), .DIN3(n9553), .DIN4(n9554), 
        .Q(n9543) );
  nnd2s1 U9609 ( .DIN1(n8649), .DIN2(n9555), .Q(n9554) );
  nnd2s1 U9610 ( .DIN1(n8590), .DIN2(n8253), .Q(n9555) );
  nnd2s1 U9611 ( .DIN1(n8037), .DIN2(n9556), .Q(n9553) );
  nnd2s1 U9612 ( .DIN1(n8044), .DIN2(n8077), .Q(n9556) );
  nnd2s1 U9613 ( .DIN1(n7853), .DIN2(n9557), .Q(n9552) );
  nnd2s1 U9614 ( .DIN1(n8627), .DIN2(n8032), .Q(n9557) );
  nor2s1 U9615 ( .DIN1(n8699), .DIN2(n8310), .Q(n8627) );
  nnd2s1 U9616 ( .DIN1(n8052), .DIN2(n9558), .Q(n9551) );
  nnd2s1 U9617 ( .DIN1(n7878), .DIN2(n8278), .Q(n9558) );
  nnd3s1 U9618 ( .DIN1(n9559), .DIN2(n9560), .DIN3(n9561), .Q(n9535) );
  nnd2s1 U9619 ( .DIN1(n8023), .DIN2(n8078), .Q(n9561) );
  nnd2s1 U9620 ( .DIN1(n8254), .DIN2(n8649), .Q(n9560) );
  nnd2s1 U9621 ( .DIN1(n8034), .DIN2(n8042), .Q(n9559) );
  nnd4s1 U9622 ( .DIN1(n9562), .DIN2(n9563), .DIN3(n9564), .DIN4(n9565), 
        .Q(n9534) );
  nnd2s1 U9623 ( .DIN1(n8271), .DIN2(n9566), .Q(n9565) );
  nnd2s1 U9624 ( .DIN1(n8590), .DIN2(n8318), .Q(n9566) );
  nnd2s1 U9625 ( .DIN1(n8310), .DIN2(n9567), .Q(n9564) );
  nnd4s1 U9626 ( .DIN1(n8318), .DIN2(n8045), .DIN3(n8284), .DIN4(n8260), 
        .Q(n9567) );
  nnd2s1 U9627 ( .DIN1(n8069), .DIN2(n8624), .Q(n9563) );
  nnd2s1 U9628 ( .DIN1(n8277), .DIN2(n7859), .Q(n8624) );
  nnd2s1 U9629 ( .DIN1(n7853), .DIN2(n8261), .Q(n9562) );
  nnd2s1 U9630 ( .DIN1(n7857), .DIN2(n7869), .Q(n8261) );
  or3s1 U9631 ( .DIN1(n9568), .DIN2(n9569), .DIN3(n9570), .Q(n5054) );
  nnd4s1 U9632 ( .DIN1(n9571), .DIN2(n8713), .DIN3(n9572), .DIN4(n9573), 
        .Q(n9570) );
  and3s1 U9633 ( .DIN1(n7882), .DIN2(n9375), .DIN3(n9364), .Q(n9573) );
  nor4s1 U9634 ( .DIN1(n9574), .DIN2(n9575), .DIN3(n9576), .DIN4(n9577), 
        .Q(n9364) );
  nnd4s1 U9635 ( .DIN1(n9578), .DIN2(n9213), .DIN3(n9579), .DIN4(n9580), 
        .Q(n9577) );
  nnd2s1 U9636 ( .DIN1(n8370), .DIN2(n7921), .Q(n9580) );
  nnd2s1 U9637 ( .DIN1(n7893), .DIN2(n8373), .Q(n9579) );
  nnd2s1 U9638 ( .DIN1(n7902), .DIN2(n9196), .Q(n9213) );
  nnd2s1 U9639 ( .DIN1(n8102), .DIN2(n8724), .Q(n9578) );
  nnd3s1 U9640 ( .DIN1(n9581), .DIN2(n9582), .DIN3(n9583), .Q(n9576) );
  nnd2s1 U9641 ( .DIN1(n7908), .DIN2(n9584), .Q(n9583) );
  nnd2s1 U9642 ( .DIN1(n7898), .DIN2(n9585), .Q(n9582) );
  nnd2s1 U9643 ( .DIN1(n8108), .DIN2(n8105), .Q(n9585) );
  nnd2s1 U9644 ( .DIN1(n8091), .DIN2(n9586), .Q(n9581) );
  nnd2s1 U9645 ( .DIN1(n8096), .DIN2(n7918), .Q(n9586) );
  nor2s1 U9646 ( .DIN1(n9132), .DIN2(n8356), .Q(n9575) );
  nor2s1 U9647 ( .DIN1(n8380), .DIN2(n8373), .Q(n9132) );
  nor2s1 U9648 ( .DIN1(n9587), .DIN2(n9126), .Q(n9574) );
  nor2s1 U9649 ( .DIN1(n8339), .DIN2(n8338), .Q(n9587) );
  nor2s1 U9650 ( .DIN1(n9588), .DIN2(n9589), .Q(n9375) );
  nnd4s1 U9651 ( .DIN1(n9590), .DIN2(n9591), .DIN3(n9239), .DIN4(n9592), 
        .Q(n9589) );
  nnd2s1 U9652 ( .DIN1(n8091), .DIN2(n8098), .Q(n9592) );
  nnd2s1 U9653 ( .DIN1(n8790), .DIN2(n7919), .Q(n8098) );
  nnd2s1 U9654 ( .DIN1(n8102), .DIN2(n7901), .Q(n9239) );
  nnd2s1 U9655 ( .DIN1(n8748), .DIN2(n8724), .Q(n9591) );
  nnd2s1 U9656 ( .DIN1(n7893), .DIN2(n8106), .Q(n9590) );
  nnd4s1 U9657 ( .DIN1(n9593), .DIN2(n9594), .DIN3(n9595), .DIN4(n9596), 
        .Q(n9588) );
  nnd2s1 U9658 ( .DIN1(n7902), .DIN2(n9597), .Q(n9596) );
  nnd2s1 U9659 ( .DIN1(n9133), .DIN2(n8734), .Q(n9597) );
  nnd2s1 U9660 ( .DIN1(n8370), .DIN2(n9598), .Q(n9595) );
  nnd2s1 U9661 ( .DIN1(n8364), .DIN2(n8379), .Q(n9598) );
  nnd2s1 U9662 ( .DIN1(n8340), .DIN2(n9599), .Q(n9594) );
  nnd3s1 U9663 ( .DIN1(n8109), .DIN2(n8105), .DIN3(n8095), .Q(n9599) );
  nnd2s1 U9664 ( .DIN1(n8357), .DIN2(n9600), .Q(n9593) );
  nnd4s1 U9665 ( .DIN1(n8347), .DIN2(n8364), .DIN3(n8737), .DIN4(n8108), 
        .Q(n9600) );
  nor2s1 U9666 ( .DIN1(n9601), .DIN2(n9602), .Q(n7882) );
  nnd4s1 U9667 ( .DIN1(n9603), .DIN2(n9604), .DIN3(n9605), .DIN4(n9606), 
        .Q(n9602) );
  nnd2s1 U9668 ( .DIN1(n7903), .DIN2(n8756), .Q(n9606) );
  nnd2s1 U9669 ( .DIN1(n8362), .DIN2(n7918), .Q(n8756) );
  nnd2s1 U9670 ( .DIN1(n7899), .DIN2(n7900), .Q(n9605) );
  nnd2s1 U9671 ( .DIN1(n7892), .DIN2(n8339), .Q(n9604) );
  nnd2s1 U9672 ( .DIN1(n8380), .DIN2(n8747), .Q(n9603) );
  nnd4s1 U9673 ( .DIN1(n9607), .DIN2(n9608), .DIN3(n9609), .DIN4(n9610), 
        .Q(n9601) );
  nnd2s1 U9674 ( .DIN1(n8090), .DIN2(n9611), .Q(n9610) );
  or2s1 U9675 ( .DIN1(n9242), .DIN2(n7902), .Q(n9611) );
  nnd2s1 U9676 ( .DIN1(n8350), .DIN2(n9612), .Q(n9609) );
  nnd2s1 U9677 ( .DIN1(n8095), .DIN2(n8359), .Q(n9612) );
  nnd2s1 U9678 ( .DIN1(n7893), .DIN2(n9613), .Q(n9608) );
  nnd2s1 U9679 ( .DIN1(n8772), .DIN2(n7919), .Q(n9613) );
  nnd2s1 U9680 ( .DIN1(n7916), .DIN2(n9614), .Q(n9607) );
  nnd3s1 U9681 ( .DIN1(n8772), .DIN2(n8768), .DIN3(n9615), .Q(n9614) );
  nnd2s1 U9682 ( .DIN1(n7903), .DIN2(n8370), .Q(n8713) );
  nnd2s1 U9683 ( .DIN1(n8748), .DIN2(n7916), .Q(n9571) );
  nnd3s1 U9684 ( .DIN1(n9616), .DIN2(n9617), .DIN3(n9618), .Q(n9569) );
  nnd2s1 U9685 ( .DIN1(n8102), .DIN2(n8349), .Q(n9618) );
  nnd2s1 U9686 ( .DIN1(n7902), .DIN2(n7899), .Q(n9617) );
  nnd2s1 U9687 ( .DIN1(n8724), .DIN2(n7891), .Q(n9616) );
  nnd4s1 U9688 ( .DIN1(n9619), .DIN2(n9620), .DIN3(n9621), .DIN4(n9622), 
        .Q(n9568) );
  nnd2s1 U9689 ( .DIN1(n9191), .DIN2(n9623), .Q(n9622) );
  nnd2s1 U9690 ( .DIN1(n8764), .DIN2(n8733), .Q(n9623) );
  nnd2s1 U9691 ( .DIN1(n7908), .DIN2(n9624), .Q(n9621) );
  nnd2s1 U9692 ( .DIN1(n9126), .DIN2(n8768), .Q(n9624) );
  nnd2s1 U9693 ( .DIN1(n8338), .DIN2(n9625), .Q(n9620) );
  nnd2s1 U9694 ( .DIN1(n8348), .DIN2(n8790), .Q(n9625) );
  nor2s1 U9695 ( .DIN1(n7892), .DIN2(n8373), .Q(n8348) );
  nnd2s1 U9696 ( .DIN1(n8339), .DIN2(n9626), .Q(n9619) );
  nnd3s1 U9697 ( .DIN1(n8767), .DIN2(n8765), .DIN3(n8096), .Q(n9626) );
  nor2s1 U9698 ( .DIN1(n7920), .DIN2(n8373), .Q(n8096) );
  nnd2s1 U9699 ( .DIN1(n9627), .DIN2(n1603), .Q(n9400) );
  xor2s1 U9700 ( .DIN1(w0[1]), .DIN2(text_in_r[97]), .Q(n9627) );
  nnd2s1 U9701 ( .DIN1(n9628), .DIN2(n9629), .Q(N226) );
  nnd2s1 U9702 ( .DIN1(n9630), .DIN2(n1624), .Q(n9629) );
  xor2s1 U9703 ( .DIN1(n9631), .DIN2(n9632), .Q(n9630) );
  xor2s1 U9704 ( .DIN1(n7628), .DIN2(n8391), .Q(n9632) );
  hi1s1 U9705 ( .DIN(n8798), .Q(n8391) );
  xor2s1 U9706 ( .DIN1(n6115), .DIN2(n5037), .Q(n8798) );
  nor3s1 U9707 ( .DIN1(n9633), .DIN2(n9634), .DIN3(n9635), .Q(n5037) );
  nnd4s1 U9708 ( .DIN1(n9341), .DIN2(n9513), .DIN3(n9092), .DIN4(n9636), 
        .Q(n9635) );
  and4s1 U9709 ( .DIN1(n9537), .DIN2(n9637), .DIN3(n9638), .DIN4(n8295), 
        .Q(n9636) );
  nnd2s1 U9710 ( .DIN1(n8049), .DIN2(n8035), .Q(n8295) );
  nnd2s1 U9711 ( .DIN1(n8052), .DIN2(n8037), .Q(n9638) );
  nnd2s1 U9712 ( .DIN1(n7853), .DIN2(n8584), .Q(n9637) );
  and4s1 U9713 ( .DIN1(n9639), .DIN2(n9640), .DIN3(n9641), .DIN4(n9642), 
        .Q(n9537) );
  and4s1 U9714 ( .DIN1(n9643), .DIN2(n9644), .DIN3(n9645), .DIN4(n9646), 
        .Q(n9642) );
  nnd2s1 U9715 ( .DIN1(n8062), .DIN2(n7853), .Q(n9646) );
  nnd2s1 U9716 ( .DIN1(n7852), .DIN2(n8072), .Q(n9645) );
  nnd2s1 U9717 ( .DIN1(n7870), .DIN2(n8584), .Q(n9644) );
  nnd2s1 U9718 ( .DIN1(n8254), .DIN2(n8257), .Q(n9643) );
  and3s1 U9719 ( .DIN1(n9647), .DIN2(n9648), .DIN3(n9649), .Q(n9641) );
  nnd2s1 U9720 ( .DIN1(n8023), .DIN2(n9650), .Q(n9649) );
  nnd3s1 U9721 ( .DIN1(n9651), .DIN2(n8260), .DIN3(n8077), .Q(n9650) );
  nnd2s1 U9722 ( .DIN1(n8078), .DIN2(n8643), .Q(n9648) );
  nnd2s1 U9723 ( .DIN1(n8281), .DIN2(n8071), .Q(n8643) );
  nnd2s1 U9724 ( .DIN1(n8037), .DIN2(n9652), .Q(n9647) );
  nnd2s1 U9725 ( .DIN1(n8252), .DIN2(n8045), .Q(n9652) );
  nnd2s1 U9726 ( .DIN1(n8316), .DIN2(n9653), .Q(n9640) );
  nnd4s1 U9727 ( .DIN1(n7877), .DIN2(n7868), .DIN3(n7878), .DIN4(n8074), 
        .Q(n9653) );
  nnd2s1 U9728 ( .DIN1(n8063), .DIN2(n8272), .Q(n9639) );
  nor3s1 U9729 ( .DIN1(n9654), .DIN2(n9655), .DIN3(n9656), .Q(n9092) );
  nnd4s1 U9730 ( .DIN1(n9512), .DIN2(n9538), .DIN3(n9342), .DIN4(n9657), 
        .Q(n9656) );
  and4s1 U9731 ( .DIN1(n9658), .DIN2(n9659), .DIN3(n9660), .DIN4(n9661), 
        .Q(n9657) );
  nnd2s1 U9732 ( .DIN1(n8069), .DIN2(n8699), .Q(n9661) );
  nnd2s1 U9733 ( .DIN1(n7866), .DIN2(n8064), .Q(n9660) );
  nnd2s1 U9734 ( .DIN1(n8023), .DIN2(n8254), .Q(n9659) );
  hi1s1 U9735 ( .DIN(n8277), .Q(n8023) );
  nnd2s1 U9736 ( .DIN1(n8030), .DIN2(n8035), .Q(n9658) );
  nor2s1 U9737 ( .DIN1(n9662), .DIN2(n9663), .Q(n9342) );
  nnd4s1 U9738 ( .DIN1(n8569), .DIN2(n9664), .DIN3(n9665), .DIN4(n9666), 
        .Q(n9663) );
  nnd2s1 U9739 ( .DIN1(n8052), .DIN2(n9340), .Q(n9666) );
  nnd2s1 U9740 ( .DIN1(n8277), .DIN2(n8071), .Q(n9340) );
  nnd2s1 U9741 ( .DIN1(n8316), .DIN2(n8699), .Q(n9665) );
  nnd2s1 U9742 ( .DIN1(n8064), .DIN2(n7875), .Q(n9664) );
  nnd2s1 U9743 ( .DIN1(n7866), .DIN2(n8584), .Q(n8569) );
  nnd4s1 U9744 ( .DIN1(n9667), .DIN2(n9668), .DIN3(n9669), .DIN4(n9670), 
        .Q(n9662) );
  nnd2s1 U9745 ( .DIN1(n8078), .DIN2(n9671), .Q(n9670) );
  nnd2s1 U9746 ( .DIN1(n8032), .DIN2(n8074), .Q(n9671) );
  hi1s1 U9747 ( .DIN(n8586), .Q(n8078) );
  nnd2s1 U9748 ( .DIN1(n8034), .DIN2(n9672), .Q(n9669) );
  nnd3s1 U9749 ( .DIN1(n7857), .DIN2(n7868), .DIN3(n7877), .Q(n9672) );
  nnd2s1 U9750 ( .DIN1(n8049), .DIN2(n9673), .Q(n9668) );
  nnd4s1 U9751 ( .DIN1(n8278), .DIN2(n8032), .DIN3(n7878), .DIN4(n8286), 
        .Q(n9673) );
  nnd2s1 U9752 ( .DIN1(n8042), .DIN2(n7862), .Q(n9667) );
  nnd2s1 U9753 ( .DIN1(n8259), .DIN2(n8312), .Q(n7862) );
  nor4s1 U9754 ( .DIN1(n9674), .DIN2(n9675), .DIN3(n9676), .DIN4(n9677), 
        .Q(n9538) );
  nnd4s1 U9755 ( .DIN1(n9678), .DIN2(n9679), .DIN3(n9680), .DIN4(n9681), 
        .Q(n9677) );
  and3s1 U9756 ( .DIN1(n9682), .DIN2(n9683), .DIN3(n9684), .Q(n9681) );
  nnd2s1 U9757 ( .DIN1(n8030), .DIN2(n9108), .Q(n9684) );
  nnd2s1 U9758 ( .DIN1(n8051), .DIN2(n8054), .Q(n9108) );
  nnd2s1 U9759 ( .DIN1(n8649), .DIN2(n9685), .Q(n9683) );
  nnd2s1 U9760 ( .DIN1(n8586), .DIN2(n8284), .Q(n9685) );
  hi1s1 U9761 ( .DIN(n7869), .Q(n8649) );
  nnd2s1 U9762 ( .DIN1(n7852), .DIN2(n9686), .Q(n9682) );
  nnd2s1 U9763 ( .DIN1(n8077), .DIN2(n8045), .Q(n9686) );
  nnd2s1 U9764 ( .DIN1(n7866), .DIN2(n8062), .Q(n9680) );
  nnd2s1 U9765 ( .DIN1(n8072), .DIN2(n9687), .Q(n9679) );
  nnd2s1 U9766 ( .DIN1(n7857), .DIN2(n7859), .Q(n9687) );
  nnd2s1 U9767 ( .DIN1(n8584), .DIN2(n9688), .Q(n9678) );
  nnd2s1 U9768 ( .DIN1(n8076), .DIN2(n8312), .Q(n9688) );
  nnd3s1 U9769 ( .DIN1(n9689), .DIN2(n9690), .DIN3(n9691), .Q(n9676) );
  nnd2s1 U9770 ( .DIN1(n8316), .DIN2(n8272), .Q(n9691) );
  nnd2s1 U9771 ( .DIN1(n8254), .DIN2(n8271), .Q(n9690) );
  nnd2s1 U9772 ( .DIN1(n8310), .DIN2(n8036), .Q(n9689) );
  nor2s1 U9773 ( .DIN1(n7868), .DIN2(n8253), .Q(n9675) );
  nor2s1 U9774 ( .DIN1(n8260), .DIN2(n8591), .Q(n9674) );
  nor4s1 U9775 ( .DIN1(n9692), .DIN2(n9693), .DIN3(n9694), .DIN4(n9695), 
        .Q(n9512) );
  nnd4s1 U9776 ( .DIN1(n9696), .DIN2(n9697), .DIN3(n9698), .DIN4(n9699), 
        .Q(n9695) );
  nnd2s1 U9777 ( .DIN1(n8063), .DIN2(n8271), .Q(n9699) );
  nnd2s1 U9778 ( .DIN1(n8022), .DIN2(n8036), .Q(n9698) );
  nnd2s1 U9779 ( .DIN1(n7853), .DIN2(n8042), .Q(n9697) );
  nnd2s1 U9780 ( .DIN1(n7870), .DIN2(n7861), .Q(n9696) );
  nnd3s1 U9781 ( .DIN1(n9700), .DIN2(n9701), .DIN3(n9702), .Q(n9694) );
  nnd2s1 U9782 ( .DIN1(n8064), .DIN2(n9703), .Q(n9702) );
  nnd2s1 U9783 ( .DIN1(n8077), .DIN2(n8586), .Q(n9703) );
  nnd2s1 U9784 ( .DIN1(n8034), .DIN2(n8679), .Q(n9701) );
  nnd2s1 U9785 ( .DIN1(n8074), .DIN2(n8051), .Q(n8679) );
  nnd2s1 U9786 ( .DIN1(n8062), .DIN2(n9704), .Q(n9700) );
  nnd2s1 U9787 ( .DIN1(n9705), .DIN2(n8586), .Q(n9704) );
  nor2s1 U9788 ( .DIN1(n7869), .DIN2(n8318), .Q(n9693) );
  and2s1 U9789 ( .DIN1(n7875), .DIN2(n9706), .Q(n9692) );
  nnd3s1 U9790 ( .DIN1(n7878), .DIN2(n8074), .DIN3(n7859), .Q(n9706) );
  nnd3s1 U9791 ( .DIN1(n8671), .DIN2(n9707), .DIN3(n9708), .Q(n9655) );
  nnd2s1 U9792 ( .DIN1(n8316), .DIN2(n8022), .Q(n9708) );
  hi1s1 U9793 ( .DIN(n8048), .Q(n8316) );
  nnd2s1 U9794 ( .DIN1(n8063), .DIN2(n7874), .Q(n9707) );
  nnd2s1 U9795 ( .DIN1(n8032), .DIN2(n7869), .Q(n7874) );
  hi1s1 U9796 ( .DIN(n8045), .Q(n8063) );
  nnd2s1 U9797 ( .DIN1(n9709), .DIN2(n9710), .Q(n8045) );
  nnd2s1 U9798 ( .DIN1(n8034), .DIN2(n8271), .Q(n8671) );
  hi1s1 U9799 ( .DIN(n8071), .Q(n8271) );
  hi1s1 U9800 ( .DIN(n8284), .Q(n8034) );
  nnd4s1 U9801 ( .DIN1(n9711), .DIN2(n9712), .DIN3(n9713), .DIN4(n9714), 
        .Q(n9654) );
  nnd2s1 U9802 ( .DIN1(n7870), .DIN2(n9715), .Q(n9714) );
  nnd2s1 U9803 ( .DIN1(n8074), .DIN2(n7869), .Q(n9715) );
  nnd3s1 U9804 ( .DIN1(sa33[7]), .DIN2(n1428), .DIN3(n9716), .Q(n7869) );
  nnd2s1 U9805 ( .DIN1(n7861), .DIN2(n9717), .Q(n9713) );
  nnd2s1 U9806 ( .DIN1(n8688), .DIN2(n8586), .Q(n9717) );
  hi1s1 U9807 ( .DIN(n8061), .Q(n8688) );
  nnd2s1 U9808 ( .DIN1(n8252), .DIN2(n8077), .Q(n8061) );
  nnd2s1 U9809 ( .DIN1(n8052), .DIN2(n9718), .Q(n9712) );
  nnd2s1 U9810 ( .DIN1(n8281), .DIN2(n8051), .Q(n9718) );
  or2s1 U9811 ( .DIN1(n8590), .DIN2(n8682), .Q(n9711) );
  nor2s1 U9812 ( .DIN1(n8584), .DIN2(n8062), .Q(n8682) );
  nor4s1 U9813 ( .DIN1(n9719), .DIN2(n9720), .DIN3(n9721), .DIN4(n9722), 
        .Q(n9513) );
  nnd4s1 U9814 ( .DIN1(n8618), .DIN2(n7846), .DIN3(n9723), .DIN4(n9724), 
        .Q(n9722) );
  nor2s1 U9815 ( .DIN1(n9725), .DIN2(n9726), .Q(n9724) );
  nor2s1 U9816 ( .DIN1(n8059), .DIN2(n8591), .Q(n9726) );
  nor2s1 U9817 ( .DIN1(n9651), .DIN2(n8032), .Q(n9725) );
  nnd2s1 U9818 ( .DIN1(n8049), .DIN2(n8022), .Q(n9723) );
  hi1s1 U9819 ( .DIN(n8252), .Q(n8049) );
  nnd2s1 U9820 ( .DIN1(n9727), .DIN2(n9728), .Q(n8252) );
  nnd2s1 U9821 ( .DIN1(n8042), .DIN2(n8036), .Q(n7846) );
  hi1s1 U9822 ( .DIN(n8278), .Q(n8042) );
  nnd2s1 U9823 ( .DIN1(n7875), .DIN2(n8699), .Q(n8618) );
  nnd3s1 U9824 ( .DIN1(n9729), .DIN2(n9730), .DIN3(n9731), .Q(n9721) );
  nnd2s1 U9825 ( .DIN1(n8021), .DIN2(n8302), .Q(n9731) );
  nnd2s1 U9826 ( .DIN1(n8278), .DIN2(n8054), .Q(n8302) );
  nnd3s1 U9827 ( .DIN1(n9732), .DIN2(n1382), .DIN3(sa33[6]), .Q(n8278) );
  nnd2s1 U9828 ( .DIN1(n8035), .DIN2(n9733), .Q(n9730) );
  nnd3s1 U9829 ( .DIN1(n8059), .DIN2(n8586), .DIN3(n9651), .Q(n9733) );
  hi1s1 U9830 ( .DIN(n7868), .Q(n8035) );
  nnd3s1 U9831 ( .DIN1(sa33[5]), .DIN2(n9732), .DIN3(sa33[6]), .Q(n7868) );
  nnd2s1 U9832 ( .DIN1(n8584), .DIN2(n9734), .Q(n9729) );
  nnd3s1 U9833 ( .DIN1(n8284), .DIN2(n8260), .DIN3(n8318), .Q(n9734) );
  nnd2s1 U9834 ( .DIN1(n9735), .DIN2(n9736), .Q(n8284) );
  hi1s1 U9835 ( .DIN(n8286), .Q(n8584) );
  nor2s1 U9836 ( .DIN1(n7859), .DIN2(n8586), .Q(n9720) );
  nnd2s1 U9837 ( .DIN1(n9728), .DIN2(n9710), .Q(n8586) );
  nor2s1 U9838 ( .DIN1(n8689), .DIN2(n8071), .Q(n9719) );
  nnd3s1 U9839 ( .DIN1(sa33[4]), .DIN2(n1382), .DIN3(n9737), .Q(n8071) );
  nor2s1 U9840 ( .DIN1(n7866), .DIN2(n8072), .Q(n8689) );
  nor2s1 U9841 ( .DIN1(n9738), .DIN2(n9739), .Q(n9341) );
  nnd4s1 U9842 ( .DIN1(n9740), .DIN2(n9741), .DIN3(n9742), .DIN4(n9743), 
        .Q(n9739) );
  nnd2s1 U9843 ( .DIN1(n8069), .DIN2(n8310), .Q(n9743) );
  hi1s1 U9844 ( .DIN(n7878), .Q(n8310) );
  nnd2s1 U9845 ( .DIN1(n9716), .DIN2(n9744), .Q(n7878) );
  hi1s1 U9846 ( .DIN(n8253), .Q(n8069) );
  nnd2s1 U9847 ( .DIN1(n8699), .DIN2(n8021), .Q(n9742) );
  hi1s1 U9848 ( .DIN(n8051), .Q(n8699) );
  nnd2s1 U9849 ( .DIN1(n7870), .DIN2(n8022), .Q(n9741) );
  hi1s1 U9850 ( .DIN(n8281), .Q(n8022) );
  nnd2s1 U9851 ( .DIN1(n7853), .DIN2(n8272), .Q(n9740) );
  hi1s1 U9852 ( .DIN(n7859), .Q(n8272) );
  hi1s1 U9853 ( .DIN(n8059), .Q(n7853) );
  nnd2s1 U9854 ( .DIN1(n9745), .DIN2(n9709), .Q(n8059) );
  nnd4s1 U9855 ( .DIN1(n9746), .DIN2(n9747), .DIN3(n9748), .DIN4(n9749), 
        .Q(n9738) );
  nnd2s1 U9856 ( .DIN1(n8064), .DIN2(n9750), .Q(n9749) );
  nnd2s1 U9857 ( .DIN1(n8318), .DIN2(n8312), .Q(n9750) );
  nnd2s1 U9858 ( .DIN1(n7852), .DIN2(n9751), .Q(n9748) );
  or2s1 U9859 ( .DIN1(n8700), .DIN2(n8052), .Q(n9751) );
  nnd2s1 U9860 ( .DIN1(n8312), .DIN2(n8253), .Q(n8700) );
  hi1s1 U9861 ( .DIN(n8074), .Q(n7852) );
  nnd3s1 U9862 ( .DIN1(sa33[5]), .DIN2(sa33[4]), .DIN3(n9737), .Q(n8074) );
  nnd2s1 U9863 ( .DIN1(n8037), .DIN2(n9752), .Q(n9747) );
  or2s1 U9864 ( .DIN1(n8303), .DIN2(n8021), .Q(n9752) );
  hi1s1 U9865 ( .DIN(n8260), .Q(n8021) );
  nnd2s1 U9866 ( .DIN1(n9753), .DIN2(n9710), .Q(n8260) );
  nnd2s1 U9867 ( .DIN1(n8590), .DIN2(n8048), .Q(n8303) );
  nnd2s1 U9868 ( .DIN1(n9727), .DIN2(n9753), .Q(n8048) );
  hi1s1 U9869 ( .DIN(n7857), .Q(n8037) );
  nnd3s1 U9870 ( .DIN1(sa33[5]), .DIN2(sa33[4]), .DIN3(n9744), .Q(n7857) );
  nnd2s1 U9871 ( .DIN1(n7861), .DIN2(n9754), .Q(n9746) );
  nnd3s1 U9872 ( .DIN1(n8318), .DIN2(n8253), .DIN3(n9705), .Q(n9754) );
  nor2s1 U9873 ( .DIN1(n8052), .DIN2(n8072), .Q(n9705) );
  hi1s1 U9874 ( .DIN(n8076), .Q(n8052) );
  nnd2s1 U9875 ( .DIN1(n9727), .DIN2(n9736), .Q(n8253) );
  hi1s1 U9876 ( .DIN(n8591), .Q(n7861) );
  nnd3s1 U9877 ( .DIN1(n9755), .DIN2(n9756), .DIN3(n9757), .Q(n9634) );
  nnd2s1 U9878 ( .DIN1(n7870), .DIN2(n8064), .Q(n9757) );
  hi1s1 U9879 ( .DIN(n7877), .Q(n8064) );
  nnd3s1 U9880 ( .DIN1(sa33[6]), .DIN2(sa33[7]), .DIN3(n9716), .Q(n7877) );
  hi1s1 U9881 ( .DIN(n8044), .Q(n7870) );
  nnd2s1 U9882 ( .DIN1(n9745), .DIN2(n9728), .Q(n8044) );
  nnd2s1 U9883 ( .DIN1(n8072), .DIN2(n8667), .Q(n9756) );
  nnd2s1 U9884 ( .DIN1(n8286), .DIN2(n8051), .Q(n8667) );
  nnd3s1 U9885 ( .DIN1(n9732), .DIN2(n1428), .DIN3(sa33[5]), .Q(n8051) );
  nnd3s1 U9886 ( .DIN1(sa33[6]), .DIN2(sa33[7]), .DIN3(n9758), .Q(n8286) );
  hi1s1 U9887 ( .DIN(n9651), .Q(n8072) );
  nnd2s1 U9888 ( .DIN1(n9736), .DIN2(n9710), .Q(n9651) );
  and2s1 U9889 ( .DIN1(sa33[0]), .DIN2(n1537), .Q(n9710) );
  nnd2s1 U9890 ( .DIN1(n8062), .DIN2(n8036), .Q(n9755) );
  hi1s1 U9891 ( .DIN(n8077), .Q(n8036) );
  nnd2s1 U9892 ( .DIN1(n9735), .DIN2(n9728), .Q(n8077) );
  and2s1 U9893 ( .DIN1(sa33[3]), .DIN2(n1529), .Q(n9728) );
  hi1s1 U9894 ( .DIN(n8054), .Q(n8062) );
  nnd2s1 U9895 ( .DIN1(n9744), .DIN2(n9758), .Q(n8054) );
  nnd4s1 U9896 ( .DIN1(n9759), .DIN2(n9760), .DIN3(n9761), .DIN4(n9762), 
        .Q(n9633) );
  nnd2s1 U9897 ( .DIN1(n8254), .DIN2(n9763), .Q(n9762) );
  nnd2s1 U9898 ( .DIN1(n8591), .DIN2(n7859), .Q(n9763) );
  hi1s1 U9899 ( .DIN(n8312), .Q(n8254) );
  nnd2s1 U9900 ( .DIN1(n9735), .DIN2(n9753), .Q(n8312) );
  nnd2s1 U9901 ( .DIN1(n8030), .DIN2(n9764), .Q(n9761) );
  nnd2s1 U9902 ( .DIN1(n7859), .DIN2(n8281), .Q(n9764) );
  nnd3s1 U9903 ( .DIN1(sa33[7]), .DIN2(n1428), .DIN3(n9758), .Q(n8281) );
  nnd2s1 U9904 ( .DIN1(n9737), .DIN2(n9758), .Q(n7859) );
  nor2s1 U9905 ( .DIN1(n1382), .DIN2(sa33[4]), .Q(n9758) );
  hi1s1 U9906 ( .DIN(n8318), .Q(n8030) );
  nnd2s1 U9907 ( .DIN1(n9736), .DIN2(n9745), .Q(n8318) );
  nor2s1 U9908 ( .DIN1(sa33[3]), .DIN2(sa33[1]), .Q(n9736) );
  nnd2s1 U9909 ( .DIN1(n7875), .DIN2(n9765), .Q(n9760) );
  nnd2s1 U9910 ( .DIN1(n8591), .DIN2(n8277), .Q(n9765) );
  nnd2s1 U9911 ( .DIN1(n9716), .DIN2(n9737), .Q(n8277) );
  nor2s1 U9912 ( .DIN1(n1428), .DIN2(sa33[7]), .Q(n9737) );
  nor2s1 U9913 ( .DIN1(sa33[5]), .DIN2(sa33[4]), .Q(n9716) );
  nnd3s1 U9914 ( .DIN1(sa33[4]), .DIN2(n1382), .DIN3(n9744), .Q(n8591) );
  nor2s1 U9915 ( .DIN1(sa33[7]), .DIN2(sa33[6]), .Q(n9744) );
  nnd2s1 U9916 ( .DIN1(n8257), .DIN2(n9766), .Q(n9759) );
  nnd2s1 U9917 ( .DIN1(n9100), .DIN2(n8076), .Q(n9766) );
  nnd2s1 U9918 ( .DIN1(n9753), .DIN2(n9745), .Q(n8076) );
  nor2s1 U9919 ( .DIN1(sa33[2]), .DIN2(sa33[0]), .Q(n9745) );
  and2s1 U9920 ( .DIN1(sa33[1]), .DIN2(sa33[3]), .Q(n9753) );
  nor2s1 U9921 ( .DIN1(n7866), .DIN2(n7875), .Q(n9100) );
  hi1s1 U9922 ( .DIN(n8590), .Q(n7875) );
  nnd2s1 U9923 ( .DIN1(n9735), .DIN2(n9709), .Q(n8590) );
  and2s1 U9924 ( .DIN1(sa33[2]), .DIN2(sa33[0]), .Q(n9735) );
  hi1s1 U9925 ( .DIN(n8259), .Q(n7866) );
  nnd2s1 U9926 ( .DIN1(n9727), .DIN2(n9709), .Q(n8259) );
  nor2s1 U9927 ( .DIN1(n1529), .DIN2(sa33[3]), .Q(n9709) );
  nor2s1 U9928 ( .DIN1(n1537), .DIN2(sa33[0]), .Q(n9727) );
  hi1s1 U9929 ( .DIN(n8032), .Q(n8257) );
  nnd3s1 U9930 ( .DIN1(n1382), .DIN2(n1428), .DIN3(n9732), .Q(n8032) );
  and2s1 U9931 ( .DIN1(sa33[7]), .DIN2(sa33[4]), .Q(n9732) );
  or3s1 U9932 ( .DIN1(n9767), .DIN2(n9768), .DIN3(n9769), .Q(n6115) );
  nnd4s1 U9933 ( .DIN1(n9472), .DIN2(n9770), .DIN3(n9309), .DIN4(n9771), 
        .Q(n9769) );
  and4s1 U9934 ( .DIN1(n9772), .DIN2(n9773), .DIN3(n9774), .DIN4(n8184), 
        .Q(n9771) );
  nnd2s1 U9935 ( .DIN1(n8197), .DIN2(n8001), .Q(n8184) );
  nnd2s1 U9936 ( .DIN1(n8224), .DIN2(n7983), .Q(n9774) );
  nnd2s1 U9937 ( .DIN1(n8005), .DIN2(n8187), .Q(n9773) );
  nor3s1 U9938 ( .DIN1(n9775), .DIN2(n9776), .DIN3(n9777), .Q(n9309) );
  nnd4s1 U9939 ( .DIN1(n9778), .DIN2(n9779), .DIN3(n9473), .DIN4(n9780), 
        .Q(n9777) );
  and3s1 U9940 ( .DIN1(n9781), .DIN2(n9782), .DIN3(n9783), .Q(n9780) );
  nnd2s1 U9941 ( .DIN1(n7997), .DIN2(n8187), .Q(n9783) );
  nnd2s1 U9942 ( .DIN1(n8197), .DIN2(n8492), .Q(n9782) );
  nnd2s1 U9943 ( .DIN1(n8213), .DIN2(n8196), .Q(n9781) );
  nor2s1 U9944 ( .DIN1(n9784), .DIN2(n9785), .Q(n9473) );
  nnd4s1 U9945 ( .DIN1(n9786), .DIN2(n9787), .DIN3(n9075), .DIN4(n9788), 
        .Q(n9785) );
  nnd2s1 U9946 ( .DIN1(n7984), .DIN2(n7993), .Q(n9788) );
  nnd2s1 U9947 ( .DIN1(n8564), .DIN2(n8540), .Q(n7993) );
  nnd2s1 U9948 ( .DIN1(n7997), .DIN2(n8963), .Q(n9075) );
  nnd2s1 U9949 ( .DIN1(n8519), .DIN2(n8493), .Q(n9787) );
  nnd2s1 U9950 ( .DIN1(n8187), .DIN2(n8001), .Q(n9786) );
  nnd4s1 U9951 ( .DIN1(n9789), .DIN2(n9790), .DIN3(n9791), .DIN4(n9792), 
        .Q(n9784) );
  nnd2s1 U9952 ( .DIN1(n8204), .DIN2(n9793), .Q(n9792) );
  nnd2s1 U9953 ( .DIN1(n8967), .DIN2(n8505), .Q(n9793) );
  nnd2s1 U9954 ( .DIN1(n8221), .DIN2(n9794), .Q(n9791) );
  nnd2s1 U9955 ( .DIN1(n8215), .DIN2(n8232), .Q(n9794) );
  nnd2s1 U9956 ( .DIN1(n8186), .DIN2(n9795), .Q(n9790) );
  nnd3s1 U9957 ( .DIN1(n8004), .DIN2(n8000), .DIN3(n7988), .Q(n9795) );
  nnd2s1 U9958 ( .DIN1(n8207), .DIN2(n9796), .Q(n9789) );
  nnd4s1 U9959 ( .DIN1(n8194), .DIN2(n8215), .DIN3(n8508), .DIN4(n8003), 
        .Q(n9796) );
  nnd3s1 U9960 ( .DIN1(n9797), .DIN2(n9798), .DIN3(n9051), .Q(n9776) );
  nnd2s1 U9961 ( .DIN1(n8186), .DIN2(n9026), .Q(n9051) );
  or2s1 U9962 ( .DIN1(n9025), .DIN2(n9059), .Q(n9798) );
  nor2s1 U9963 ( .DIN1(n8224), .DIN2(n8963), .Q(n9059) );
  nnd2s1 U9964 ( .DIN1(n8225), .DIN2(n8009), .Q(n9797) );
  nnd2s1 U9965 ( .DIN1(n8215), .DIN2(n7999), .Q(n8009) );
  nnd4s1 U9966 ( .DIN1(n9799), .DIN2(n9800), .DIN3(n9801), .DIN4(n9802), 
        .Q(n9775) );
  nnd2s1 U9967 ( .DIN1(n8493), .DIN2(n9325), .Q(n9802) );
  nnd2s1 U9968 ( .DIN1(n8539), .DIN2(n8237), .Q(n9325) );
  nnd2s1 U9969 ( .DIN1(n8005), .DIN2(n9803), .Q(n9801) );
  nnd2s1 U9970 ( .DIN1(n7999), .DIN2(n8232), .Q(n9803) );
  nnd2s1 U9971 ( .DIN1(n8185), .DIN2(n9804), .Q(n9800) );
  nnd2s1 U9972 ( .DIN1(n8212), .DIN2(n8237), .Q(n9804) );
  nnd2s1 U9973 ( .DIN1(n7992), .DIN2(n9805), .Q(n9799) );
  nnd2s1 U9974 ( .DIN1(n9067), .DIN2(n8958), .Q(n9805) );
  hi1s1 U9975 ( .DIN(n8223), .Q(n9067) );
  nnd2s1 U9976 ( .DIN1(n8535), .DIN2(n8236), .Q(n8223) );
  nor2s1 U9977 ( .DIN1(n9806), .DIN2(n9807), .Q(n9472) );
  nnd4s1 U9978 ( .DIN1(n9808), .DIN2(n9809), .DIN3(n9810), .DIN4(n9811), 
        .Q(n9807) );
  nnd2s1 U9979 ( .DIN1(n8198), .DIN2(n8527), .Q(n9811) );
  nnd2s1 U9980 ( .DIN1(n8212), .DIN2(n9025), .Q(n8527) );
  nnd2s1 U9981 ( .DIN1(n8494), .DIN2(n7982), .Q(n9810) );
  nnd2s1 U9982 ( .DIN1(n8005), .DIN2(n8185), .Q(n9809) );
  nnd2s1 U9983 ( .DIN1(n8233), .DIN2(n8518), .Q(n9808) );
  nnd4s1 U9984 ( .DIN1(n9812), .DIN2(n9813), .DIN3(n9814), .DIN4(n9815), 
        .Q(n9806) );
  nnd2s1 U9985 ( .DIN1(n7981), .DIN2(n9816), .Q(n9815) );
  or2s1 U9986 ( .DIN1(n9078), .DIN2(n8204), .Q(n9816) );
  nnd2s1 U9987 ( .DIN1(n8199), .DIN2(n9817), .Q(n9814) );
  nnd2s1 U9988 ( .DIN1(n7988), .DIN2(n8209), .Q(n9817) );
  nnd2s1 U9989 ( .DIN1(n8187), .DIN2(n9818), .Q(n9813) );
  nnd2s1 U9990 ( .DIN1(n8545), .DIN2(n8540), .Q(n9818) );
  nnd2s1 U9991 ( .DIN1(n7992), .DIN2(n9819), .Q(n9812) );
  nnd3s1 U9992 ( .DIN1(n8545), .DIN2(n8539), .DIN3(n9820), .Q(n9819) );
  nnd4s1 U9993 ( .DIN1(n8543), .DIN2(n9821), .DIN3(n9822), .DIN4(n9823), 
        .Q(n9768) );
  nnd2s1 U9994 ( .DIN1(n8492), .DIN2(n8494), .Q(n9823) );
  nnd2s1 U9995 ( .DIN1(n7982), .DIN2(n8963), .Q(n9822) );
  nnd2s1 U9996 ( .DIN1(n8204), .DIN2(n8198), .Q(n9821) );
  nnd2s1 U9997 ( .DIN1(n8207), .DIN2(n8196), .Q(n8543) );
  nnd4s1 U9998 ( .DIN1(n9824), .DIN2(n9825), .DIN3(n9826), .DIN4(n9827), 
        .Q(n9767) );
  nnd2s1 U9999 ( .DIN1(n8562), .DIN2(n9828), .Q(n9827) );
  nnd2s1 U10000 ( .DIN1(n9317), .DIN2(n8237), .Q(n9828) );
  nor2s1 U10001 ( .DIN1(n7997), .DIN2(n8001), .Q(n9317) );
  nnd2s1 U10002 ( .DIN1(n8213), .DIN2(n9829), .Q(n9826) );
  nnd2s1 U10003 ( .DIN1(n8500), .DIN2(n7990), .Q(n9829) );
  nnd2s1 U10004 ( .DIN1(n7992), .DIN2(n9830), .Q(n9825) );
  nnd2s1 U10005 ( .DIN1(n9025), .DIN2(n8540), .Q(n9830) );
  nnd2s1 U10006 ( .DIN1(n8230), .DIN2(n9046), .Q(n9824) );
  xor2s1 U10007 ( .DIN1(n5702), .DIN2(n5077), .Q(n7628) );
  nor4s1 U10008 ( .DIN1(n9831), .DIN2(n9832), .DIN3(n9833), .DIN4(n9834), 
        .Q(n5077) );
  nnd4s1 U10009 ( .DIN1(n8399), .DIN2(n9835), .DIN3(n9836), .DIN4(n9837), 
        .Q(n9834) );
  nnd2s1 U10010 ( .DIN1(n8129), .DIN2(n8934), .Q(n9837) );
  nnd2s1 U10011 ( .DIN1(n8453), .DIN2(n7838), .Q(n8934) );
  nnd2s1 U10012 ( .DIN1(n8170), .DIN2(n7840), .Q(n9836) );
  nnd2s1 U10013 ( .DIN1(n8149), .DIN2(n8422), .Q(n7840) );
  nnd2s1 U10014 ( .DIN1(n8883), .DIN2(n8140), .Q(n9835) );
  nnd2s1 U10015 ( .DIN1(n8163), .DIN2(n7820), .Q(n8399) );
  nnd4s1 U10016 ( .DIN1(n9838), .DIN2(n9839), .DIN3(n9840), .DIN4(n9841), 
        .Q(n9833) );
  nnd2s1 U10017 ( .DIN1(n7811), .DIN2(n9842), .Q(n9841) );
  nnd2s1 U10018 ( .DIN1(n7962), .DIN2(n8137), .Q(n9842) );
  nnd2s1 U10019 ( .DIN1(n8128), .DIN2(n9843), .Q(n9840) );
  nnd2s1 U10020 ( .DIN1(n8457), .DIN2(n8449), .Q(n9843) );
  or2s1 U10021 ( .DIN1(n8169), .DIN2(n8151), .Q(n9839) );
  nor2s1 U10022 ( .DIN1(n7831), .DIN2(n8140), .Q(n8151) );
  nnd2s1 U10023 ( .DIN1(n8433), .DIN2(n8161), .Q(n9838) );
  nnd2s1 U10024 ( .DIN1(n8146), .DIN2(n7961), .Q(n8161) );
  nnd3s1 U10025 ( .DIN1(n9269), .DIN2(n9277), .DIN3(n7802), .Q(n9832) );
  nor4s1 U10026 ( .DIN1(n9844), .DIN2(n9845), .DIN3(n9846), .DIN4(n9847), 
        .Q(n7802) );
  nnd4s1 U10027 ( .DIN1(n9848), .DIN2(n9849), .DIN3(n9850), .DIN4(n9851), 
        .Q(n9847) );
  nnd2s1 U10028 ( .DIN1(n7835), .DIN2(n7819), .Q(n9851) );
  nor2s1 U10029 ( .DIN1(n9852), .DIN2(n8853), .Q(n9850) );
  nor2s1 U10030 ( .DIN1(n8149), .DIN2(n7837), .Q(n8853) );
  nor2s1 U10031 ( .DIN1(n8137), .DIN2(n8173), .Q(n9852) );
  nnd2s1 U10032 ( .DIN1(n8160), .DIN2(n7818), .Q(n9849) );
  nnd2s1 U10033 ( .DIN1(n8129), .DIN2(n8147), .Q(n9848) );
  hi1s1 U10034 ( .DIN(n7833), .Q(n8129) );
  nnd3s1 U10035 ( .DIN1(n9853), .DIN2(n9854), .DIN3(n9855), .Q(n9846) );
  nnd2s1 U10036 ( .DIN1(n8140), .DIN2(n8440), .Q(n9855) );
  nnd2s1 U10037 ( .DIN1(n8146), .DIN2(n8137), .Q(n8440) );
  nnd2s1 U10038 ( .DIN1(n7820), .DIN2(n9856), .Q(n9854) );
  nnd3s1 U10039 ( .DIN1(n8450), .DIN2(n8818), .DIN3(n8457), .Q(n9856) );
  nnd2s1 U10040 ( .DIN1(n8139), .DIN2(n9857), .Q(n9853) );
  nnd3s1 U10041 ( .DIN1(n8452), .DIN2(n8817), .DIN3(n8420), .Q(n9857) );
  nor2s1 U10042 ( .DIN1(n8420), .DIN2(n8154), .Q(n9845) );
  nor2s1 U10043 ( .DIN1(n8924), .DIN2(n8419), .Q(n9844) );
  nor2s1 U10044 ( .DIN1(n7959), .DIN2(n7839), .Q(n8924) );
  and4s1 U10045 ( .DIN1(n9858), .DIN2(n9859), .DIN3(n9860), .DIN4(n9861), 
        .Q(n9277) );
  and4s1 U10046 ( .DIN1(n9862), .DIN2(n8867), .DIN3(n9863), .DIN4(n9864), 
        .Q(n9861) );
  nnd2s1 U10047 ( .DIN1(n8163), .DIN2(n8883), .Q(n9864) );
  nnd2s1 U10048 ( .DIN1(n7819), .DIN2(n7948), .Q(n9863) );
  nnd2s1 U10049 ( .DIN1(n7831), .DIN2(n8888), .Q(n8867) );
  nnd2s1 U10050 ( .DIN1(n7811), .DIN2(n7835), .Q(n9862) );
  and3s1 U10051 ( .DIN1(n9865), .DIN2(n9866), .DIN3(n9867), .Q(n9860) );
  nnd2s1 U10052 ( .DIN1(n8160), .DIN2(n9868), .Q(n9867) );
  nnd2s1 U10053 ( .DIN1(n7966), .DIN2(n8146), .Q(n9868) );
  nnd2s1 U10054 ( .DIN1(n7810), .DIN2(n9869), .Q(n9866) );
  nnd2s1 U10055 ( .DIN1(n7833), .DIN2(n7966), .Q(n9869) );
  nnd2s1 U10056 ( .DIN1(n8130), .DIN2(n8916), .Q(n9865) );
  nnd2s1 U10057 ( .DIN1(n8149), .DIN2(n8169), .Q(n8916) );
  nnd2s1 U10058 ( .DIN1(n7963), .DIN2(n9870), .Q(n9859) );
  nnd3s1 U10059 ( .DIN1(n8169), .DIN2(n7965), .DIN3(n7834), .Q(n9870) );
  hi1s1 U10060 ( .DIN(n7837), .Q(n7963) );
  or2s1 U10061 ( .DIN1(n8146), .DIN2(n9454), .Q(n9858) );
  nor2s1 U10062 ( .DIN1(n7821), .DIN2(n7839), .Q(n9454) );
  nor4s1 U10063 ( .DIN1(n9871), .DIN2(n9872), .DIN3(n9873), .DIN4(n9874), 
        .Q(n9269) );
  nnd4s1 U10064 ( .DIN1(n9875), .DIN2(n9876), .DIN3(n9877), .DIN4(n9878), 
        .Q(n9874) );
  nor2s1 U10065 ( .DIN1(n9879), .DIN2(n9880), .Q(n9878) );
  nor2s1 U10066 ( .DIN1(n8450), .DIN2(n7961), .Q(n9880) );
  nor2s1 U10067 ( .DIN1(n8452), .DIN2(n7966), .Q(n9879) );
  nnd2s1 U10068 ( .DIN1(n8147), .DIN2(n8409), .Q(n9877) );
  or2s1 U10069 ( .DIN1(n8854), .DIN2(n8414), .Q(n9876) );
  nor2s1 U10070 ( .DIN1(n7835), .DIN2(n8409), .Q(n8414) );
  nnd2s1 U10071 ( .DIN1(n7809), .DIN2(n7817), .Q(n9875) );
  nnd3s1 U10072 ( .DIN1(n9881), .DIN2(n9882), .DIN3(n9883), .Q(n9873) );
  nnd2s1 U10073 ( .DIN1(n7810), .DIN2(n8473), .Q(n9883) );
  nnd2s1 U10074 ( .DIN1(n7961), .DIN2(n8422), .Q(n8473) );
  hi1s1 U10075 ( .DIN(n8173), .Q(n7810) );
  nnd2s1 U10076 ( .DIN1(n7948), .DIN2(n9884), .Q(n9882) );
  nnd2s1 U10077 ( .DIN1(n8817), .DIN2(n8152), .Q(n9884) );
  nnd2s1 U10078 ( .DIN1(n8139), .DIN2(n9885), .Q(n9881) );
  nnd2s1 U10079 ( .DIN1(n7830), .DIN2(n8854), .Q(n9885) );
  nor2s1 U10080 ( .DIN1(n9886), .DIN2(n7834), .Q(n9872) );
  nor2s1 U10081 ( .DIN1(n7811), .DIN2(n8130), .Q(n9886) );
  nor2s1 U10082 ( .DIN1(n9887), .DIN2(n7952), .Q(n9871) );
  nor2s1 U10083 ( .DIN1(n7817), .DIN2(n7959), .Q(n9887) );
  nnd4s1 U10084 ( .DIN1(n9411), .DIN2(n9888), .DIN3(n9889), .DIN4(n9890), 
        .Q(n9831) );
  nnd2s1 U10085 ( .DIN1(n7809), .DIN2(n8147), .Q(n9890) );
  nnd2s1 U10086 ( .DIN1(n8130), .DIN2(n7835), .Q(n9889) );
  nnd2s1 U10087 ( .DIN1(n8432), .DIN2(n8160), .Q(n9888) );
  nor3s1 U10088 ( .DIN1(n9891), .DIN2(n9892), .DIN3(n9893), .Q(n9411) );
  nnd4s1 U10089 ( .DIN1(n7805), .DIN2(n9278), .DIN3(n9273), .DIN4(n9894), 
        .Q(n9893) );
  and3s1 U10090 ( .DIN1(n9895), .DIN2(n9896), .DIN3(n9897), .Q(n9894) );
  nnd2s1 U10091 ( .DIN1(n8128), .DIN2(n8160), .Q(n9897) );
  nnd2s1 U10092 ( .DIN1(n7812), .DIN2(n8147), .Q(n9896) );
  hi1s1 U10093 ( .DIN(n8449), .Q(n8147) );
  hi1s1 U10094 ( .DIN(n7966), .Q(n7812) );
  nnd2s1 U10095 ( .DIN1(n8433), .DIN2(n7827), .Q(n9895) );
  hi1s1 U10096 ( .DIN(n8154), .Q(n7827) );
  and4s1 U10097 ( .DIN1(n9898), .DIN2(n9899), .DIN3(n9900), .DIN4(n9901), 
        .Q(n9273) );
  and4s1 U10098 ( .DIN1(n9902), .DIN2(n9903), .DIN3(n8832), .DIN4(n8407), 
        .Q(n9901) );
  nnd2s1 U10099 ( .DIN1(n7821), .DIN2(n7948), .Q(n8407) );
  nnd2s1 U10100 ( .DIN1(n8130), .DIN2(n7809), .Q(n8832) );
  nnd2s1 U10101 ( .DIN1(n7959), .DIN2(n7835), .Q(n9903) );
  nnd2s1 U10102 ( .DIN1(n8128), .DIN2(n8433), .Q(n9902) );
  and3s1 U10103 ( .DIN1(n9904), .DIN2(n9905), .DIN3(n9906), .Q(n9900) );
  nnd2s1 U10104 ( .DIN1(n7822), .DIN2(n9423), .Q(n9906) );
  nnd2s1 U10105 ( .DIN1(n8418), .DIN2(n8173), .Q(n9423) );
  nnd2s1 U10106 ( .DIN1(n7819), .DIN2(n9907), .Q(n9905) );
  nnd2s1 U10107 ( .DIN1(n8861), .DIN2(n8154), .Q(n9907) );
  nor2s1 U10108 ( .DIN1(n8432), .DIN2(n8409), .Q(n8861) );
  hi1s1 U10109 ( .DIN(n8149), .Q(n8409) );
  nnd2s1 U10110 ( .DIN1(n8888), .DIN2(n9908), .Q(n9904) );
  nnd2s1 U10111 ( .DIN1(n8453), .DIN2(n7837), .Q(n9908) );
  nnd2s1 U10112 ( .DIN1(n8432), .DIN2(n9909), .Q(n9899) );
  nnd2s1 U10113 ( .DIN1(n8475), .DIN2(n7830), .Q(n9909) );
  nnd2s1 U10114 ( .DIN1(n8140), .DIN2(n9910), .Q(n9898) );
  nnd3s1 U10115 ( .DIN1(n7962), .DIN2(n7834), .DIN3(n7966), .Q(n9910) );
  and4s1 U10116 ( .DIN1(n9911), .DIN2(n9912), .DIN3(n9913), .DIN4(n9914), 
        .Q(n9278) );
  nor4s1 U10117 ( .DIN1(n9915), .DIN2(n9916), .DIN3(n9917), .DIN4(n9918), 
        .Q(n9914) );
  nor2s1 U10118 ( .DIN1(n9919), .DIN2(n7961), .Q(n9918) );
  nor2s1 U10119 ( .DIN1(n8130), .DIN2(n8160), .Q(n9919) );
  nor2s1 U10120 ( .DIN1(n9920), .DIN2(n8422), .Q(n9917) );
  nor2s1 U10121 ( .DIN1(n7817), .DIN2(n7821), .Q(n9920) );
  hi1s1 U10122 ( .DIN(n7830), .Q(n7821) );
  nnd3s1 U10123 ( .DIN1(n9921), .DIN2(n1362), .DIN3(sa11[1]), .Q(n7830) );
  nor2s1 U10124 ( .DIN1(n9922), .DIN2(n8173), .Q(n9916) );
  nor2s1 U10125 ( .DIN1(n7947), .DIN2(n8432), .Q(n9922) );
  nnd3s1 U10126 ( .DIN1(n9923), .DIN2(n9924), .DIN3(n9925), .Q(n9915) );
  nnd2s1 U10127 ( .DIN1(n7817), .DIN2(n8883), .Q(n9925) );
  nnd2s1 U10128 ( .DIN1(n7818), .DIN2(n9926), .Q(n9924) );
  nnd2s1 U10129 ( .DIN1(n8152), .DIN2(n8420), .Q(n9926) );
  nnd2s1 U10130 ( .DIN1(n7831), .DIN2(n9303), .Q(n9923) );
  nnd2s1 U10131 ( .DIN1(n8146), .DIN2(n8149), .Q(n9303) );
  nnd2s1 U10132 ( .DIN1(n9927), .DIN2(n9928), .Q(n8149) );
  hi1s1 U10133 ( .DIN(n8457), .Q(n7831) );
  and3s1 U10134 ( .DIN1(n9929), .DIN2(n9930), .DIN3(n9931), .Q(n9913) );
  nnd2s1 U10135 ( .DIN1(n8170), .DIN2(n8139), .Q(n9931) );
  hi1s1 U10136 ( .DIN(n7962), .Q(n8139) );
  nnd2s1 U10137 ( .DIN1(n7947), .DIN2(n8163), .Q(n9930) );
  nnd2s1 U10138 ( .DIN1(n7822), .DIN2(n7839), .Q(n9929) );
  nnd2s1 U10139 ( .DIN1(n7959), .DIN2(n7809), .Q(n9912) );
  nnd2s1 U10140 ( .DIN1(n7835), .DIN2(n8140), .Q(n9911) );
  hi1s1 U10141 ( .DIN(n8450), .Q(n8140) );
  hi1s1 U10142 ( .DIN(n8878), .Q(n7835) );
  nnd2s1 U10143 ( .DIN1(n9927), .DIN2(n9932), .Q(n8878) );
  nor4s1 U10144 ( .DIN1(n9933), .DIN2(n9934), .DIN3(n9935), .DIN4(n9936), 
        .Q(n7805) );
  nnd4s1 U10145 ( .DIN1(n9937), .DIN2(n9938), .DIN3(n9939), .DIN4(n9940), 
        .Q(n9936) );
  nnd2s1 U10146 ( .DIN1(n8163), .DIN2(n7818), .Q(n9940) );
  hi1s1 U10147 ( .DIN(n8854), .Q(n8163) );
  nnd2s1 U10148 ( .DIN1(n7811), .DIN2(n7820), .Q(n9939) );
  hi1s1 U10149 ( .DIN(n8422), .Q(n7820) );
  nnd2s1 U10150 ( .DIN1(n9941), .DIN2(n9928), .Q(n8422) );
  hi1s1 U10151 ( .DIN(n8418), .Q(n7811) );
  nnd3s1 U10152 ( .DIN1(n1362), .DIN2(n1429), .DIN3(n9921), .Q(n8418) );
  nnd2s1 U10153 ( .DIN1(n7947), .DIN2(n7839), .Q(n9938) );
  hi1s1 U10154 ( .DIN(n8420), .Q(n7839) );
  hi1s1 U10155 ( .DIN(n8169), .Q(n7947) );
  nnd2s1 U10156 ( .DIN1(n7809), .DIN2(n7819), .Q(n9937) );
  hi1s1 U10157 ( .DIN(n8146), .Q(n7809) );
  nnd2s1 U10158 ( .DIN1(n9942), .DIN2(n9943), .Q(n8146) );
  nnd3s1 U10159 ( .DIN1(n9944), .DIN2(n9945), .DIN3(n9946), .Q(n9935) );
  nnd2s1 U10160 ( .DIN1(n8128), .DIN2(n9947), .Q(n9946) );
  nnd3s1 U10161 ( .DIN1(n8173), .DIN2(n8450), .DIN3(n8420), .Q(n9947) );
  nnd3s1 U10162 ( .DIN1(n9948), .DIN2(n1443), .DIN3(sa11[0]), .Q(n8420) );
  nnd3s1 U10163 ( .DIN1(sa11[0]), .DIN2(n1429), .DIN3(n9949), .Q(n8173) );
  hi1s1 U10164 ( .DIN(n8825), .Q(n8128) );
  nnd2s1 U10165 ( .DIN1(n7822), .DIN2(n9950), .Q(n9945) );
  nnd2s1 U10166 ( .DIN1(n8449), .DIN2(n8854), .Q(n9950) );
  nnd3s1 U10167 ( .DIN1(n1362), .DIN2(n1429), .DIN3(n9949), .Q(n8449) );
  hi1s1 U10168 ( .DIN(n7952), .Q(n7822) );
  nnd2s1 U10169 ( .DIN1(n8160), .DIN2(n9951), .Q(n9944) );
  nnd2s1 U10170 ( .DIN1(n7833), .DIN2(n8419), .Q(n9951) );
  nnd2s1 U10171 ( .DIN1(n9942), .DIN2(n9928), .Q(n7833) );
  hi1s1 U10172 ( .DIN(n8817), .Q(n8160) );
  nnd3s1 U10173 ( .DIN1(sa11[0]), .DIN2(n1429), .DIN3(n9921), .Q(n8817) );
  nor2s1 U10174 ( .DIN1(n8154), .DIN2(n7838), .Q(n9934) );
  nnd2s1 U10175 ( .DIN1(n9927), .DIN2(n9952), .Q(n8154) );
  and2s1 U10176 ( .DIN1(n8433), .DIN2(n9953), .Q(n9933) );
  nnd4s1 U10177 ( .DIN1(n7966), .DIN2(n7962), .DIN3(n8169), .DIN4(n7965), 
        .Q(n9953) );
  nnd2s1 U10178 ( .DIN1(n9943), .DIN2(n9954), .Q(n8169) );
  nnd2s1 U10179 ( .DIN1(n9954), .DIN2(n9928), .Q(n7962) );
  nor2s1 U10180 ( .DIN1(n1518), .DIN2(n1400), .Q(n9928) );
  nnd2s1 U10181 ( .DIN1(n9952), .DIN2(n9941), .Q(n7966) );
  hi1s1 U10182 ( .DIN(n8152), .Q(n8433) );
  nnd3s1 U10183 ( .DIN1(sa11[1]), .DIN2(n1362), .DIN3(n9949), .Q(n8152) );
  nnd3s1 U10184 ( .DIN1(n9955), .DIN2(n9956), .DIN3(n9957), .Q(n9892) );
  nnd2s1 U10185 ( .DIN1(n7959), .DIN2(n7818), .Q(n9957) );
  hi1s1 U10186 ( .DIN(n7834), .Q(n7818) );
  hi1s1 U10187 ( .DIN(n8475), .Q(n7959) );
  nnd3s1 U10188 ( .DIN1(sa11[2]), .DIN2(n1362), .DIN3(n9958), .Q(n8475) );
  nnd2s1 U10189 ( .DIN1(n8888), .DIN2(n7817), .Q(n9956) );
  hi1s1 U10190 ( .DIN(n7838), .Q(n7817) );
  nnd3s1 U10191 ( .DIN1(sa11[1]), .DIN2(sa11[0]), .DIN3(n9949), .Q(n7838) );
  and2s1 U10192 ( .DIN1(sa11[3]), .DIN2(sa11[2]), .Q(n9949) );
  hi1s1 U10193 ( .DIN(n7961), .Q(n8888) );
  nnd2s1 U10194 ( .DIN1(n8130), .DIN2(n7948), .Q(n9955) );
  hi1s1 U10195 ( .DIN(n8137), .Q(n7948) );
  nnd2s1 U10196 ( .DIN1(n9952), .DIN2(n9954), .Q(n8137) );
  hi1s1 U10197 ( .DIN(n8818), .Q(n8130) );
  nnd4s1 U10198 ( .DIN1(n9959), .DIN2(n9960), .DIN3(n9961), .DIN4(n9962), 
        .Q(n9891) );
  nnd2s1 U10199 ( .DIN1(n8883), .DIN2(n9963), .Q(n9962) );
  nnd2s1 U10200 ( .DIN1(n8457), .DIN2(n7837), .Q(n9963) );
  nnd3s1 U10201 ( .DIN1(sa11[2]), .DIN2(sa11[0]), .DIN3(n9958), .Q(n7837) );
  hi1s1 U10202 ( .DIN(n8419), .Q(n8883) );
  nnd2s1 U10203 ( .DIN1(n9932), .DIN2(n9954), .Q(n8419) );
  and2s1 U10204 ( .DIN1(sa11[4]), .DIN2(sa11[6]), .Q(n9954) );
  nnd2s1 U10205 ( .DIN1(n8432), .DIN2(n9964), .Q(n9961) );
  nnd4s1 U10206 ( .DIN1(n8457), .DIN2(n8854), .DIN3(n8450), .DIN4(n8818), 
        .Q(n9964) );
  nnd3s1 U10207 ( .DIN1(sa11[0]), .DIN2(n9948), .DIN3(sa11[2]), .Q(n8818) );
  nnd3s1 U10208 ( .DIN1(n9921), .DIN2(sa11[0]), .DIN3(sa11[1]), .Q(n8450) );
  and2s1 U10209 ( .DIN1(sa11[3]), .DIN2(n1443), .Q(n9921) );
  nnd3s1 U10210 ( .DIN1(sa11[0]), .DIN2(n1443), .DIN3(n9958), .Q(n8854) );
  nnd3s1 U10211 ( .DIN1(n1362), .DIN2(n1443), .DIN3(n9948), .Q(n8457) );
  hi1s1 U10212 ( .DIN(n7965), .Q(n8432) );
  nnd2s1 U10213 ( .DIN1(n9932), .DIN2(n9942), .Q(n7965) );
  nnd2s1 U10214 ( .DIN1(n8170), .DIN2(n8858), .Q(n9960) );
  nnd2s1 U10215 ( .DIN1(n8825), .DIN2(n7834), .Q(n8858) );
  nnd2s1 U10216 ( .DIN1(n9943), .DIN2(n9941), .Q(n7834) );
  nnd2s1 U10217 ( .DIN1(n9932), .DIN2(n9941), .Q(n8825) );
  and2s1 U10218 ( .DIN1(sa11[6]), .DIN2(n1530), .Q(n9941) );
  nor2s1 U10219 ( .DIN1(sa11[7]), .DIN2(sa11[5]), .Q(n9932) );
  hi1s1 U10220 ( .DIN(n8453), .Q(n8170) );
  nnd3s1 U10221 ( .DIN1(n9948), .DIN2(n1362), .DIN3(sa11[2]), .Q(n8453) );
  nor2s1 U10222 ( .DIN1(sa11[3]), .DIN2(sa11[1]), .Q(n9948) );
  nnd2s1 U10223 ( .DIN1(n7819), .DIN2(n8442), .Q(n9959) );
  nnd2s1 U10224 ( .DIN1(n7952), .DIN2(n7961), .Q(n8442) );
  nnd2s1 U10225 ( .DIN1(n9942), .DIN2(n9952), .Q(n7961) );
  nor2s1 U10226 ( .DIN1(n1518), .DIN2(sa11[5]), .Q(n9952) );
  nor2s1 U10227 ( .DIN1(sa11[6]), .DIN2(sa11[4]), .Q(n9942) );
  nnd2s1 U10228 ( .DIN1(n9927), .DIN2(n9943), .Q(n7952) );
  nor2s1 U10229 ( .DIN1(n1400), .DIN2(sa11[7]), .Q(n9943) );
  nor2s1 U10230 ( .DIN1(n1530), .DIN2(sa11[6]), .Q(n9927) );
  hi1s1 U10231 ( .DIN(n8452), .Q(n7819) );
  nnd3s1 U10232 ( .DIN1(n1362), .DIN2(n1443), .DIN3(n9958), .Q(n8452) );
  nor2s1 U10233 ( .DIN1(n1429), .DIN2(sa11[3]), .Q(n9958) );
  hi1s1 U10234 ( .DIN(n9406), .Q(n5702) );
  or4s1 U10235 ( .DIN1(n9965), .DIN2(n9966), .DIN3(n9967), .DIN4(n9968), 
        .Q(n9406) );
  nnd4s1 U10236 ( .DIN1(n8482), .DIN2(n9969), .DIN3(n9970), .DIN4(n9971), 
        .Q(n9968) );
  nnd2s1 U10237 ( .DIN1(n8185), .DIN2(n9078), .Q(n9971) );
  nnd2s1 U10238 ( .DIN1(n8539), .DIN2(n8540), .Q(n9078) );
  nnd2s1 U10239 ( .DIN1(n8233), .DIN2(n9046), .Q(n9970) );
  nnd2s1 U10240 ( .DIN1(n8209), .DIN2(n8508), .Q(n9046) );
  nnd2s1 U10241 ( .DIN1(n9026), .DIN2(n8199), .Q(n9969) );
  nnd2s1 U10242 ( .DIN1(n8225), .DIN2(n8963), .Q(n8482) );
  nnd4s1 U10243 ( .DIN1(n9972), .DIN2(n9973), .DIN3(n9974), .DIN4(n9975), 
        .Q(n9967) );
  nnd2s1 U10244 ( .DIN1(n8005), .DIN2(n9976), .Q(n9975) );
  nnd2s1 U10245 ( .DIN1(n8000), .DIN2(n8194), .Q(n9976) );
  nnd2s1 U10246 ( .DIN1(n8197), .DIN2(n9977), .Q(n9974) );
  nnd2s1 U10247 ( .DIN1(n8545), .DIN2(n8535), .Q(n9977) );
  or2s1 U10248 ( .DIN1(n8232), .DIN2(n8211), .Q(n9973) );
  nor2s1 U10249 ( .DIN1(n8213), .DIN2(n8199), .Q(n8211) );
  nnd2s1 U10250 ( .DIN1(n8519), .DIN2(n8222), .Q(n9972) );
  nnd2s1 U10251 ( .DIN1(n8206), .DIN2(n7999), .Q(n8222) );
  nnd3s1 U10252 ( .DIN1(n9308), .DIN2(n9778), .DIN3(n9770), .Q(n9966) );
  nor4s1 U10253 ( .DIN1(n9978), .DIN2(n9979), .DIN3(n9980), .DIN4(n9981), 
        .Q(n9770) );
  nnd4s1 U10254 ( .DIN1(n9982), .DIN2(n9983), .DIN3(n9984), .DIN4(n9985), 
        .Q(n9981) );
  nnd2s1 U10255 ( .DIN1(n7992), .DIN2(n7982), .Q(n9985) );
  nor2s1 U10256 ( .DIN1(n9986), .DIN2(n8995), .Q(n9984) );
  nor2s1 U10257 ( .DIN1(n8209), .DIN2(n9025), .Q(n8995) );
  nor2s1 U10258 ( .DIN1(n8194), .DIN2(n8236), .Q(n9986) );
  nnd2s1 U10259 ( .DIN1(n8221), .DIN2(n8494), .Q(n9983) );
  nnd2s1 U10260 ( .DIN1(n8185), .DIN2(n8207), .Q(n9982) );
  hi1s1 U10261 ( .DIN(n8500), .Q(n8185) );
  nnd3s1 U10262 ( .DIN1(n9987), .DIN2(n9988), .DIN3(n9989), .Q(n9980) );
  nnd2s1 U10263 ( .DIN1(n8199), .DIN2(n8526), .Q(n9989) );
  nnd2s1 U10264 ( .DIN1(n8206), .DIN2(n8194), .Q(n8526) );
  nnd2s1 U10265 ( .DIN1(n8963), .DIN2(n9990), .Q(n9988) );
  nnd3s1 U10266 ( .DIN1(n8536), .DIN2(n8959), .DIN3(n8545), .Q(n9990) );
  nnd2s1 U10267 ( .DIN1(n8196), .DIN2(n9991), .Q(n9987) );
  nnd3s1 U10268 ( .DIN1(n8538), .DIN2(n8958), .DIN3(n8506), .Q(n9991) );
  nor2s1 U10269 ( .DIN1(n8506), .DIN2(n8215), .Q(n9979) );
  nor2s1 U10270 ( .DIN1(n9068), .DIN2(n8505), .Q(n9978) );
  nor2s1 U10271 ( .DIN1(n7997), .DIN2(n8230), .Q(n9068) );
  and4s1 U10272 ( .DIN1(n9992), .DIN2(n9993), .DIN3(n9994), .DIN4(n9995), 
        .Q(n9778) );
  and4s1 U10273 ( .DIN1(n9996), .DIN2(n9009), .DIN3(n9997), .DIN4(n9998), 
        .Q(n9995) );
  nnd2s1 U10274 ( .DIN1(n8225), .DIN2(n9026), .Q(n9998) );
  nnd2s1 U10275 ( .DIN1(n7982), .DIN2(n7984), .Q(n9997) );
  nnd2s1 U10276 ( .DIN1(n8213), .DIN2(n9031), .Q(n9009) );
  nnd2s1 U10277 ( .DIN1(n8005), .DIN2(n7992), .Q(n9996) );
  and3s1 U10278 ( .DIN1(n9999), .DIN2(n10000), .DIN3(n10001), .Q(n9994) );
  nnd2s1 U10279 ( .DIN1(n8221), .DIN2(n10002), .Q(n10001) );
  nnd2s1 U10280 ( .DIN1(n8004), .DIN2(n8206), .Q(n10002) );
  nnd2s1 U10281 ( .DIN1(n7983), .DIN2(n10003), .Q(n10000) );
  nnd2s1 U10282 ( .DIN1(n8500), .DIN2(n8004), .Q(n10003) );
  nnd2s1 U10283 ( .DIN1(n8186), .DIN2(n9060), .Q(n9999) );
  nnd2s1 U10284 ( .DIN1(n8209), .DIN2(n8232), .Q(n9060) );
  nnd2s1 U10285 ( .DIN1(n8001), .DIN2(n10004), .Q(n9993) );
  nnd3s1 U10286 ( .DIN1(n8232), .DIN2(n8003), .DIN3(n7990), .Q(n10004) );
  hi1s1 U10287 ( .DIN(n9025), .Q(n8001) );
  or2s1 U10288 ( .DIN1(n8206), .DIN2(n9820), .Q(n9992) );
  nor2s1 U10289 ( .DIN1(n8204), .DIN2(n8230), .Q(n9820) );
  nor4s1 U10290 ( .DIN1(n10005), .DIN2(n10006), .DIN3(n10007), .DIN4(n10008), 
        .Q(n9308) );
  nnd4s1 U10291 ( .DIN1(n10009), .DIN2(n10010), .DIN3(n10011), .DIN4(n10012), 
        .Q(n10008) );
  nor2s1 U10292 ( .DIN1(n10013), .DIN2(n10014), .Q(n10012) );
  nor2s1 U10293 ( .DIN1(n8536), .DIN2(n7999), .Q(n10014) );
  nor2s1 U10294 ( .DIN1(n8538), .DIN2(n8004), .Q(n10013) );
  nnd2s1 U10295 ( .DIN1(n8207), .DIN2(n8493), .Q(n10011) );
  or2s1 U10296 ( .DIN1(n8996), .DIN2(n8499), .Q(n10010) );
  nor2s1 U10297 ( .DIN1(n7992), .DIN2(n8493), .Q(n8499) );
  nnd2s1 U10298 ( .DIN1(n8224), .DIN2(n8492), .Q(n10009) );
  nnd3s1 U10299 ( .DIN1(n10015), .DIN2(n10016), .DIN3(n10017), .Q(n10007) );
  nnd2s1 U10300 ( .DIN1(n7983), .DIN2(n8561), .Q(n10017) );
  nnd2s1 U10301 ( .DIN1(n7999), .DIN2(n8508), .Q(n8561) );
  hi1s1 U10302 ( .DIN(n8236), .Q(n7983) );
  nnd2s1 U10303 ( .DIN1(n7984), .DIN2(n10018), .Q(n10016) );
  nnd2s1 U10304 ( .DIN1(n8958), .DIN2(n8212), .Q(n10018) );
  nnd2s1 U10305 ( .DIN1(n8196), .DIN2(n10019), .Q(n10015) );
  nnd2s1 U10306 ( .DIN1(n8237), .DIN2(n8996), .Q(n10019) );
  nor2s1 U10307 ( .DIN1(n10020), .DIN2(n7990), .Q(n10006) );
  nor2s1 U10308 ( .DIN1(n8005), .DIN2(n8186), .Q(n10020) );
  nor2s1 U10309 ( .DIN1(n10021), .DIN2(n7988), .Q(n10005) );
  nor2s1 U10310 ( .DIN1(n8492), .DIN2(n7997), .Q(n10021) );
  nnd4s1 U10311 ( .DIN1(n9470), .DIN2(n10022), .DIN3(n10023), .DIN4(n10024), 
        .Q(n9965) );
  nnd2s1 U10312 ( .DIN1(n8224), .DIN2(n8207), .Q(n10024) );
  nnd2s1 U10313 ( .DIN1(n8186), .DIN2(n7992), .Q(n10023) );
  nnd2s1 U10314 ( .DIN1(n8518), .DIN2(n8221), .Q(n10022) );
  nor3s1 U10315 ( .DIN1(n10025), .DIN2(n10026), .DIN3(n10027), .Q(n9470) );
  nnd4s1 U10316 ( .DIN1(n9772), .DIN2(n9779), .DIN3(n9313), .DIN4(n10028), 
        .Q(n10027) );
  and3s1 U10317 ( .DIN1(n10029), .DIN2(n10030), .DIN3(n10031), .Q(n10028) );
  nnd2s1 U10318 ( .DIN1(n8197), .DIN2(n8221), .Q(n10031) );
  nnd2s1 U10319 ( .DIN1(n8187), .DIN2(n8207), .Q(n10030) );
  hi1s1 U10320 ( .DIN(n8535), .Q(n8207) );
  hi1s1 U10321 ( .DIN(n8004), .Q(n8187) );
  nnd2s1 U10322 ( .DIN1(n8519), .DIN2(n8562), .Q(n10029) );
  hi1s1 U10323 ( .DIN(n8215), .Q(n8562) );
  and4s1 U10324 ( .DIN1(n10032), .DIN2(n10033), .DIN3(n10034), .DIN4(n10035), 
        .Q(n9313) );
  and4s1 U10325 ( .DIN1(n10036), .DIN2(n10037), .DIN3(n8974), .DIN4(n8490), 
        .Q(n10035) );
  nnd2s1 U10326 ( .DIN1(n8204), .DIN2(n7984), .Q(n8490) );
  nnd2s1 U10327 ( .DIN1(n8186), .DIN2(n8224), .Q(n8974) );
  nnd2s1 U10328 ( .DIN1(n7997), .DIN2(n7992), .Q(n10037) );
  nnd2s1 U10329 ( .DIN1(n8197), .DIN2(n8519), .Q(n10036) );
  and3s1 U10330 ( .DIN1(n10038), .DIN2(n10039), .DIN3(n10040), .Q(n10034) );
  nnd2s1 U10331 ( .DIN1(n8198), .DIN2(n9484), .Q(n10040) );
  nnd2s1 U10332 ( .DIN1(n8504), .DIN2(n8236), .Q(n9484) );
  nnd2s1 U10333 ( .DIN1(n7982), .DIN2(n10041), .Q(n10039) );
  nnd2s1 U10334 ( .DIN1(n9003), .DIN2(n8215), .Q(n10041) );
  nor2s1 U10335 ( .DIN1(n8518), .DIN2(n8493), .Q(n9003) );
  hi1s1 U10336 ( .DIN(n8209), .Q(n8493) );
  nnd2s1 U10337 ( .DIN1(n9031), .DIN2(n10042), .Q(n10038) );
  nnd2s1 U10338 ( .DIN1(n8539), .DIN2(n9025), .Q(n10042) );
  nnd2s1 U10339 ( .DIN1(n8518), .DIN2(n10043), .Q(n10033) );
  nnd2s1 U10340 ( .DIN1(n8564), .DIN2(n8237), .Q(n10043) );
  nnd2s1 U10341 ( .DIN1(n8199), .DIN2(n10044), .Q(n10032) );
  nnd3s1 U10342 ( .DIN1(n8000), .DIN2(n7990), .DIN3(n8004), .Q(n10044) );
  and4s1 U10343 ( .DIN1(n10045), .DIN2(n10046), .DIN3(n10047), .DIN4(n10048), 
        .Q(n9779) );
  nor4s1 U10344 ( .DIN1(n10049), .DIN2(n10050), .DIN3(n10051), .DIN4(n10052), 
        .Q(n10048) );
  nor2s1 U10345 ( .DIN1(n10053), .DIN2(n7999), .Q(n10052) );
  nor2s1 U10346 ( .DIN1(n8186), .DIN2(n8221), .Q(n10053) );
  nor2s1 U10347 ( .DIN1(n10054), .DIN2(n8508), .Q(n10051) );
  nor2s1 U10348 ( .DIN1(n8492), .DIN2(n8204), .Q(n10054) );
  hi1s1 U10349 ( .DIN(n8237), .Q(n8204) );
  nnd3s1 U10350 ( .DIN1(n10055), .DIN2(n1363), .DIN3(sa00[1]), .Q(n8237) );
  nor2s1 U10351 ( .DIN1(n10056), .DIN2(n8236), .Q(n10050) );
  nor2s1 U10352 ( .DIN1(n7981), .DIN2(n8518), .Q(n10056) );
  nnd3s1 U10353 ( .DIN1(n10057), .DIN2(n10058), .DIN3(n10059), .Q(n10049) );
  nnd2s1 U10354 ( .DIN1(n8492), .DIN2(n9026), .Q(n10059) );
  nnd2s1 U10355 ( .DIN1(n8494), .DIN2(n10060), .Q(n10058) );
  nnd2s1 U10356 ( .DIN1(n8212), .DIN2(n8506), .Q(n10060) );
  nnd2s1 U10357 ( .DIN1(n8213), .DIN2(n9324), .Q(n10057) );
  nnd2s1 U10358 ( .DIN1(n8206), .DIN2(n8209), .Q(n9324) );
  nnd2s1 U10359 ( .DIN1(n10061), .DIN2(n10062), .Q(n8209) );
  hi1s1 U10360 ( .DIN(n8545), .Q(n8213) );
  and3s1 U10361 ( .DIN1(n10063), .DIN2(n10064), .DIN3(n10065), .Q(n10047) );
  nnd2s1 U10362 ( .DIN1(n8233), .DIN2(n8196), .Q(n10065) );
  hi1s1 U10363 ( .DIN(n8000), .Q(n8196) );
  nnd2s1 U10364 ( .DIN1(n7981), .DIN2(n8225), .Q(n10064) );
  nnd2s1 U10365 ( .DIN1(n8198), .DIN2(n8230), .Q(n10063) );
  nnd2s1 U10366 ( .DIN1(n7997), .DIN2(n8224), .Q(n10046) );
  nnd2s1 U10367 ( .DIN1(n7992), .DIN2(n8199), .Q(n10045) );
  hi1s1 U10368 ( .DIN(n8536), .Q(n8199) );
  hi1s1 U10369 ( .DIN(n9020), .Q(n7992) );
  nnd2s1 U10370 ( .DIN1(n10061), .DIN2(n10066), .Q(n9020) );
  nor4s1 U10371 ( .DIN1(n10067), .DIN2(n10068), .DIN3(n10069), .DIN4(n10070), 
        .Q(n9772) );
  nnd4s1 U10372 ( .DIN1(n10071), .DIN2(n10072), .DIN3(n10073), .DIN4(n10074), 
        .Q(n10070) );
  nnd2s1 U10373 ( .DIN1(n8225), .DIN2(n8494), .Q(n10074) );
  hi1s1 U10374 ( .DIN(n8996), .Q(n8225) );
  nnd2s1 U10375 ( .DIN1(n8005), .DIN2(n8963), .Q(n10073) );
  hi1s1 U10376 ( .DIN(n8508), .Q(n8963) );
  nnd2s1 U10377 ( .DIN1(n10075), .DIN2(n10062), .Q(n8508) );
  hi1s1 U10378 ( .DIN(n8504), .Q(n8005) );
  nnd3s1 U10379 ( .DIN1(n1363), .DIN2(n1430), .DIN3(n10055), .Q(n8504) );
  nnd2s1 U10380 ( .DIN1(n7981), .DIN2(n8230), .Q(n10072) );
  hi1s1 U10381 ( .DIN(n8506), .Q(n8230) );
  hi1s1 U10382 ( .DIN(n8232), .Q(n7981) );
  nnd2s1 U10383 ( .DIN1(n8224), .DIN2(n7982), .Q(n10071) );
  hi1s1 U10384 ( .DIN(n8206), .Q(n8224) );
  nnd2s1 U10385 ( .DIN1(n10076), .DIN2(n10077), .Q(n8206) );
  nnd3s1 U10386 ( .DIN1(n10078), .DIN2(n10079), .DIN3(n10080), .Q(n10069) );
  nnd2s1 U10387 ( .DIN1(n8197), .DIN2(n10081), .Q(n10080) );
  nnd3s1 U10388 ( .DIN1(n8236), .DIN2(n8536), .DIN3(n8506), .Q(n10081) );
  nnd3s1 U10389 ( .DIN1(n10082), .DIN2(n1444), .DIN3(sa00[0]), .Q(n8506) );
  nnd3s1 U10390 ( .DIN1(sa00[0]), .DIN2(n1430), .DIN3(n10083), .Q(n8236) );
  hi1s1 U10391 ( .DIN(n8967), .Q(n8197) );
  nnd2s1 U10392 ( .DIN1(n8198), .DIN2(n10084), .Q(n10079) );
  nnd2s1 U10393 ( .DIN1(n8535), .DIN2(n8996), .Q(n10084) );
  nnd3s1 U10394 ( .DIN1(n1363), .DIN2(n1430), .DIN3(n10083), .Q(n8535) );
  hi1s1 U10395 ( .DIN(n7988), .Q(n8198) );
  nnd2s1 U10396 ( .DIN1(n8221), .DIN2(n10085), .Q(n10078) );
  nnd2s1 U10397 ( .DIN1(n8500), .DIN2(n8505), .Q(n10085) );
  nnd2s1 U10398 ( .DIN1(n10076), .DIN2(n10062), .Q(n8500) );
  hi1s1 U10399 ( .DIN(n8958), .Q(n8221) );
  nnd3s1 U10400 ( .DIN1(sa00[0]), .DIN2(n1430), .DIN3(n10055), .Q(n8958) );
  nor2s1 U10401 ( .DIN1(n8215), .DIN2(n8540), .Q(n10068) );
  nnd2s1 U10402 ( .DIN1(n10061), .DIN2(n10086), .Q(n8215) );
  and2s1 U10403 ( .DIN1(n8519), .DIN2(n10087), .Q(n10067) );
  nnd4s1 U10404 ( .DIN1(n8004), .DIN2(n8000), .DIN3(n8232), .DIN4(n8003), 
        .Q(n10087) );
  nnd2s1 U10405 ( .DIN1(n10077), .DIN2(n10088), .Q(n8232) );
  nnd2s1 U10406 ( .DIN1(n10088), .DIN2(n10062), .Q(n8000) );
  nor2s1 U10407 ( .DIN1(n1519), .DIN2(n1401), .Q(n10062) );
  nnd2s1 U10408 ( .DIN1(n10086), .DIN2(n10075), .Q(n8004) );
  hi1s1 U10409 ( .DIN(n8212), .Q(n8519) );
  nnd3s1 U10410 ( .DIN1(sa00[1]), .DIN2(n1363), .DIN3(n10083), .Q(n8212) );
  nnd3s1 U10411 ( .DIN1(n10089), .DIN2(n10090), .DIN3(n10091), .Q(n10026) );
  nnd2s1 U10412 ( .DIN1(n7997), .DIN2(n8494), .Q(n10091) );
  hi1s1 U10413 ( .DIN(n7990), .Q(n8494) );
  hi1s1 U10414 ( .DIN(n8564), .Q(n7997) );
  nnd3s1 U10415 ( .DIN1(sa00[2]), .DIN2(n1363), .DIN3(n10092), .Q(n8564) );
  nnd2s1 U10416 ( .DIN1(n9031), .DIN2(n8492), .Q(n10090) );
  hi1s1 U10417 ( .DIN(n8540), .Q(n8492) );
  nnd3s1 U10418 ( .DIN1(sa00[1]), .DIN2(sa00[0]), .DIN3(n10083), .Q(n8540) );
  and2s1 U10419 ( .DIN1(sa00[3]), .DIN2(sa00[2]), .Q(n10083) );
  hi1s1 U10420 ( .DIN(n7999), .Q(n9031) );
  nnd2s1 U10421 ( .DIN1(n8186), .DIN2(n7984), .Q(n10089) );
  hi1s1 U10422 ( .DIN(n8194), .Q(n7984) );
  nnd2s1 U10423 ( .DIN1(n10086), .DIN2(n10088), .Q(n8194) );
  hi1s1 U10424 ( .DIN(n8959), .Q(n8186) );
  nnd4s1 U10425 ( .DIN1(n10093), .DIN2(n10094), .DIN3(n10095), .DIN4(n10096), 
        .Q(n10025) );
  nnd2s1 U10426 ( .DIN1(n9026), .DIN2(n10097), .Q(n10096) );
  nnd2s1 U10427 ( .DIN1(n8545), .DIN2(n9025), .Q(n10097) );
  nnd3s1 U10428 ( .DIN1(sa00[2]), .DIN2(sa00[0]), .DIN3(n10092), .Q(n9025) );
  hi1s1 U10429 ( .DIN(n8505), .Q(n9026) );
  nnd2s1 U10430 ( .DIN1(n10066), .DIN2(n10088), .Q(n8505) );
  and2s1 U10431 ( .DIN1(sa00[4]), .DIN2(sa00[6]), .Q(n10088) );
  nnd2s1 U10432 ( .DIN1(n8518), .DIN2(n10098), .Q(n10095) );
  nnd4s1 U10433 ( .DIN1(n8545), .DIN2(n8996), .DIN3(n8536), .DIN4(n8959), 
        .Q(n10098) );
  nnd3s1 U10434 ( .DIN1(sa00[0]), .DIN2(n10082), .DIN3(sa00[2]), .Q(n8959) );
  nnd3s1 U10435 ( .DIN1(n10055), .DIN2(sa00[0]), .DIN3(sa00[1]), .Q(n8536) );
  and2s1 U10436 ( .DIN1(sa00[3]), .DIN2(n1444), .Q(n10055) );
  nnd3s1 U10437 ( .DIN1(sa00[0]), .DIN2(n1444), .DIN3(n10092), .Q(n8996) );
  nnd3s1 U10438 ( .DIN1(n1363), .DIN2(n1444), .DIN3(n10082), .Q(n8545) );
  hi1s1 U10439 ( .DIN(n8003), .Q(n8518) );
  nnd2s1 U10440 ( .DIN1(n10066), .DIN2(n10076), .Q(n8003) );
  nnd2s1 U10441 ( .DIN1(n8233), .DIN2(n9000), .Q(n10094) );
  nnd2s1 U10442 ( .DIN1(n8967), .DIN2(n7990), .Q(n9000) );
  nnd2s1 U10443 ( .DIN1(n10077), .DIN2(n10075), .Q(n7990) );
  nnd2s1 U10444 ( .DIN1(n10066), .DIN2(n10075), .Q(n8967) );
  and2s1 U10445 ( .DIN1(sa00[6]), .DIN2(n1531), .Q(n10075) );
  nor2s1 U10446 ( .DIN1(sa00[7]), .DIN2(sa00[5]), .Q(n10066) );
  hi1s1 U10447 ( .DIN(n8539), .Q(n8233) );
  nnd3s1 U10448 ( .DIN1(n10082), .DIN2(n1363), .DIN3(sa00[2]), .Q(n8539) );
  nor2s1 U10449 ( .DIN1(sa00[3]), .DIN2(sa00[1]), .Q(n10082) );
  nnd2s1 U10450 ( .DIN1(n7982), .DIN2(n8528), .Q(n10093) );
  nnd2s1 U10451 ( .DIN1(n7988), .DIN2(n7999), .Q(n8528) );
  nnd2s1 U10452 ( .DIN1(n10076), .DIN2(n10086), .Q(n7999) );
  nor2s1 U10453 ( .DIN1(n1519), .DIN2(sa00[5]), .Q(n10086) );
  nor2s1 U10454 ( .DIN1(sa00[6]), .DIN2(sa00[4]), .Q(n10076) );
  nnd2s1 U10455 ( .DIN1(n10061), .DIN2(n10077), .Q(n7988) );
  nor2s1 U10456 ( .DIN1(n1401), .DIN2(sa00[7]), .Q(n10077) );
  nor2s1 U10457 ( .DIN1(n1531), .DIN2(sa00[6]), .Q(n10061) );
  hi1s1 U10458 ( .DIN(n8538), .Q(n7982) );
  nnd3s1 U10459 ( .DIN1(n1363), .DIN2(n1444), .DIN3(n10092), .Q(n8538) );
  nor2s1 U10460 ( .DIN1(n1430), .DIN2(sa00[3]), .Q(n10092) );
  xor2s1 U10461 ( .DIN1(n1473), .DIN2(n5053), .Q(n9631) );
  hi1s1 U10462 ( .DIN(n7712), .Q(n5053) );
  or4s1 U10463 ( .DIN1(n10099), .DIN2(n10100), .DIN3(n10101), .DIN4(n10102), 
        .Q(n7712) );
  nnd4s1 U10464 ( .DIN1(n8714), .DIN2(n10103), .DIN3(n10104), .DIN4(n10105), 
        .Q(n10102) );
  nnd2s1 U10465 ( .DIN1(n8339), .DIN2(n9242), .Q(n10105) );
  nnd2s1 U10466 ( .DIN1(n8768), .DIN2(n7919), .Q(n9242) );
  nnd2s1 U10467 ( .DIN1(n8380), .DIN2(n7921), .Q(n10104) );
  nnd2s1 U10468 ( .DIN1(n8359), .DIN2(n8737), .Q(n7921) );
  nnd2s1 U10469 ( .DIN1(n9191), .DIN2(n8350), .Q(n10103) );
  nnd2s1 U10470 ( .DIN1(n8373), .DIN2(n7901), .Q(n8714) );
  nnd4s1 U10471 ( .DIN1(n10106), .DIN2(n10107), .DIN3(n10108), .DIN4(n10109), 
        .Q(n10101) );
  nnd2s1 U10472 ( .DIN1(n7892), .DIN2(n10110), .Q(n10109) );
  nnd2s1 U10473 ( .DIN1(n8105), .DIN2(n8347), .Q(n10110) );
  nnd2s1 U10474 ( .DIN1(n8338), .DIN2(n10111), .Q(n10108) );
  nnd2s1 U10475 ( .DIN1(n8772), .DIN2(n8764), .Q(n10111) );
  or2s1 U10476 ( .DIN1(n8379), .DIN2(n8361), .Q(n10107) );
  nor2s1 U10477 ( .DIN1(n7912), .DIN2(n8350), .Q(n8361) );
  nnd2s1 U10478 ( .DIN1(n8748), .DIN2(n8371), .Q(n10106) );
  nnd2s1 U10479 ( .DIN1(n8356), .DIN2(n8104), .Q(n8371) );
  nnd3s1 U10480 ( .DIN1(n9365), .DIN2(n9373), .DIN3(n7883), .Q(n10100) );
  nor4s1 U10481 ( .DIN1(n10112), .DIN2(n10113), .DIN3(n10114), .DIN4(n10115), 
        .Q(n7883) );
  nnd4s1 U10482 ( .DIN1(n10116), .DIN2(n10117), .DIN3(n10118), .DIN4(n10119), 
        .Q(n10115) );
  nnd2s1 U10483 ( .DIN1(n7916), .DIN2(n7900), .Q(n10119) );
  nor2s1 U10484 ( .DIN1(n10120), .DIN2(n9161), .Q(n10118) );
  nor2s1 U10485 ( .DIN1(n8359), .DIN2(n7918), .Q(n9161) );
  nor2s1 U10486 ( .DIN1(n8347), .DIN2(n8383), .Q(n10120) );
  nnd2s1 U10487 ( .DIN1(n8370), .DIN2(n7899), .Q(n10117) );
  nnd2s1 U10488 ( .DIN1(n8339), .DIN2(n8357), .Q(n10116) );
  hi1s1 U10489 ( .DIN(n7914), .Q(n8339) );
  nnd3s1 U10490 ( .DIN1(n10121), .DIN2(n10122), .DIN3(n10123), .Q(n10114) );
  nnd2s1 U10491 ( .DIN1(n8350), .DIN2(n8755), .Q(n10123) );
  nnd2s1 U10492 ( .DIN1(n8356), .DIN2(n8347), .Q(n8755) );
  nnd2s1 U10493 ( .DIN1(n7901), .DIN2(n10124), .Q(n10122) );
  nnd3s1 U10494 ( .DIN1(n8765), .DIN2(n9126), .DIN3(n8772), .Q(n10124) );
  nnd2s1 U10495 ( .DIN1(n8349), .DIN2(n10125), .Q(n10121) );
  nnd3s1 U10496 ( .DIN1(n8767), .DIN2(n9125), .DIN3(n8735), .Q(n10125) );
  nor2s1 U10497 ( .DIN1(n8735), .DIN2(n8364), .Q(n10113) );
  nor2s1 U10498 ( .DIN1(n9232), .DIN2(n8734), .Q(n10112) );
  nor2s1 U10499 ( .DIN1(n8102), .DIN2(n7920), .Q(n9232) );
  and4s1 U10500 ( .DIN1(n10126), .DIN2(n10127), .DIN3(n10128), .DIN4(n10129), 
        .Q(n9373) );
  and4s1 U10501 ( .DIN1(n10130), .DIN2(n9175), .DIN3(n10131), .DIN4(n10132), 
        .Q(n10129) );
  nnd2s1 U10502 ( .DIN1(n8373), .DIN2(n9191), .Q(n10132) );
  nnd2s1 U10503 ( .DIN1(n7900), .DIN2(n8091), .Q(n10131) );
  nnd2s1 U10504 ( .DIN1(n7912), .DIN2(n9196), .Q(n9175) );
  nnd2s1 U10505 ( .DIN1(n7892), .DIN2(n7916), .Q(n10130) );
  and3s1 U10506 ( .DIN1(n10133), .DIN2(n10134), .DIN3(n10135), .Q(n10128) );
  nnd2s1 U10507 ( .DIN1(n8370), .DIN2(n10136), .Q(n10135) );
  nnd2s1 U10508 ( .DIN1(n8109), .DIN2(n8356), .Q(n10136) );
  nnd2s1 U10509 ( .DIN1(n7891), .DIN2(n10137), .Q(n10134) );
  nnd2s1 U10510 ( .DIN1(n7914), .DIN2(n8109), .Q(n10137) );
  nnd2s1 U10511 ( .DIN1(n8340), .DIN2(n9224), .Q(n10133) );
  nnd2s1 U10512 ( .DIN1(n8359), .DIN2(n8379), .Q(n9224) );
  nnd2s1 U10513 ( .DIN1(n8106), .DIN2(n10138), .Q(n10127) );
  nnd3s1 U10514 ( .DIN1(n8379), .DIN2(n8108), .DIN3(n7915), .Q(n10138) );
  hi1s1 U10515 ( .DIN(n7918), .Q(n8106) );
  or2s1 U10516 ( .DIN1(n8356), .DIN2(n9615), .Q(n10126) );
  nor2s1 U10517 ( .DIN1(n7902), .DIN2(n7920), .Q(n9615) );
  nor4s1 U10518 ( .DIN1(n10139), .DIN2(n10140), .DIN3(n10141), .DIN4(n10142), 
        .Q(n9365) );
  nnd4s1 U10519 ( .DIN1(n10143), .DIN2(n10144), .DIN3(n10145), .DIN4(n10146), 
        .Q(n10142) );
  nor2s1 U10520 ( .DIN1(n10147), .DIN2(n10148), .Q(n10146) );
  nor2s1 U10521 ( .DIN1(n8765), .DIN2(n8104), .Q(n10148) );
  nor2s1 U10522 ( .DIN1(n8767), .DIN2(n8109), .Q(n10147) );
  nnd2s1 U10523 ( .DIN1(n8357), .DIN2(n8724), .Q(n10145) );
  or2s1 U10524 ( .DIN1(n9162), .DIN2(n8729), .Q(n10144) );
  nor2s1 U10525 ( .DIN1(n7916), .DIN2(n8724), .Q(n8729) );
  nnd2s1 U10526 ( .DIN1(n7890), .DIN2(n7898), .Q(n10143) );
  nnd3s1 U10527 ( .DIN1(n10149), .DIN2(n10150), .DIN3(n10151), .Q(n10141) );
  nnd2s1 U10528 ( .DIN1(n7891), .DIN2(n8788), .Q(n10151) );
  nnd2s1 U10529 ( .DIN1(n8104), .DIN2(n8737), .Q(n8788) );
  hi1s1 U10530 ( .DIN(n8383), .Q(n7891) );
  nnd2s1 U10531 ( .DIN1(n8091), .DIN2(n10152), .Q(n10150) );
  nnd2s1 U10532 ( .DIN1(n9125), .DIN2(n8362), .Q(n10152) );
  nnd2s1 U10533 ( .DIN1(n8349), .DIN2(n10153), .Q(n10149) );
  nnd2s1 U10534 ( .DIN1(n7911), .DIN2(n9162), .Q(n10153) );
  nor2s1 U10535 ( .DIN1(n10154), .DIN2(n7915), .Q(n10140) );
  nor2s1 U10536 ( .DIN1(n7892), .DIN2(n8340), .Q(n10154) );
  nor2s1 U10537 ( .DIN1(n10155), .DIN2(n8095), .Q(n10139) );
  nor2s1 U10538 ( .DIN1(n7898), .DIN2(n8102), .Q(n10155) );
  nnd4s1 U10539 ( .DIN1(n9572), .DIN2(n10156), .DIN3(n10157), .DIN4(n10158), 
        .Q(n10099) );
  nnd2s1 U10540 ( .DIN1(n7890), .DIN2(n8357), .Q(n10158) );
  nnd2s1 U10541 ( .DIN1(n8340), .DIN2(n7916), .Q(n10157) );
  nnd2s1 U10542 ( .DIN1(n8747), .DIN2(n8370), .Q(n10156) );
  nor3s1 U10543 ( .DIN1(n10159), .DIN2(n10160), .DIN3(n10161), .Q(n9572) );
  nnd4s1 U10544 ( .DIN1(n7886), .DIN2(n9374), .DIN3(n9369), .DIN4(n10162), 
        .Q(n10161) );
  and3s1 U10545 ( .DIN1(n10163), .DIN2(n10164), .DIN3(n10165), .Q(n10162) );
  nnd2s1 U10546 ( .DIN1(n8338), .DIN2(n8370), .Q(n10165) );
  nnd2s1 U10547 ( .DIN1(n7893), .DIN2(n8357), .Q(n10164) );
  hi1s1 U10548 ( .DIN(n8764), .Q(n8357) );
  hi1s1 U10549 ( .DIN(n8109), .Q(n7893) );
  nnd2s1 U10550 ( .DIN1(n8748), .DIN2(n7908), .Q(n10163) );
  hi1s1 U10551 ( .DIN(n8364), .Q(n7908) );
  and4s1 U10552 ( .DIN1(n10166), .DIN2(n10167), .DIN3(n10168), .DIN4(n10169), 
        .Q(n9369) );
  and4s1 U10553 ( .DIN1(n10170), .DIN2(n10171), .DIN3(n9140), .DIN4(n8722), 
        .Q(n10169) );
  nnd2s1 U10554 ( .DIN1(n7902), .DIN2(n8091), .Q(n8722) );
  nnd2s1 U10555 ( .DIN1(n8340), .DIN2(n7890), .Q(n9140) );
  nnd2s1 U10556 ( .DIN1(n8102), .DIN2(n7916), .Q(n10171) );
  nnd2s1 U10557 ( .DIN1(n8338), .DIN2(n8748), .Q(n10170) );
  and3s1 U10558 ( .DIN1(n10172), .DIN2(n10173), .DIN3(n10174), .Q(n10168) );
  nnd2s1 U10559 ( .DIN1(n7903), .DIN2(n9584), .Q(n10174) );
  nnd2s1 U10560 ( .DIN1(n8733), .DIN2(n8383), .Q(n9584) );
  nnd2s1 U10561 ( .DIN1(n7900), .DIN2(n10175), .Q(n10173) );
  nnd2s1 U10562 ( .DIN1(n9169), .DIN2(n8364), .Q(n10175) );
  nor2s1 U10563 ( .DIN1(n8747), .DIN2(n8724), .Q(n9169) );
  hi1s1 U10564 ( .DIN(n8359), .Q(n8724) );
  nnd2s1 U10565 ( .DIN1(n9196), .DIN2(n10176), .Q(n10172) );
  nnd2s1 U10566 ( .DIN1(n8768), .DIN2(n7918), .Q(n10176) );
  nnd2s1 U10567 ( .DIN1(n8747), .DIN2(n10177), .Q(n10167) );
  nnd2s1 U10568 ( .DIN1(n8790), .DIN2(n7911), .Q(n10177) );
  nnd2s1 U10569 ( .DIN1(n8350), .DIN2(n10178), .Q(n10166) );
  nnd3s1 U10570 ( .DIN1(n8105), .DIN2(n7915), .DIN3(n8109), .Q(n10178) );
  and4s1 U10571 ( .DIN1(n10179), .DIN2(n10180), .DIN3(n10181), .DIN4(n10182), 
        .Q(n9374) );
  nor4s1 U10572 ( .DIN1(n10183), .DIN2(n10184), .DIN3(n10185), .DIN4(n10186), 
        .Q(n10182) );
  nor2s1 U10573 ( .DIN1(n10187), .DIN2(n8104), .Q(n10186) );
  nor2s1 U10574 ( .DIN1(n8340), .DIN2(n8370), .Q(n10187) );
  nor2s1 U10575 ( .DIN1(n10188), .DIN2(n8737), .Q(n10185) );
  nor2s1 U10576 ( .DIN1(n7898), .DIN2(n7902), .Q(n10188) );
  hi1s1 U10577 ( .DIN(n7911), .Q(n7902) );
  nnd3s1 U10578 ( .DIN1(n10189), .DIN2(n1364), .DIN3(sa22[1]), .Q(n7911) );
  nor2s1 U10579 ( .DIN1(n10190), .DIN2(n8383), .Q(n10184) );
  nor2s1 U10580 ( .DIN1(n8090), .DIN2(n8747), .Q(n10190) );
  nnd3s1 U10581 ( .DIN1(n10191), .DIN2(n10192), .DIN3(n10193), .Q(n10183) );
  nnd2s1 U10582 ( .DIN1(n7898), .DIN2(n9191), .Q(n10193) );
  nnd2s1 U10583 ( .DIN1(n7899), .DIN2(n10194), .Q(n10192) );
  nnd2s1 U10584 ( .DIN1(n8362), .DIN2(n8735), .Q(n10194) );
  nnd2s1 U10585 ( .DIN1(n7912), .DIN2(n9399), .Q(n10191) );
  nnd2s1 U10586 ( .DIN1(n8356), .DIN2(n8359), .Q(n9399) );
  nnd2s1 U10587 ( .DIN1(n10195), .DIN2(n10196), .Q(n8359) );
  hi1s1 U10588 ( .DIN(n8772), .Q(n7912) );
  and3s1 U10589 ( .DIN1(n10197), .DIN2(n10198), .DIN3(n10199), .Q(n10181) );
  nnd2s1 U10590 ( .DIN1(n8380), .DIN2(n8349), .Q(n10199) );
  hi1s1 U10591 ( .DIN(n8105), .Q(n8349) );
  nnd2s1 U10592 ( .DIN1(n8090), .DIN2(n8373), .Q(n10198) );
  nnd2s1 U10593 ( .DIN1(n7903), .DIN2(n7920), .Q(n10197) );
  nnd2s1 U10594 ( .DIN1(n8102), .DIN2(n7890), .Q(n10180) );
  nnd2s1 U10595 ( .DIN1(n7916), .DIN2(n8350), .Q(n10179) );
  hi1s1 U10596 ( .DIN(n8765), .Q(n8350) );
  hi1s1 U10597 ( .DIN(n9186), .Q(n7916) );
  nnd2s1 U10598 ( .DIN1(n10195), .DIN2(n10200), .Q(n9186) );
  nor4s1 U10599 ( .DIN1(n10201), .DIN2(n10202), .DIN3(n10203), .DIN4(n10204), 
        .Q(n7886) );
  nnd4s1 U10600 ( .DIN1(n10205), .DIN2(n10206), .DIN3(n10207), .DIN4(n10208), 
        .Q(n10204) );
  nnd2s1 U10601 ( .DIN1(n8373), .DIN2(n7899), .Q(n10208) );
  hi1s1 U10602 ( .DIN(n9162), .Q(n8373) );
  nnd2s1 U10603 ( .DIN1(n7892), .DIN2(n7901), .Q(n10207) );
  hi1s1 U10604 ( .DIN(n8737), .Q(n7901) );
  nnd2s1 U10605 ( .DIN1(n10209), .DIN2(n10196), .Q(n8737) );
  hi1s1 U10606 ( .DIN(n8733), .Q(n7892) );
  nnd3s1 U10607 ( .DIN1(n1364), .DIN2(n1431), .DIN3(n10189), .Q(n8733) );
  nnd2s1 U10608 ( .DIN1(n8090), .DIN2(n7920), .Q(n10206) );
  hi1s1 U10609 ( .DIN(n8735), .Q(n7920) );
  hi1s1 U10610 ( .DIN(n8379), .Q(n8090) );
  nnd2s1 U10611 ( .DIN1(n7890), .DIN2(n7900), .Q(n10205) );
  hi1s1 U10612 ( .DIN(n8356), .Q(n7890) );
  nnd2s1 U10613 ( .DIN1(n10210), .DIN2(n10211), .Q(n8356) );
  nnd3s1 U10614 ( .DIN1(n10212), .DIN2(n10213), .DIN3(n10214), .Q(n10203) );
  nnd2s1 U10615 ( .DIN1(n8338), .DIN2(n10215), .Q(n10214) );
  nnd3s1 U10616 ( .DIN1(n8383), .DIN2(n8765), .DIN3(n8735), .Q(n10215) );
  nnd3s1 U10617 ( .DIN1(n10216), .DIN2(n1445), .DIN3(sa22[0]), .Q(n8735) );
  nnd3s1 U10618 ( .DIN1(sa22[0]), .DIN2(n1431), .DIN3(n10217), .Q(n8383) );
  hi1s1 U10619 ( .DIN(n9133), .Q(n8338) );
  nnd2s1 U10620 ( .DIN1(n7903), .DIN2(n10218), .Q(n10213) );
  nnd2s1 U10621 ( .DIN1(n8764), .DIN2(n9162), .Q(n10218) );
  nnd3s1 U10622 ( .DIN1(n1364), .DIN2(n1431), .DIN3(n10217), .Q(n8764) );
  hi1s1 U10623 ( .DIN(n8095), .Q(n7903) );
  nnd2s1 U10624 ( .DIN1(n8370), .DIN2(n10219), .Q(n10212) );
  nnd2s1 U10625 ( .DIN1(n7914), .DIN2(n8734), .Q(n10219) );
  nnd2s1 U10626 ( .DIN1(n10210), .DIN2(n10196), .Q(n7914) );
  hi1s1 U10627 ( .DIN(n9125), .Q(n8370) );
  nnd3s1 U10628 ( .DIN1(sa22[0]), .DIN2(n1431), .DIN3(n10189), .Q(n9125) );
  nor2s1 U10629 ( .DIN1(n8364), .DIN2(n7919), .Q(n10202) );
  nnd2s1 U10630 ( .DIN1(n10195), .DIN2(n10220), .Q(n8364) );
  and2s1 U10631 ( .DIN1(n8748), .DIN2(n10221), .Q(n10201) );
  nnd4s1 U10632 ( .DIN1(n8109), .DIN2(n8105), .DIN3(n8379), .DIN4(n8108), 
        .Q(n10221) );
  nnd2s1 U10633 ( .DIN1(n10211), .DIN2(n10222), .Q(n8379) );
  nnd2s1 U10634 ( .DIN1(n10222), .DIN2(n10196), .Q(n8105) );
  nor2s1 U10635 ( .DIN1(n1520), .DIN2(n1402), .Q(n10196) );
  nnd2s1 U10636 ( .DIN1(n10220), .DIN2(n10209), .Q(n8109) );
  hi1s1 U10637 ( .DIN(n8362), .Q(n8748) );
  nnd3s1 U10638 ( .DIN1(sa22[1]), .DIN2(n1364), .DIN3(n10217), .Q(n8362) );
  nnd3s1 U10639 ( .DIN1(n10223), .DIN2(n10224), .DIN3(n10225), .Q(n10160) );
  nnd2s1 U10640 ( .DIN1(n8102), .DIN2(n7899), .Q(n10225) );
  hi1s1 U10641 ( .DIN(n7915), .Q(n7899) );
  hi1s1 U10642 ( .DIN(n8790), .Q(n8102) );
  nnd3s1 U10643 ( .DIN1(sa22[2]), .DIN2(n1364), .DIN3(n10226), .Q(n8790) );
  nnd2s1 U10644 ( .DIN1(n9196), .DIN2(n7898), .Q(n10224) );
  hi1s1 U10645 ( .DIN(n7919), .Q(n7898) );
  nnd3s1 U10646 ( .DIN1(sa22[1]), .DIN2(sa22[0]), .DIN3(n10217), .Q(n7919) );
  and2s1 U10647 ( .DIN1(sa22[3]), .DIN2(sa22[2]), .Q(n10217) );
  hi1s1 U10648 ( .DIN(n8104), .Q(n9196) );
  nnd2s1 U10649 ( .DIN1(n8340), .DIN2(n8091), .Q(n10223) );
  hi1s1 U10650 ( .DIN(n8347), .Q(n8091) );
  nnd2s1 U10651 ( .DIN1(n10220), .DIN2(n10222), .Q(n8347) );
  hi1s1 U10652 ( .DIN(n9126), .Q(n8340) );
  nnd4s1 U10653 ( .DIN1(n10227), .DIN2(n10228), .DIN3(n10229), .DIN4(n10230), 
        .Q(n10159) );
  nnd2s1 U10654 ( .DIN1(n9191), .DIN2(n10231), .Q(n10230) );
  nnd2s1 U10655 ( .DIN1(n8772), .DIN2(n7918), .Q(n10231) );
  nnd3s1 U10656 ( .DIN1(sa22[2]), .DIN2(sa22[0]), .DIN3(n10226), .Q(n7918) );
  hi1s1 U10657 ( .DIN(n8734), .Q(n9191) );
  nnd2s1 U10658 ( .DIN1(n10200), .DIN2(n10222), .Q(n8734) );
  and2s1 U10659 ( .DIN1(sa22[4]), .DIN2(sa22[6]), .Q(n10222) );
  nnd2s1 U10660 ( .DIN1(n8747), .DIN2(n10232), .Q(n10229) );
  nnd4s1 U10661 ( .DIN1(n8772), .DIN2(n9162), .DIN3(n8765), .DIN4(n9126), 
        .Q(n10232) );
  nnd3s1 U10662 ( .DIN1(sa22[0]), .DIN2(n10216), .DIN3(sa22[2]), .Q(n9126) );
  nnd3s1 U10663 ( .DIN1(n10189), .DIN2(sa22[0]), .DIN3(sa22[1]), .Q(n8765) );
  and2s1 U10664 ( .DIN1(sa22[3]), .DIN2(n1445), .Q(n10189) );
  nnd3s1 U10665 ( .DIN1(sa22[0]), .DIN2(n1445), .DIN3(n10226), .Q(n9162) );
  nnd3s1 U10666 ( .DIN1(n1364), .DIN2(n1445), .DIN3(n10216), .Q(n8772) );
  hi1s1 U10667 ( .DIN(n8108), .Q(n8747) );
  nnd2s1 U10668 ( .DIN1(n10200), .DIN2(n10210), .Q(n8108) );
  nnd2s1 U10669 ( .DIN1(n8380), .DIN2(n9166), .Q(n10228) );
  nnd2s1 U10670 ( .DIN1(n9133), .DIN2(n7915), .Q(n9166) );
  nnd2s1 U10671 ( .DIN1(n10211), .DIN2(n10209), .Q(n7915) );
  nnd2s1 U10672 ( .DIN1(n10200), .DIN2(n10209), .Q(n9133) );
  and2s1 U10673 ( .DIN1(sa22[6]), .DIN2(n1532), .Q(n10209) );
  nor2s1 U10674 ( .DIN1(sa22[7]), .DIN2(sa22[5]), .Q(n10200) );
  hi1s1 U10675 ( .DIN(n8768), .Q(n8380) );
  nnd3s1 U10676 ( .DIN1(n10216), .DIN2(n1364), .DIN3(sa22[2]), .Q(n8768) );
  nor2s1 U10677 ( .DIN1(sa22[3]), .DIN2(sa22[1]), .Q(n10216) );
  nnd2s1 U10678 ( .DIN1(n7900), .DIN2(n8757), .Q(n10227) );
  nnd2s1 U10679 ( .DIN1(n8095), .DIN2(n8104), .Q(n8757) );
  nnd2s1 U10680 ( .DIN1(n10210), .DIN2(n10220), .Q(n8104) );
  nor2s1 U10681 ( .DIN1(n1520), .DIN2(sa22[5]), .Q(n10220) );
  nor2s1 U10682 ( .DIN1(sa22[6]), .DIN2(sa22[4]), .Q(n10210) );
  nnd2s1 U10683 ( .DIN1(n10195), .DIN2(n10211), .Q(n8095) );
  nor2s1 U10684 ( .DIN1(n1402), .DIN2(sa22[7]), .Q(n10211) );
  nor2s1 U10685 ( .DIN1(n1532), .DIN2(sa22[6]), .Q(n10195) );
  hi1s1 U10686 ( .DIN(n8767), .Q(n7900) );
  nnd3s1 U10687 ( .DIN1(n1364), .DIN2(n1445), .DIN3(n10226), .Q(n8767) );
  nor2s1 U10688 ( .DIN1(n1431), .DIN2(sa22[3]), .Q(n10226) );
  nnd2s1 U10689 ( .DIN1(n10233), .DIN2(n1603), .Q(n9628) );
  xor2s1 U10690 ( .DIN1(w0[0]), .DIN2(text_in_r[96]), .Q(n10233) );
  nnd2s1 U10691 ( .DIN1(n10234), .DIN2(n10235), .Q(N217) );
  nnd2s1 U10692 ( .DIN1(n10236), .DIN2(n1624), .Q(n10235) );
  xor2s1 U10693 ( .DIN1(n10237), .DIN2(n10238), .Q(n10236) );
  xor2s1 U10694 ( .DIN1(n10239), .DIN2(n10240), .Q(n10238) );
  xor2s1 U10695 ( .DIN1(w1[31]), .DIN2(n10241), .Q(n10237) );
  nnd2s1 U10696 ( .DIN1(n10242), .DIN2(n1603), .Q(n10234) );
  xor2s1 U10697 ( .DIN1(w1[31]), .DIN2(text_in_r[95]), .Q(n10242) );
  nnd2s1 U10698 ( .DIN1(n10243), .DIN2(n10244), .Q(N216) );
  nnd2s1 U10699 ( .DIN1(n10245), .DIN2(n1624), .Q(n10244) );
  xor2s1 U10700 ( .DIN1(n10246), .DIN2(n10247), .Q(n10245) );
  xor2s1 U10701 ( .DIN1(n10248), .DIN2(n10249), .Q(n10247) );
  xor2s1 U10702 ( .DIN1(n5075), .DIN2(w1[30]), .Q(n10246) );
  nnd2s1 U10703 ( .DIN1(n10250), .DIN2(n1603), .Q(n10243) );
  xor2s1 U10704 ( .DIN1(w1[30]), .DIN2(text_in_r[94]), .Q(n10250) );
  nnd2s1 U10705 ( .DIN1(n10251), .DIN2(n10252), .Q(N215) );
  nnd2s1 U10706 ( .DIN1(n10253), .DIN2(n1625), .Q(n10252) );
  xor2s1 U10707 ( .DIN1(n10254), .DIN2(n10255), .Q(n10253) );
  xor2s1 U10708 ( .DIN1(n10256), .DIN2(n10257), .Q(n10255) );
  xor2s1 U10709 ( .DIN1(n1485), .DIN2(n5074), .Q(n10254) );
  nnd2s1 U10710 ( .DIN1(n10258), .DIN2(n1603), .Q(n10251) );
  xor2s1 U10711 ( .DIN1(w1[29]), .DIN2(text_in_r[93]), .Q(n10258) );
  nnd3s1 U10712 ( .DIN1(n10259), .DIN2(n10260), .DIN3(n10261), .Q(N214) );
  nnd2s1 U10713 ( .DIN1(n1599), .DIN2(n10262), .Q(n10261) );
  xor2s1 U10714 ( .DIN1(w1[28]), .DIN2(text_in_r[92]), .Q(n10262) );
  nnd2s1 U10715 ( .DIN1(n10263), .DIN2(n10264), .Q(n10260) );
  nnd2s1 U10716 ( .DIN1(n10265), .DIN2(n10266), .Q(n10263) );
  nnd2s1 U10717 ( .DIN1(n10267), .DIN2(n10268), .Q(n10266) );
  nnd2s1 U10718 ( .DIN1(n10269), .DIN2(n10270), .Q(n10265) );
  nnd2s1 U10719 ( .DIN1(n10271), .DIN2(n10272), .Q(n10259) );
  nnd2s1 U10720 ( .DIN1(n10273), .DIN2(n10274), .Q(n10272) );
  nnd2s1 U10721 ( .DIN1(n10269), .DIN2(n10268), .Q(n10274) );
  nnd2s1 U10722 ( .DIN1(n10270), .DIN2(n10267), .Q(n10273) );
  hi1s1 U10723 ( .DIN(n10268), .Q(n10270) );
  xor2s1 U10724 ( .DIN1(n10275), .DIN2(n10276), .Q(n10268) );
  xor2s1 U10725 ( .DIN1(n1541), .DIN2(n5073), .Q(n10275) );
  nnd3s1 U10726 ( .DIN1(n10277), .DIN2(n10278), .DIN3(n10279), .Q(N213) );
  nnd2s1 U10727 ( .DIN1(n1598), .DIN2(n10280), .Q(n10279) );
  xor2s1 U10728 ( .DIN1(w1[27]), .DIN2(text_in_r[91]), .Q(n10280) );
  nnd2s1 U10729 ( .DIN1(n10281), .DIN2(n10282), .Q(n10278) );
  nnd2s1 U10730 ( .DIN1(n10283), .DIN2(n10284), .Q(n10281) );
  nnd2s1 U10731 ( .DIN1(n10285), .DIN2(n10286), .Q(n10284) );
  nnd2s1 U10732 ( .DIN1(n10287), .DIN2(n10288), .Q(n10283) );
  nnd2s1 U10733 ( .DIN1(n10289), .DIN2(n10290), .Q(n10277) );
  nnd2s1 U10734 ( .DIN1(n10291), .DIN2(n10292), .Q(n10290) );
  nnd2s1 U10735 ( .DIN1(n10287), .DIN2(n10286), .Q(n10292) );
  nnd2s1 U10736 ( .DIN1(n10288), .DIN2(n10285), .Q(n10291) );
  hi1s1 U10737 ( .DIN(n10286), .Q(n10288) );
  xor2s1 U10738 ( .DIN1(n10293), .DIN2(n10276), .Q(n10286) );
  xor2s1 U10739 ( .DIN1(n5072), .DIN2(w1[27]), .Q(n10293) );
  nnd2s1 U10740 ( .DIN1(n10294), .DIN2(n10295), .Q(N212) );
  nnd2s1 U10741 ( .DIN1(n10296), .DIN2(n1625), .Q(n10295) );
  xor2s1 U10742 ( .DIN1(n10297), .DIN2(n10298), .Q(n10296) );
  xor2s1 U10743 ( .DIN1(n10299), .DIN2(n10300), .Q(n10298) );
  xor2s1 U10744 ( .DIN1(w1[26]), .DIN2(n10301), .Q(n10297) );
  nnd2s1 U10745 ( .DIN1(n10302), .DIN2(n1602), .Q(n10294) );
  xor2s1 U10746 ( .DIN1(w1[26]), .DIN2(text_in_r[90]), .Q(n10302) );
  nnd2s1 U10747 ( .DIN1(n10303), .DIN2(n10304), .Q(N211) );
  nnd2s1 U10748 ( .DIN1(n10305), .DIN2(n1625), .Q(n10304) );
  xor2s1 U10749 ( .DIN1(n10306), .DIN2(n10307), .Q(n10305) );
  xnr2s1 U10750 ( .DIN1(n10308), .DIN2(n10309), .Q(n10307) );
  xor2s1 U10751 ( .DIN1(n10310), .DIN2(n10276), .Q(n10306) );
  xor2s1 U10752 ( .DIN1(n5070), .DIN2(w1[25]), .Q(n10310) );
  nnd2s1 U10753 ( .DIN1(n10311), .DIN2(n1602), .Q(n10303) );
  xor2s1 U10754 ( .DIN1(w1[25]), .DIN2(text_in_r[89]), .Q(n10311) );
  nnd2s1 U10755 ( .DIN1(n10312), .DIN2(n10313), .Q(N210) );
  nnd2s1 U10756 ( .DIN1(n10314), .DIN2(n1626), .Q(n10313) );
  xor2s1 U10757 ( .DIN1(n10315), .DIN2(n10316), .Q(n10314) );
  xor2s1 U10758 ( .DIN1(n10276), .DIN2(n10317), .Q(n10316) );
  xor2s1 U10759 ( .DIN1(n1486), .DIN2(n5069), .Q(n10315) );
  nnd2s1 U10760 ( .DIN1(n10318), .DIN2(n1602), .Q(n10312) );
  xor2s1 U10761 ( .DIN1(w1[24]), .DIN2(text_in_r[88]), .Q(n10318) );
  nnd2s1 U10762 ( .DIN1(n10319), .DIN2(n10320), .Q(N201) );
  nnd2s1 U10763 ( .DIN1(n10321), .DIN2(n1626), .Q(n10320) );
  xor2s1 U10764 ( .DIN1(n10322), .DIN2(n10323), .Q(n10321) );
  xor2s1 U10765 ( .DIN1(n5701), .DIN2(n10324), .Q(n10323) );
  xor2s1 U10766 ( .DIN1(n5075), .DIN2(n10325), .Q(n10322) );
  xor2s1 U10767 ( .DIN1(n1487), .DIN2(n5051), .Q(n10325) );
  nnd2s1 U10768 ( .DIN1(n10326), .DIN2(n1602), .Q(n10319) );
  xor2s1 U10769 ( .DIN1(w1[23]), .DIN2(text_in_r[87]), .Q(n10326) );
  nnd3s1 U10770 ( .DIN1(n10327), .DIN2(n10328), .DIN3(n10329), .Q(N200) );
  nnd2s1 U10771 ( .DIN1(n1599), .DIN2(n10330), .Q(n10329) );
  xor2s1 U10772 ( .DIN1(w1[22]), .DIN2(text_in_r[86]), .Q(n10330) );
  nnd2s1 U10773 ( .DIN1(n10331), .DIN2(n10332), .Q(n10328) );
  nnd2s1 U10774 ( .DIN1(n10333), .DIN2(n10334), .Q(n10331) );
  nnd2s1 U10775 ( .DIN1(n10335), .DIN2(n10336), .Q(n10334) );
  nnd2s1 U10776 ( .DIN1(n10337), .DIN2(n10338), .Q(n10333) );
  nnd2s1 U10777 ( .DIN1(n10248), .DIN2(n10339), .Q(n10327) );
  nnd2s1 U10778 ( .DIN1(n10340), .DIN2(n10341), .Q(n10339) );
  nnd2s1 U10779 ( .DIN1(n10337), .DIN2(n10336), .Q(n10341) );
  nnd2s1 U10780 ( .DIN1(n10338), .DIN2(n10335), .Q(n10340) );
  hi1s1 U10781 ( .DIN(n10336), .Q(n10338) );
  xnr2s1 U10782 ( .DIN1(n5074), .DIN2(n10342), .Q(n10336) );
  xor2s1 U10783 ( .DIN1(w1[22]), .DIN2(n5050), .Q(n10342) );
  nnd3s1 U10784 ( .DIN1(n10343), .DIN2(n10344), .DIN3(n10345), .Q(N199) );
  nnd2s1 U10785 ( .DIN1(n1598), .DIN2(n10346), .Q(n10345) );
  xor2s1 U10786 ( .DIN1(w1[21]), .DIN2(text_in_r[85]), .Q(n10346) );
  nnd2s1 U10787 ( .DIN1(n10347), .DIN2(n10348), .Q(n10344) );
  nnd2s1 U10788 ( .DIN1(n10349), .DIN2(n10350), .Q(n10347) );
  nnd2s1 U10789 ( .DIN1(n10351), .DIN2(n10352), .Q(n10350) );
  nnd2s1 U10790 ( .DIN1(n10353), .DIN2(n10354), .Q(n10349) );
  nnd2s1 U10791 ( .DIN1(n10256), .DIN2(n10355), .Q(n10343) );
  nnd2s1 U10792 ( .DIN1(n10356), .DIN2(n10357), .Q(n10355) );
  nnd2s1 U10793 ( .DIN1(n10353), .DIN2(n10352), .Q(n10357) );
  nnd2s1 U10794 ( .DIN1(n10354), .DIN2(n10351), .Q(n10356) );
  hi1s1 U10795 ( .DIN(n10352), .Q(n10354) );
  xor2s1 U10796 ( .DIN1(n10358), .DIN2(n10359), .Q(n10352) );
  xor2s1 U10797 ( .DIN1(w1[21]), .DIN2(n5049), .Q(n10359) );
  nnd2s1 U10798 ( .DIN1(n10360), .DIN2(n10361), .Q(N198) );
  nnd2s1 U10799 ( .DIN1(n10362), .DIN2(n1627), .Q(n10361) );
  xor2s1 U10800 ( .DIN1(n10363), .DIN2(n10364), .Q(n10362) );
  xor2s1 U10801 ( .DIN1(n10365), .DIN2(n10366), .Q(n10364) );
  xor2s1 U10802 ( .DIN1(n5698), .DIN2(n10264), .Q(n10366) );
  hi1s1 U10803 ( .DIN(n10271), .Q(n10264) );
  xor2s1 U10804 ( .DIN1(n5072), .DIN2(n10367), .Q(n10363) );
  xor2s1 U10805 ( .DIN1(n1488), .DIN2(n5048), .Q(n10367) );
  nnd2s1 U10806 ( .DIN1(n10368), .DIN2(n1602), .Q(n10360) );
  xor2s1 U10807 ( .DIN1(w1[20]), .DIN2(text_in_r[84]), .Q(n10368) );
  nnd2s1 U10808 ( .DIN1(n10369), .DIN2(n10370), .Q(N197) );
  nnd2s1 U10809 ( .DIN1(n10371), .DIN2(n1627), .Q(n10370) );
  xor2s1 U10810 ( .DIN1(n10372), .DIN2(n10373), .Q(n10371) );
  xor2s1 U10811 ( .DIN1(n10365), .DIN2(n10374), .Q(n10373) );
  xor2s1 U10812 ( .DIN1(n5425), .DIN2(n10282), .Q(n10374) );
  xor2s1 U10813 ( .DIN1(n10301), .DIN2(n10375), .Q(n10372) );
  xnr2s1 U10814 ( .DIN1(w1[19]), .DIN2(n5047), .Q(n10375) );
  nnd2s1 U10815 ( .DIN1(n10376), .DIN2(n1602), .Q(n10369) );
  xor2s1 U10816 ( .DIN1(w1[19]), .DIN2(text_in_r[83]), .Q(n10376) );
  nnd2s1 U10817 ( .DIN1(n10377), .DIN2(n10378), .Q(N196) );
  nnd2s1 U10818 ( .DIN1(n10379), .DIN2(n1627), .Q(n10378) );
  xor2s1 U10819 ( .DIN1(n10380), .DIN2(n10381), .Q(n10379) );
  xor2s1 U10820 ( .DIN1(n5424), .DIN2(n10382), .Q(n10381) );
  xor2s1 U10821 ( .DIN1(n5070), .DIN2(n10383), .Q(n10380) );
  xor2s1 U10822 ( .DIN1(n1489), .DIN2(n5046), .Q(n10383) );
  nnd2s1 U10823 ( .DIN1(n10384), .DIN2(n1602), .Q(n10377) );
  xor2s1 U10824 ( .DIN1(w1[18]), .DIN2(text_in_r[82]), .Q(n10384) );
  nnd2s1 U10825 ( .DIN1(n10385), .DIN2(n10386), .Q(N195) );
  nnd2s1 U10826 ( .DIN1(n10387), .DIN2(n1628), .Q(n10386) );
  xor2s1 U10827 ( .DIN1(n10388), .DIN2(n10389), .Q(n10387) );
  xor2s1 U10828 ( .DIN1(n10365), .DIN2(n10390), .Q(n10389) );
  xor2s1 U10829 ( .DIN1(n5423), .DIN2(n10309), .Q(n10390) );
  xnr2s1 U10830 ( .DIN1(n5069), .DIN2(n10391), .Q(n10388) );
  xor2s1 U10831 ( .DIN1(w1[17]), .DIN2(n5045), .Q(n10391) );
  nnd2s1 U10832 ( .DIN1(n10392), .DIN2(n1602), .Q(n10385) );
  xor2s1 U10833 ( .DIN1(w1[17]), .DIN2(text_in_r[81]), .Q(n10392) );
  nnd2s1 U10834 ( .DIN1(n10393), .DIN2(n10394), .Q(N194) );
  nnd2s1 U10835 ( .DIN1(n10395), .DIN2(n1628), .Q(n10394) );
  xor2s1 U10836 ( .DIN1(n10396), .DIN2(n10397), .Q(n10395) );
  xor2s1 U10837 ( .DIN1(n10317), .DIN2(n10365), .Q(n10397) );
  xor2s1 U10838 ( .DIN1(n5076), .DIN2(n5052), .Q(n10365) );
  xor2s1 U10839 ( .DIN1(n1490), .DIN2(n5422), .Q(n10396) );
  nnd2s1 U10840 ( .DIN1(n10398), .DIN2(n1602), .Q(n10393) );
  xor2s1 U10841 ( .DIN1(w1[16]), .DIN2(text_in_r[80]), .Q(n10398) );
  nnd2s1 U10842 ( .DIN1(n10399), .DIN2(n10400), .Q(N185) );
  nnd2s1 U10843 ( .DIN1(n10401), .DIN2(n1628), .Q(n10400) );
  xor2s1 U10844 ( .DIN1(n10402), .DIN2(n10403), .Q(n10401) );
  xor2s1 U10845 ( .DIN1(n10248), .DIN2(n10276), .Q(n10403) );
  hi1s1 U10846 ( .DIN(n10332), .Q(n10248) );
  xor2s1 U10847 ( .DIN1(n5028), .DIN2(n10404), .Q(n10332) );
  hi1s1 U10848 ( .DIN(n5051), .Q(n10404) );
  xor2s1 U10849 ( .DIN1(n1491), .DIN2(n5029), .Q(n10402) );
  nnd2s1 U10850 ( .DIN1(n10405), .DIN2(n1602), .Q(n10399) );
  xor2s1 U10851 ( .DIN1(w1[15]), .DIN2(text_in_r[79]), .Q(n10405) );
  nnd2s1 U10852 ( .DIN1(n10406), .DIN2(n10407), .Q(N184) );
  nnd2s1 U10853 ( .DIN1(n10408), .DIN2(n1629), .Q(n10407) );
  xor2s1 U10854 ( .DIN1(n10409), .DIN2(n10410), .Q(n10408) );
  xnr2s1 U10855 ( .DIN1(w1[14]), .DIN2(n5028), .Q(n10410) );
  xor2s1 U10856 ( .DIN1(n10348), .DIN2(n10240), .Q(n10409) );
  hi1s1 U10857 ( .DIN(n10256), .Q(n10348) );
  xnr2s1 U10858 ( .DIN1(n10411), .DIN2(n5050), .Q(n10256) );
  hi1s1 U10859 ( .DIN(n10412), .Q(n5050) );
  nnd2s1 U10860 ( .DIN1(n10413), .DIN2(n1602), .Q(n10406) );
  xor2s1 U10861 ( .DIN1(w1[14]), .DIN2(text_in_r[78]), .Q(n10413) );
  nnd2s1 U10862 ( .DIN1(n10414), .DIN2(n10415), .Q(N183) );
  nnd2s1 U10863 ( .DIN1(n10416), .DIN2(n1629), .Q(n10415) );
  xor2s1 U10864 ( .DIN1(n10417), .DIN2(n10418), .Q(n10416) );
  xor2s1 U10865 ( .DIN1(n10249), .DIN2(n10271), .Q(n10418) );
  xnr2s1 U10866 ( .DIN1(n10419), .DIN2(n5049), .Q(n10271) );
  hi1s1 U10867 ( .DIN(n10420), .Q(n5049) );
  xor2s1 U10868 ( .DIN1(n1492), .DIN2(n5027), .Q(n10417) );
  hi1s1 U10869 ( .DIN(n10411), .Q(n5027) );
  nnd2s1 U10870 ( .DIN1(n10421), .DIN2(n1601), .Q(n10414) );
  xor2s1 U10871 ( .DIN1(w1[13]), .DIN2(text_in_r[77]), .Q(n10421) );
  nnd2s1 U10872 ( .DIN1(n10422), .DIN2(n10423), .Q(N182) );
  nnd2s1 U10873 ( .DIN1(n10424), .DIN2(n1629), .Q(n10423) );
  xor2s1 U10874 ( .DIN1(n10425), .DIN2(n10426), .Q(n10424) );
  xor2s1 U10875 ( .DIN1(n10257), .DIN2(n10289), .Q(n10426) );
  hi1s1 U10876 ( .DIN(n10282), .Q(n10289) );
  xor2s1 U10877 ( .DIN1(n5025), .DIN2(n10427), .Q(n10282) );
  hi1s1 U10878 ( .DIN(n5048), .Q(n10427) );
  xor2s1 U10879 ( .DIN1(n10428), .DIN2(n10239), .Q(n10425) );
  xor2s1 U10880 ( .DIN1(n1493), .DIN2(n5026), .Q(n10428) );
  hi1s1 U10881 ( .DIN(n10419), .Q(n5026) );
  nnd2s1 U10882 ( .DIN1(n10429), .DIN2(n1601), .Q(n10422) );
  xor2s1 U10883 ( .DIN1(w1[12]), .DIN2(text_in_r[76]), .Q(n10429) );
  nnd3s1 U10884 ( .DIN1(n10430), .DIN2(n10431), .DIN3(n10432), .Q(N181) );
  nnd2s1 U10885 ( .DIN1(n1599), .DIN2(n10433), .Q(n10432) );
  xor2s1 U10886 ( .DIN1(w1[11]), .DIN2(text_in_r[75]), .Q(n10433) );
  nnd2s1 U10887 ( .DIN1(n10434), .DIN2(n10435), .Q(n10431) );
  nnd2s1 U10888 ( .DIN1(n10436), .DIN2(n10437), .Q(n10434) );
  nnd2s1 U10889 ( .DIN1(n10267), .DIN2(n10382), .Q(n10437) );
  nnd2s1 U10890 ( .DIN1(n10299), .DIN2(n10269), .Q(n10436) );
  nnd2s1 U10891 ( .DIN1(n10438), .DIN2(n10439), .Q(n10430) );
  nnd2s1 U10892 ( .DIN1(n10440), .DIN2(n10441), .Q(n10439) );
  nnd2s1 U10893 ( .DIN1(n10269), .DIN2(n10382), .Q(n10441) );
  and2s1 U10894 ( .DIN1(n10442), .DIN2(n1642), .Q(n10269) );
  nnd2s1 U10895 ( .DIN1(n10299), .DIN2(n10267), .Q(n10440) );
  nor2s1 U10896 ( .DIN1(n10442), .DIN2(n1594), .Q(n10267) );
  hi1s1 U10897 ( .DIN(n10382), .Q(n10299) );
  xor2s1 U10898 ( .DIN1(n5047), .DIN2(n10443), .Q(n10382) );
  hi1s1 U10899 ( .DIN(n10435), .Q(n10438) );
  xor2s1 U10900 ( .DIN1(n10444), .DIN2(n10239), .Q(n10435) );
  xor2s1 U10901 ( .DIN1(n5025), .DIN2(w1[11]), .Q(n10444) );
  nnd2s1 U10902 ( .DIN1(n10445), .DIN2(n10446), .Q(N180) );
  nnd2s1 U10903 ( .DIN1(n10447), .DIN2(n1630), .Q(n10446) );
  xor2s1 U10904 ( .DIN1(n10448), .DIN2(n10449), .Q(n10447) );
  xor2s1 U10905 ( .DIN1(n10450), .DIN2(n10309), .Q(n10449) );
  xnr2s1 U10906 ( .DIN1(n5046), .DIN2(n5023), .Q(n10309) );
  xor2s1 U10907 ( .DIN1(w1[10]), .DIN2(n5024), .Q(n10448) );
  nnd2s1 U10908 ( .DIN1(n10451), .DIN2(n1601), .Q(n10445) );
  xor2s1 U10909 ( .DIN1(w1[10]), .DIN2(text_in_r[74]), .Q(n10451) );
  nnd2s1 U10910 ( .DIN1(n10452), .DIN2(n10453), .Q(N179) );
  nnd2s1 U10911 ( .DIN1(n10454), .DIN2(n1626), .Q(n10453) );
  xor2s1 U10912 ( .DIN1(n10455), .DIN2(n10456), .Q(n10454) );
  xor2s1 U10913 ( .DIN1(n10239), .DIN2(n10457), .Q(n10456) );
  xnr2s1 U10914 ( .DIN1(w1[9]), .DIN2(n5023), .Q(n10457) );
  xnr2s1 U10915 ( .DIN1(n10317), .DIN2(n10300), .Q(n10455) );
  xor2s1 U10916 ( .DIN1(n5045), .DIN2(n5022), .Q(n10317) );
  nnd2s1 U10917 ( .DIN1(n10458), .DIN2(n1601), .Q(n10452) );
  xor2s1 U10918 ( .DIN1(w1[9]), .DIN2(text_in_r[73]), .Q(n10458) );
  nnd2s1 U10919 ( .DIN1(n10459), .DIN2(n10460), .Q(N178) );
  nnd2s1 U10920 ( .DIN1(n10461), .DIN2(n1630), .Q(n10460) );
  xor2s1 U10921 ( .DIN1(n10462), .DIN2(n10463), .Q(n10461) );
  xor2s1 U10922 ( .DIN1(n10239), .DIN2(n10308), .Q(n10463) );
  hi1s1 U10923 ( .DIN(n10324), .Q(n10239) );
  xnr2s1 U10924 ( .DIN1(n5052), .DIN2(n5029), .Q(n10324) );
  xor2s1 U10925 ( .DIN1(n1494), .DIN2(n5022), .Q(n10462) );
  nnd2s1 U10926 ( .DIN1(n10464), .DIN2(n1601), .Q(n10459) );
  xor2s1 U10927 ( .DIN1(w1[8]), .DIN2(text_in_r[72]), .Q(n10464) );
  nnd3s1 U10928 ( .DIN1(n10465), .DIN2(n10466), .DIN3(n10467), .Q(N169) );
  nnd2s1 U10929 ( .DIN1(n1599), .DIN2(n10468), .Q(n10467) );
  xor2s1 U10930 ( .DIN1(w1[7]), .DIN2(text_in_r[71]), .Q(n10468) );
  nnd2s1 U10931 ( .DIN1(n10469), .DIN2(n10470), .Q(n10466) );
  nnd2s1 U10932 ( .DIN1(n10471), .DIN2(n10472), .Q(n10469) );
  nnd2s1 U10933 ( .DIN1(n10335), .DIN2(n10473), .Q(n10472) );
  nnd2s1 U10934 ( .DIN1(n10276), .DIN2(n10337), .Q(n10471) );
  nnd2s1 U10935 ( .DIN1(n10474), .DIN2(n10475), .Q(n10465) );
  nnd2s1 U10936 ( .DIN1(n10476), .DIN2(n10477), .Q(n10475) );
  nnd2s1 U10937 ( .DIN1(n10337), .DIN2(n10473), .Q(n10477) );
  nor2s1 U10938 ( .DIN1(n5700), .DIN2(n1595), .Q(n10337) );
  nnd2s1 U10939 ( .DIN1(n10276), .DIN2(n10335), .Q(n10476) );
  and2s1 U10940 ( .DIN1(n5700), .DIN2(n1643), .Q(n10335) );
  hi1s1 U10941 ( .DIN(n10473), .Q(n10276) );
  xor2s1 U10942 ( .DIN1(n5701), .DIN2(n5076), .Q(n10473) );
  hi1s1 U10943 ( .DIN(n10241), .Q(n5076) );
  or3s1 U10944 ( .DIN1(n10478), .DIN2(n10479), .DIN3(n10480), .Q(n10241) );
  nnd4s1 U10945 ( .DIN1(n10481), .DIN2(n10482), .DIN3(n10483), .DIN4(n10484), 
        .Q(n10480) );
  and4s1 U10946 ( .DIN1(n10485), .DIN2(n10486), .DIN3(n10487), .DIN4(n10488), 
        .Q(n10484) );
  nnd2s1 U10947 ( .DIN1(n10489), .DIN2(n10490), .Q(n10487) );
  nnd2s1 U10948 ( .DIN1(n10491), .DIN2(n10492), .Q(n10486) );
  nnd4s1 U10949 ( .DIN1(n10493), .DIN2(n10494), .DIN3(n10495), .DIN4(n10496), 
        .Q(n10479) );
  nnd2s1 U10950 ( .DIN1(n10497), .DIN2(n10498), .Q(n10496) );
  nnd2s1 U10951 ( .DIN1(n10499), .DIN2(n10500), .Q(n10495) );
  nnd2s1 U10952 ( .DIN1(n10501), .DIN2(n10502), .Q(n10494) );
  nnd4s1 U10953 ( .DIN1(n10503), .DIN2(n10504), .DIN3(n10505), .DIN4(n10506), 
        .Q(n10478) );
  nnd2s1 U10954 ( .DIN1(n10507), .DIN2(n10508), .Q(n10506) );
  nnd2s1 U10955 ( .DIN1(n10509), .DIN2(n10510), .Q(n10508) );
  nnd2s1 U10956 ( .DIN1(n10511), .DIN2(n10512), .Q(n10505) );
  nnd2s1 U10957 ( .DIN1(n10513), .DIN2(n10514), .Q(n10512) );
  nnd2s1 U10958 ( .DIN1(n10515), .DIN2(n10516), .Q(n10504) );
  nnd2s1 U10959 ( .DIN1(n10517), .DIN2(n10518), .Q(n10516) );
  nnd2s1 U10960 ( .DIN1(n10519), .DIN2(n10520), .Q(n10503) );
  hi1s1 U10961 ( .DIN(n10470), .Q(n10474) );
  xnr2s1 U10962 ( .DIN1(n5052), .DIN2(n10521), .Q(n10470) );
  xnr2s1 U10963 ( .DIN1(w1[7]), .DIN2(n5028), .Q(n10521) );
  or3s1 U10964 ( .DIN1(n10522), .DIN2(n10523), .DIN3(n10524), .Q(n5028) );
  nnd4s1 U10965 ( .DIN1(n10525), .DIN2(n10526), .DIN3(n10527), .DIN4(n10528), 
        .Q(n10524) );
  and3s1 U10966 ( .DIN1(n10529), .DIN2(n10530), .DIN3(n10531), .Q(n10528) );
  nnd2s1 U10967 ( .DIN1(n10532), .DIN2(n10533), .Q(n10525) );
  nnd3s1 U10968 ( .DIN1(n10534), .DIN2(n10535), .DIN3(n10536), .Q(n10523) );
  or2s1 U10969 ( .DIN1(n10537), .DIN2(n10538), .Q(n10536) );
  or2s1 U10970 ( .DIN1(n10539), .DIN2(n10540), .Q(n10535) );
  nnd2s1 U10971 ( .DIN1(n10541), .DIN2(n10542), .Q(n10534) );
  nnd3s1 U10972 ( .DIN1(n10543), .DIN2(n10544), .DIN3(n10545), .Q(n10522) );
  nnd2s1 U10973 ( .DIN1(n10546), .DIN2(n10547), .Q(n10545) );
  nnd2s1 U10974 ( .DIN1(n10548), .DIN2(n10549), .Q(n10547) );
  nnd2s1 U10975 ( .DIN1(n10550), .DIN2(n10551), .Q(n10544) );
  nnd2s1 U10976 ( .DIN1(n10552), .DIN2(n10553), .Q(n10551) );
  hi1s1 U10977 ( .DIN(n10554), .Q(n10553) );
  nnd2s1 U10978 ( .DIN1(n10555), .DIN2(n10556), .Q(n10543) );
  nnd2s1 U10979 ( .DIN1(n10557), .DIN2(n10558), .Q(n10556) );
  nor3s1 U10980 ( .DIN1(n10559), .DIN2(n10560), .DIN3(n10561), .Q(n5052) );
  nnd4s1 U10981 ( .DIN1(n10562), .DIN2(n10563), .DIN3(n10564), .DIN4(n10565), 
        .Q(n10561) );
  and4s1 U10982 ( .DIN1(n10566), .DIN2(n10567), .DIN3(n10568), .DIN4(n10569), 
        .Q(n10565) );
  nnd2s1 U10983 ( .DIN1(n10570), .DIN2(n10571), .Q(n10568) );
  nnd2s1 U10984 ( .DIN1(n10572), .DIN2(n10573), .Q(n10567) );
  nnd4s1 U10985 ( .DIN1(n10574), .DIN2(n10575), .DIN3(n10576), .DIN4(n10577), 
        .Q(n10560) );
  nnd2s1 U10986 ( .DIN1(n10578), .DIN2(n10579), .Q(n10577) );
  nnd2s1 U10987 ( .DIN1(n10580), .DIN2(n10581), .Q(n10576) );
  nnd2s1 U10988 ( .DIN1(n10582), .DIN2(n10583), .Q(n10575) );
  nnd4s1 U10989 ( .DIN1(n10584), .DIN2(n10585), .DIN3(n10586), .DIN4(n10587), 
        .Q(n10559) );
  nnd2s1 U10990 ( .DIN1(n10588), .DIN2(n10589), .Q(n10587) );
  nnd2s1 U10991 ( .DIN1(n10590), .DIN2(n10591), .Q(n10589) );
  nnd2s1 U10992 ( .DIN1(n10592), .DIN2(n10593), .Q(n10586) );
  nnd2s1 U10993 ( .DIN1(n10594), .DIN2(n10595), .Q(n10593) );
  nnd2s1 U10994 ( .DIN1(n10596), .DIN2(n10597), .Q(n10585) );
  nnd2s1 U10995 ( .DIN1(n10598), .DIN2(n10599), .Q(n10597) );
  nnd2s1 U10996 ( .DIN1(n10600), .DIN2(n10601), .Q(n10584) );
  nnd3s1 U10997 ( .DIN1(n10602), .DIN2(n10603), .DIN3(n10604), .Q(N168) );
  nnd2s1 U10998 ( .DIN1(n1599), .DIN2(n10605), .Q(n10604) );
  xor2s1 U10999 ( .DIN1(w1[6]), .DIN2(text_in_r[70]), .Q(n10605) );
  nnd2s1 U11000 ( .DIN1(n10606), .DIN2(n10607), .Q(n10603) );
  nnd2s1 U11001 ( .DIN1(n10608), .DIN2(n10609), .Q(n10606) );
  nnd2s1 U11002 ( .DIN1(n10351), .DIN2(n10610), .Q(n10609) );
  nnd2s1 U11003 ( .DIN1(n10240), .DIN2(n10353), .Q(n10608) );
  nnd2s1 U11004 ( .DIN1(n10611), .DIN2(n10612), .Q(n10602) );
  nnd2s1 U11005 ( .DIN1(n10613), .DIN2(n10614), .Q(n10612) );
  nnd2s1 U11006 ( .DIN1(n10353), .DIN2(n10610), .Q(n10614) );
  nor2s1 U11007 ( .DIN1(n10615), .DIN2(n1596), .Q(n10353) );
  nnd2s1 U11008 ( .DIN1(n10240), .DIN2(n10351), .Q(n10613) );
  nor2s1 U11009 ( .DIN1(n5699), .DIN2(n1595), .Q(n10351) );
  hi1s1 U11010 ( .DIN(n10615), .Q(n5699) );
  hi1s1 U11011 ( .DIN(n10610), .Q(n10240) );
  xor2s1 U11012 ( .DIN1(n5700), .DIN2(n10616), .Q(n10610) );
  hi1s1 U11013 ( .DIN(n5075), .Q(n10616) );
  or3s1 U11014 ( .DIN1(n10617), .DIN2(n10618), .DIN3(n10619), .Q(n5075) );
  nnd4s1 U11015 ( .DIN1(n10620), .DIN2(n10621), .DIN3(n10622), .DIN4(n10623), 
        .Q(n10619) );
  and3s1 U11016 ( .DIN1(n10624), .DIN2(n10625), .DIN3(n10626), .Q(n10623) );
  nnd2s1 U11017 ( .DIN1(n10627), .DIN2(n10499), .Q(n10621) );
  nnd2s1 U11018 ( .DIN1(n10490), .DIN2(n10628), .Q(n10620) );
  nnd3s1 U11019 ( .DIN1(n10629), .DIN2(n10630), .DIN3(n10631), .Q(n10618) );
  or2s1 U11020 ( .DIN1(n10632), .DIN2(n10633), .Q(n10631) );
  or2s1 U11021 ( .DIN1(n10514), .DIN2(n10634), .Q(n10630) );
  nnd2s1 U11022 ( .DIN1(n10515), .DIN2(n10635), .Q(n10629) );
  nnd3s1 U11023 ( .DIN1(n10636), .DIN2(n10637), .DIN3(n10638), .Q(n10617) );
  nnd2s1 U11024 ( .DIN1(n10639), .DIN2(n10640), .Q(n10638) );
  nnd2s1 U11025 ( .DIN1(n10641), .DIN2(n10642), .Q(n10640) );
  nnd2s1 U11026 ( .DIN1(n10643), .DIN2(n10644), .Q(n10637) );
  nnd2s1 U11027 ( .DIN1(n10645), .DIN2(n10646), .Q(n10644) );
  nnd2s1 U11028 ( .DIN1(n10491), .DIN2(n10647), .Q(n10636) );
  nnd2s1 U11029 ( .DIN1(n10648), .DIN2(n10649), .Q(n10647) );
  hi1s1 U11030 ( .DIN(n10650), .Q(n10649) );
  or3s1 U11031 ( .DIN1(n10651), .DIN2(n10652), .DIN3(n10653), .Q(n5700) );
  nnd4s1 U11032 ( .DIN1(n10654), .DIN2(n10655), .DIN3(n10656), .DIN4(n10657), 
        .Q(n10653) );
  and3s1 U11033 ( .DIN1(n10658), .DIN2(n10659), .DIN3(n10660), .Q(n10657) );
  nnd2s1 U11034 ( .DIN1(n10661), .DIN2(n10662), .Q(n10655) );
  nnd2s1 U11035 ( .DIN1(n10663), .DIN2(n10664), .Q(n10654) );
  nnd3s1 U11036 ( .DIN1(n10665), .DIN2(n10666), .DIN3(n10667), .Q(n10652) );
  or2s1 U11037 ( .DIN1(n10668), .DIN2(n10669), .Q(n10667) );
  or2s1 U11038 ( .DIN1(n10670), .DIN2(n10671), .Q(n10666) );
  nnd2s1 U11039 ( .DIN1(n10672), .DIN2(n10673), .Q(n10665) );
  nnd3s1 U11040 ( .DIN1(n10674), .DIN2(n10675), .DIN3(n10676), .Q(n10651) );
  nnd2s1 U11041 ( .DIN1(n10677), .DIN2(n10678), .Q(n10676) );
  nnd2s1 U11042 ( .DIN1(n10679), .DIN2(n10680), .Q(n10678) );
  nnd2s1 U11043 ( .DIN1(n10681), .DIN2(n10682), .Q(n10675) );
  nnd2s1 U11044 ( .DIN1(n10683), .DIN2(n10684), .Q(n10682) );
  nnd2s1 U11045 ( .DIN1(n10685), .DIN2(n10686), .Q(n10674) );
  nnd2s1 U11046 ( .DIN1(n10687), .DIN2(n10688), .Q(n10686) );
  hi1s1 U11047 ( .DIN(n10689), .Q(n10688) );
  hi1s1 U11048 ( .DIN(n10607), .Q(n10611) );
  xor2s1 U11049 ( .DIN1(n5051), .DIN2(n10690), .Q(n10607) );
  xor2s1 U11050 ( .DIN1(n1542), .DIN2(n10411), .Q(n10690) );
  or3s1 U11051 ( .DIN1(n10691), .DIN2(n10692), .DIN3(n10693), .Q(n10411) );
  nnd4s1 U11052 ( .DIN1(n10694), .DIN2(n10695), .DIN3(n10531), .DIN4(n10696), 
        .Q(n10693) );
  and4s1 U11053 ( .DIN1(n10697), .DIN2(n10698), .DIN3(n10699), .DIN4(n10700), 
        .Q(n10696) );
  nnd2s1 U11054 ( .DIN1(n10532), .DIN2(n10701), .Q(n10700) );
  nnd2s1 U11055 ( .DIN1(n10546), .DIN2(n10702), .Q(n10699) );
  nnd2s1 U11056 ( .DIN1(n10703), .DIN2(n10555), .Q(n10698) );
  nor2s1 U11057 ( .DIN1(n10704), .DIN2(n10705), .Q(n10531) );
  nnd4s1 U11058 ( .DIN1(n10706), .DIN2(n10707), .DIN3(n10708), .DIN4(n10709), 
        .Q(n10705) );
  nnd2s1 U11059 ( .DIN1(n10710), .DIN2(n10711), .Q(n10709) );
  nnd3s1 U11060 ( .DIN1(n10712), .DIN2(n10558), .DIN3(n10713), .Q(n10711) );
  nnd2s1 U11061 ( .DIN1(n10714), .DIN2(n10715), .Q(n10708) );
  nnd2s1 U11062 ( .DIN1(n10703), .DIN2(n10716), .Q(n10707) );
  nnd2s1 U11063 ( .DIN1(n10717), .DIN2(n10701), .Q(n10706) );
  nnd4s1 U11064 ( .DIN1(n10718), .DIN2(n10719), .DIN3(n10720), .DIN4(n10721), 
        .Q(n10704) );
  nnd2s1 U11065 ( .DIN1(n10722), .DIN2(n10723), .Q(n10721) );
  nnd2s1 U11066 ( .DIN1(n10724), .DIN2(n10725), .Q(n10723) );
  nnd2s1 U11067 ( .DIN1(n10702), .DIN2(n10726), .Q(n10720) );
  nnd2s1 U11068 ( .DIN1(n10727), .DIN2(n10728), .Q(n10726) );
  nnd2s1 U11069 ( .DIN1(n10729), .DIN2(n10730), .Q(n10719) );
  nnd2s1 U11070 ( .DIN1(n10731), .DIN2(n10549), .Q(n10730) );
  nnd2s1 U11071 ( .DIN1(n10732), .DIN2(n10733), .Q(n10718) );
  nnd2s1 U11072 ( .DIN1(n10558), .DIN2(n10734), .Q(n10733) );
  nnd4s1 U11073 ( .DIN1(n10735), .DIN2(n10736), .DIN3(n10737), .DIN4(n10738), 
        .Q(n10692) );
  or2s1 U11074 ( .DIN1(n10739), .DIN2(n10740), .Q(n10738) );
  nnd2s1 U11075 ( .DIN1(n10717), .DIN2(n10741), .Q(n10737) );
  nnd2s1 U11076 ( .DIN1(n10742), .DIN2(n10743), .Q(n10736) );
  nnd2s1 U11077 ( .DIN1(n10714), .DIN2(n10744), .Q(n10735) );
  nnd4s1 U11078 ( .DIN1(n10745), .DIN2(n10746), .DIN3(n10747), .DIN4(n10748), 
        .Q(n10691) );
  nnd2s1 U11079 ( .DIN1(n10749), .DIN2(n10750), .Q(n10748) );
  nnd2s1 U11080 ( .DIN1(n10712), .DIN2(n10751), .Q(n10750) );
  nnd2s1 U11081 ( .DIN1(n10752), .DIN2(n10753), .Q(n10747) );
  nnd2s1 U11082 ( .DIN1(n10548), .DIN2(n10754), .Q(n10753) );
  nnd2s1 U11083 ( .DIN1(n10541), .DIN2(n10755), .Q(n10746) );
  nnd2s1 U11084 ( .DIN1(n10756), .DIN2(n10757), .Q(n10755) );
  nnd2s1 U11085 ( .DIN1(n10758), .DIN2(n10759), .Q(n10745) );
  or3s1 U11086 ( .DIN1(n10760), .DIN2(n10761), .DIN3(n10762), .Q(n5051) );
  nnd4s1 U11087 ( .DIN1(n10763), .DIN2(n10764), .DIN3(n10765), .DIN4(n10766), 
        .Q(n10762) );
  and3s1 U11088 ( .DIN1(n10767), .DIN2(n10768), .DIN3(n10769), .Q(n10766) );
  nnd2s1 U11089 ( .DIN1(n10770), .DIN2(n10580), .Q(n10764) );
  nnd2s1 U11090 ( .DIN1(n10571), .DIN2(n10771), .Q(n10763) );
  nnd3s1 U11091 ( .DIN1(n10772), .DIN2(n10773), .DIN3(n10774), .Q(n10761) );
  or2s1 U11092 ( .DIN1(n10775), .DIN2(n10776), .Q(n10774) );
  or2s1 U11093 ( .DIN1(n10595), .DIN2(n10777), .Q(n10773) );
  nnd2s1 U11094 ( .DIN1(n10596), .DIN2(n10778), .Q(n10772) );
  nnd3s1 U11095 ( .DIN1(n10779), .DIN2(n10780), .DIN3(n10781), .Q(n10760) );
  nnd2s1 U11096 ( .DIN1(n10782), .DIN2(n10783), .Q(n10781) );
  nnd2s1 U11097 ( .DIN1(n10784), .DIN2(n10785), .Q(n10783) );
  nnd2s1 U11098 ( .DIN1(n10786), .DIN2(n10787), .Q(n10780) );
  nnd2s1 U11099 ( .DIN1(n10788), .DIN2(n10789), .Q(n10787) );
  nnd2s1 U11100 ( .DIN1(n10572), .DIN2(n10790), .Q(n10779) );
  nnd2s1 U11101 ( .DIN1(n10791), .DIN2(n10792), .Q(n10790) );
  hi1s1 U11102 ( .DIN(n10793), .Q(n10792) );
  nnd2s1 U11103 ( .DIN1(n10794), .DIN2(n10795), .Q(N167) );
  nnd2s1 U11104 ( .DIN1(n10796), .DIN2(n1631), .Q(n10795) );
  xor2s1 U11105 ( .DIN1(n10797), .DIN2(n10798), .Q(n10796) );
  xnr2s1 U11106 ( .DIN1(n5698), .DIN2(n10249), .Q(n10798) );
  xnr2s1 U11107 ( .DIN1(n10615), .DIN2(n5074), .Q(n10249) );
  nor3s1 U11108 ( .DIN1(n10799), .DIN2(n10800), .DIN3(n10801), .Q(n5074) );
  nnd4s1 U11109 ( .DIN1(n10802), .DIN2(n10803), .DIN3(n10626), .DIN4(n10804), 
        .Q(n10801) );
  and4s1 U11110 ( .DIN1(n10805), .DIN2(n10806), .DIN3(n10807), .DIN4(n10488), 
        .Q(n10804) );
  nnd2s1 U11111 ( .DIN1(n10808), .DIN2(n10643), .Q(n10488) );
  nnd2s1 U11112 ( .DIN1(n10639), .DIN2(n10809), .Q(n10807) );
  nnd2s1 U11113 ( .DIN1(n10810), .DIN2(n10492), .Q(n10806) );
  nor2s1 U11114 ( .DIN1(n10811), .DIN2(n10812), .Q(n10626) );
  nnd4s1 U11115 ( .DIN1(n10813), .DIN2(n10814), .DIN3(n10815), .DIN4(n10816), 
        .Q(n10812) );
  or2s1 U11116 ( .DIN1(n10817), .DIN2(n10818), .Q(n10816) );
  nnd2s1 U11117 ( .DIN1(n10810), .DIN2(n10819), .Q(n10815) );
  nnd2s1 U11118 ( .DIN1(n10808), .DIN2(n10490), .Q(n10814) );
  nnd2s1 U11119 ( .DIN1(n10502), .DIN2(n10820), .Q(n10813) );
  nnd4s1 U11120 ( .DIN1(n10821), .DIN2(n10822), .DIN3(n10823), .DIN4(n10824), 
        .Q(n10811) );
  nnd2s1 U11121 ( .DIN1(n10501), .DIN2(n10825), .Q(n10824) );
  nnd2s1 U11122 ( .DIN1(n10645), .DIN2(n10826), .Q(n10825) );
  nnd2s1 U11123 ( .DIN1(n10827), .DIN2(n10828), .Q(n10823) );
  nnd2s1 U11124 ( .DIN1(n10641), .DIN2(n10829), .Q(n10828) );
  nnd2s1 U11125 ( .DIN1(n10809), .DIN2(n10830), .Q(n10822) );
  nnd2s1 U11126 ( .DIN1(n10831), .DIN2(n10832), .Q(n10830) );
  nnd2s1 U11127 ( .DIN1(n10511), .DIN2(n10833), .Q(n10821) );
  nnd3s1 U11128 ( .DIN1(n10834), .DIN2(n10645), .DIN3(n10835), .Q(n10833) );
  nnd4s1 U11129 ( .DIN1(n10836), .DIN2(n10837), .DIN3(n10838), .DIN4(n10839), 
        .Q(n10800) );
  nnd2s1 U11130 ( .DIN1(n10840), .DIN2(n10841), .Q(n10839) );
  nnd2s1 U11131 ( .DIN1(n10502), .DIN2(n10842), .Q(n10838) );
  nnd2s1 U11132 ( .DIN1(n10489), .DIN2(n10843), .Q(n10837) );
  nnd2s1 U11133 ( .DIN1(n10627), .DIN2(n10820), .Q(n10836) );
  nnd4s1 U11134 ( .DIN1(n10844), .DIN2(n10845), .DIN3(n10846), .DIN4(n10847), 
        .Q(n10799) );
  nnd2s1 U11135 ( .DIN1(n10519), .DIN2(n10848), .Q(n10847) );
  nnd2s1 U11136 ( .DIN1(n10642), .DIN2(n10849), .Q(n10848) );
  nnd2s1 U11137 ( .DIN1(n10850), .DIN2(n10851), .Q(n10846) );
  nnd2s1 U11138 ( .DIN1(n10515), .DIN2(n10852), .Q(n10845) );
  nnd2s1 U11139 ( .DIN1(n10853), .DIN2(n10510), .Q(n10852) );
  nnd2s1 U11140 ( .DIN1(n10499), .DIN2(n10854), .Q(n10844) );
  or3s1 U11141 ( .DIN1(n10855), .DIN2(n10856), .DIN3(n10857), .Q(n10615) );
  nnd4s1 U11142 ( .DIN1(n10858), .DIN2(n10859), .DIN3(n10660), .DIN4(n10860), 
        .Q(n10857) );
  and4s1 U11143 ( .DIN1(n10861), .DIN2(n10862), .DIN3(n10863), .DIN4(n10864), 
        .Q(n10860) );
  nnd2s1 U11144 ( .DIN1(n10677), .DIN2(n10865), .Q(n10863) );
  nnd2s1 U11145 ( .DIN1(n10866), .DIN2(n10867), .Q(n10862) );
  nor2s1 U11146 ( .DIN1(n10868), .DIN2(n10869), .Q(n10660) );
  nnd4s1 U11147 ( .DIN1(n10870), .DIN2(n10871), .DIN3(n10872), .DIN4(n10873), 
        .Q(n10869) );
  or2s1 U11148 ( .DIN1(n10874), .DIN2(n10875), .Q(n10873) );
  nnd2s1 U11149 ( .DIN1(n10866), .DIN2(n10876), .Q(n10872) );
  nnd2s1 U11150 ( .DIN1(n10877), .DIN2(n10663), .Q(n10871) );
  nnd2s1 U11151 ( .DIN1(n10878), .DIN2(n10879), .Q(n10870) );
  nnd4s1 U11152 ( .DIN1(n10880), .DIN2(n10881), .DIN3(n10882), .DIN4(n10883), 
        .Q(n10868) );
  nnd2s1 U11153 ( .DIN1(n10884), .DIN2(n10885), .Q(n10883) );
  nnd2s1 U11154 ( .DIN1(n10683), .DIN2(n10886), .Q(n10885) );
  nnd2s1 U11155 ( .DIN1(n10887), .DIN2(n10888), .Q(n10882) );
  nnd2s1 U11156 ( .DIN1(n10679), .DIN2(n10889), .Q(n10888) );
  nnd2s1 U11157 ( .DIN1(n10865), .DIN2(n10890), .Q(n10881) );
  nnd2s1 U11158 ( .DIN1(n10891), .DIN2(n10892), .Q(n10890) );
  nnd2s1 U11159 ( .DIN1(n10893), .DIN2(n10894), .Q(n10880) );
  nnd3s1 U11160 ( .DIN1(n10895), .DIN2(n10683), .DIN3(n10896), .Q(n10894) );
  nnd4s1 U11161 ( .DIN1(n10897), .DIN2(n10898), .DIN3(n10899), .DIN4(n10900), 
        .Q(n10856) );
  nnd2s1 U11162 ( .DIN1(n10901), .DIN2(n10902), .Q(n10900) );
  nnd2s1 U11163 ( .DIN1(n10878), .DIN2(n10903), .Q(n10899) );
  nnd2s1 U11164 ( .DIN1(n10904), .DIN2(n10905), .Q(n10898) );
  nnd2s1 U11165 ( .DIN1(n10661), .DIN2(n10879), .Q(n10897) );
  nnd4s1 U11166 ( .DIN1(n10906), .DIN2(n10907), .DIN3(n10908), .DIN4(n10909), 
        .Q(n10855) );
  nnd2s1 U11167 ( .DIN1(n10910), .DIN2(n10911), .Q(n10909) );
  nnd2s1 U11168 ( .DIN1(n10680), .DIN2(n10912), .Q(n10911) );
  nnd2s1 U11169 ( .DIN1(n10913), .DIN2(n10914), .Q(n10908) );
  nnd2s1 U11170 ( .DIN1(n10672), .DIN2(n10915), .Q(n10907) );
  nnd2s1 U11171 ( .DIN1(n10916), .DIN2(n10917), .Q(n10915) );
  nnd2s1 U11172 ( .DIN1(n10662), .DIN2(n10918), .Q(n10906) );
  xor2s1 U11173 ( .DIN1(n10412), .DIN2(n10919), .Q(n10797) );
  xor2s1 U11174 ( .DIN1(n1495), .DIN2(n10419), .Q(n10919) );
  or3s1 U11175 ( .DIN1(n10920), .DIN2(n10921), .DIN3(n10922), .Q(n10419) );
  nnd4s1 U11176 ( .DIN1(n10923), .DIN2(n10924), .DIN3(n10925), .DIN4(n10926), 
        .Q(n10922) );
  and4s1 U11177 ( .DIN1(n10927), .DIN2(n10928), .DIN3(n10929), .DIN4(n10930), 
        .Q(n10926) );
  nnd2s1 U11178 ( .DIN1(n10532), .DIN2(n10931), .Q(n10930) );
  nnd2s1 U11179 ( .DIN1(n10932), .DIN2(n10933), .Q(n10931) );
  nnd2s1 U11180 ( .DIN1(n10934), .DIN2(n10935), .Q(n10929) );
  nnd2s1 U11181 ( .DIN1(n10548), .DIN2(n10734), .Q(n10935) );
  nnd2s1 U11182 ( .DIN1(n10555), .DIN2(n10936), .Q(n10928) );
  nnd2s1 U11183 ( .DIN1(n10937), .DIN2(n10938), .Q(n10927) );
  nnd2s1 U11184 ( .DIN1(n10939), .DIN2(n10940), .Q(n10938) );
  nnd2s1 U11185 ( .DIN1(n10714), .DIN2(n10941), .Q(n10925) );
  nnd2s1 U11186 ( .DIN1(n10533), .DIN2(n10759), .Q(n10924) );
  nnd2s1 U11187 ( .DIN1(n10702), .DIN2(n10741), .Q(n10923) );
  nnd3s1 U11188 ( .DIN1(n10694), .DIN2(n10942), .DIN3(n10529), .Q(n10921) );
  nor4s1 U11189 ( .DIN1(n10943), .DIN2(n10944), .DIN3(n10945), .DIN4(n10946), 
        .Q(n10529) );
  nnd4s1 U11190 ( .DIN1(n10947), .DIN2(n10948), .DIN3(n10949), .DIN4(n10950), 
        .Q(n10946) );
  nnd2s1 U11191 ( .DIN1(n10752), .DIN2(n10951), .Q(n10950) );
  nnd2s1 U11192 ( .DIN1(n10532), .DIN2(n10934), .Q(n10949) );
  nnd2s1 U11193 ( .DIN1(n10703), .DIN2(n10550), .Q(n10948) );
  nnd2s1 U11194 ( .DIN1(n10729), .DIN2(n10952), .Q(n10947) );
  nnd3s1 U11195 ( .DIN1(n10953), .DIN2(n10954), .DIN3(n10955), .Q(n10945) );
  nnd2s1 U11196 ( .DIN1(n10732), .DIN2(n10956), .Q(n10955) );
  nnd2s1 U11197 ( .DIN1(n10957), .DIN2(n10958), .Q(n10956) );
  nnd2s1 U11198 ( .DIN1(n10758), .DIN2(n10959), .Q(n10954) );
  nnd2s1 U11199 ( .DIN1(n10960), .DIN2(n10961), .Q(n10959) );
  nnd2s1 U11200 ( .DIN1(n10710), .DIN2(n10962), .Q(n10953) );
  nnd2s1 U11201 ( .DIN1(n10963), .DIN2(n10754), .Q(n10962) );
  nor2s1 U11202 ( .DIN1(n10731), .DIN2(n10964), .Q(n10944) );
  and2s1 U11203 ( .DIN1(n10716), .DIN2(n10965), .Q(n10943) );
  nnd3s1 U11204 ( .DIN1(n10558), .DIN2(n10966), .DIN3(n10548), .Q(n10965) );
  nor3s1 U11205 ( .DIN1(n10967), .DIN2(n10968), .DIN3(n10969), .Q(n10694) );
  nnd4s1 U11206 ( .DIN1(n10970), .DIN2(n10971), .DIN3(n10530), .DIN4(n10972), 
        .Q(n10969) );
  and3s1 U11207 ( .DIN1(n10973), .DIN2(n10974), .DIN3(n10975), .Q(n10972) );
  nnd2s1 U11208 ( .DIN1(n10703), .DIN2(n10701), .Q(n10974) );
  nnd2s1 U11209 ( .DIN1(n10752), .DIN2(n10702), .Q(n10973) );
  nor2s1 U11210 ( .DIN1(n10976), .DIN2(n10977), .Q(n10530) );
  nnd4s1 U11211 ( .DIN1(n10978), .DIN2(n10979), .DIN3(n10980), .DIN4(n10981), 
        .Q(n10977) );
  nnd2s1 U11212 ( .DIN1(n10546), .DIN2(n10982), .Q(n10981) );
  nnd2s1 U11213 ( .DIN1(n10541), .DIN2(n10983), .Q(n10980) );
  nnd2s1 U11214 ( .DIN1(n10934), .DIN2(n10941), .Q(n10979) );
  nnd2s1 U11215 ( .DIN1(n10710), .DIN2(n10722), .Q(n10978) );
  nnd4s1 U11216 ( .DIN1(n10984), .DIN2(n10985), .DIN3(n10986), .DIN4(n10987), 
        .Q(n10976) );
  nnd2s1 U11217 ( .DIN1(n10742), .DIN2(n10988), .Q(n10987) );
  nnd2s1 U11218 ( .DIN1(n10932), .DIN2(n10940), .Q(n10988) );
  nnd2s1 U11219 ( .DIN1(n10532), .DIN2(n10983), .Q(n10986) );
  nnd2s1 U11220 ( .DIN1(n10732), .DIN2(n10989), .Q(n10985) );
  nnd2s1 U11221 ( .DIN1(n10557), .DIN2(n10731), .Q(n10989) );
  nnd2s1 U11222 ( .DIN1(n10990), .DIN2(n10991), .Q(n10984) );
  nnd3s1 U11223 ( .DIN1(n10739), .DIN2(n10933), .DIN3(n10992), .Q(n10991) );
  nnd3s1 U11224 ( .DIN1(n10993), .DIN2(n10994), .DIN3(n10995), .Q(n10968) );
  nnd2s1 U11225 ( .DIN1(n10996), .DIN2(n10717), .Q(n10995) );
  nnd2s1 U11226 ( .DIN1(n10742), .DIN2(n10997), .Q(n10994) );
  nnd3s1 U11227 ( .DIN1(n10998), .DIN2(n10728), .DIN3(n10540), .Q(n10997) );
  nor2s1 U11228 ( .DIN1(n10550), .DIN2(n10749), .Q(n10540) );
  nnd2s1 U11229 ( .DIN1(n10990), .DIN2(n10550), .Q(n10993) );
  nnd3s1 U11230 ( .DIN1(n10999), .DIN2(n11000), .DIN3(n11001), .Q(n10967) );
  nnd2s1 U11231 ( .DIN1(n10546), .DIN2(n11002), .Q(n11001) );
  nnd2s1 U11232 ( .DIN1(n11003), .DIN2(n10539), .Q(n11002) );
  nnd2s1 U11233 ( .DIN1(n10758), .DIN2(n11004), .Q(n11000) );
  nnd2s1 U11234 ( .DIN1(n10754), .DIN2(n10958), .Q(n11004) );
  nnd2s1 U11235 ( .DIN1(n10533), .DIN2(n11005), .Q(n10999) );
  nnd2s1 U11236 ( .DIN1(n10731), .DIN2(n10958), .Q(n11005) );
  nnd3s1 U11237 ( .DIN1(n11006), .DIN2(n11007), .DIN3(n11008), .Q(n10920) );
  or3s1 U11238 ( .DIN1(n11009), .DIN2(n11010), .DIN3(n11011), .Q(n10412) );
  nnd4s1 U11239 ( .DIN1(n11012), .DIN2(n11013), .DIN3(n10769), .DIN4(n11014), 
        .Q(n11011) );
  and4s1 U11240 ( .DIN1(n11015), .DIN2(n11016), .DIN3(n11017), .DIN4(n10569), 
        .Q(n11014) );
  nnd2s1 U11241 ( .DIN1(n11018), .DIN2(n10786), .Q(n10569) );
  nnd2s1 U11242 ( .DIN1(n10782), .DIN2(n11019), .Q(n11017) );
  nnd2s1 U11243 ( .DIN1(n11020), .DIN2(n10573), .Q(n11016) );
  nor2s1 U11244 ( .DIN1(n11021), .DIN2(n11022), .Q(n10769) );
  nnd4s1 U11245 ( .DIN1(n11023), .DIN2(n11024), .DIN3(n11025), .DIN4(n11026), 
        .Q(n11022) );
  or2s1 U11246 ( .DIN1(n11027), .DIN2(n11028), .Q(n11026) );
  nnd2s1 U11247 ( .DIN1(n11020), .DIN2(n11029), .Q(n11025) );
  nnd2s1 U11248 ( .DIN1(n11018), .DIN2(n10571), .Q(n11024) );
  nnd2s1 U11249 ( .DIN1(n10583), .DIN2(n11030), .Q(n11023) );
  nnd4s1 U11250 ( .DIN1(n11031), .DIN2(n11032), .DIN3(n11033), .DIN4(n11034), 
        .Q(n11021) );
  nnd2s1 U11251 ( .DIN1(n10582), .DIN2(n11035), .Q(n11034) );
  nnd2s1 U11252 ( .DIN1(n10788), .DIN2(n11036), .Q(n11035) );
  nnd2s1 U11253 ( .DIN1(n11037), .DIN2(n11038), .Q(n11033) );
  nnd2s1 U11254 ( .DIN1(n10784), .DIN2(n11039), .Q(n11038) );
  nnd2s1 U11255 ( .DIN1(n11019), .DIN2(n11040), .Q(n11032) );
  nnd2s1 U11256 ( .DIN1(n11041), .DIN2(n11042), .Q(n11040) );
  nnd2s1 U11257 ( .DIN1(n10592), .DIN2(n11043), .Q(n11031) );
  nnd3s1 U11258 ( .DIN1(n11044), .DIN2(n10788), .DIN3(n11045), .Q(n11043) );
  nnd4s1 U11259 ( .DIN1(n11046), .DIN2(n11047), .DIN3(n11048), .DIN4(n11049), 
        .Q(n11010) );
  nnd2s1 U11260 ( .DIN1(n11050), .DIN2(n11051), .Q(n11049) );
  nnd2s1 U11261 ( .DIN1(n10583), .DIN2(n11052), .Q(n11048) );
  nnd2s1 U11262 ( .DIN1(n10570), .DIN2(n11053), .Q(n11047) );
  nnd2s1 U11263 ( .DIN1(n10770), .DIN2(n11030), .Q(n11046) );
  nnd4s1 U11264 ( .DIN1(n11054), .DIN2(n11055), .DIN3(n11056), .DIN4(n11057), 
        .Q(n11009) );
  nnd2s1 U11265 ( .DIN1(n10600), .DIN2(n11058), .Q(n11057) );
  nnd2s1 U11266 ( .DIN1(n10785), .DIN2(n11059), .Q(n11058) );
  nnd2s1 U11267 ( .DIN1(n11060), .DIN2(n11061), .Q(n11056) );
  nnd2s1 U11268 ( .DIN1(n10596), .DIN2(n11062), .Q(n11055) );
  nnd2s1 U11269 ( .DIN1(n11063), .DIN2(n10591), .Q(n11062) );
  nnd2s1 U11270 ( .DIN1(n10580), .DIN2(n11064), .Q(n11054) );
  nnd2s1 U11271 ( .DIN1(n11065), .DIN2(n1601), .Q(n10794) );
  xor2s1 U11272 ( .DIN1(w1[5]), .DIN2(text_in_r[69]), .Q(n11065) );
  nnd2s1 U11273 ( .DIN1(n11066), .DIN2(n11067), .Q(N166) );
  nnd2s1 U11274 ( .DIN1(n11068), .DIN2(n1631), .Q(n11067) );
  xor2s1 U11275 ( .DIN1(n11069), .DIN2(n11070), .Q(n11068) );
  xor2s1 U11276 ( .DIN1(n11071), .DIN2(n11072), .Q(n11070) );
  xnr2s1 U11277 ( .DIN1(n5425), .DIN2(n10257), .Q(n11072) );
  xnr2s1 U11278 ( .DIN1(n5698), .DIN2(n5073), .Q(n10257) );
  hi1s1 U11279 ( .DIN(n10358), .Q(n5073) );
  or3s1 U11280 ( .DIN1(n11073), .DIN2(n11074), .DIN3(n11075), .Q(n10358) );
  nnd4s1 U11281 ( .DIN1(n10802), .DIN2(n11076), .DIN3(n10624), .DIN4(n11077), 
        .Q(n11075) );
  and3s1 U11282 ( .DIN1(n11078), .DIN2(n11079), .DIN3(n11080), .Q(n11077) );
  nor4s1 U11283 ( .DIN1(n11081), .DIN2(n11082), .DIN3(n11083), .DIN4(n11084), 
        .Q(n10624) );
  nnd4s1 U11284 ( .DIN1(n11085), .DIN2(n11086), .DIN3(n11087), .DIN4(n11088), 
        .Q(n11084) );
  nnd2s1 U11285 ( .DIN1(n10627), .DIN2(n10497), .Q(n11088) );
  nnd2s1 U11286 ( .DIN1(n10810), .DIN2(n11089), .Q(n11086) );
  nnd2s1 U11287 ( .DIN1(n10827), .DIN2(n10498), .Q(n11085) );
  nnd3s1 U11288 ( .DIN1(n11090), .DIN2(n11091), .DIN3(n11092), .Q(n11083) );
  nnd2s1 U11289 ( .DIN1(n10840), .DIN2(n11093), .Q(n11092) );
  nnd2s1 U11290 ( .DIN1(n11094), .DIN2(n10513), .Q(n11093) );
  nnd2s1 U11291 ( .DIN1(n10511), .DIN2(n11095), .Q(n11091) );
  nnd2s1 U11292 ( .DIN1(n11096), .DIN2(n10849), .Q(n11095) );
  nnd2s1 U11293 ( .DIN1(n10808), .DIN2(n11097), .Q(n11090) );
  nnd2s1 U11294 ( .DIN1(n11098), .DIN2(n10510), .Q(n11097) );
  nor2s1 U11295 ( .DIN1(n11099), .DIN2(n11100), .Q(n11082) );
  and2s1 U11296 ( .DIN1(n10490), .DIN2(n11101), .Q(n11081) );
  nnd3s1 U11297 ( .DIN1(n11102), .DIN2(n10645), .DIN3(n10642), .Q(n11101) );
  nor3s1 U11298 ( .DIN1(n11103), .DIN2(n11104), .DIN3(n11105), .Q(n10802) );
  nnd4s1 U11299 ( .DIN1(n11106), .DIN2(n11107), .DIN3(n10625), .DIN4(n11108), 
        .Q(n11105) );
  and3s1 U11300 ( .DIN1(n11109), .DIN2(n11110), .DIN3(n11111), .Q(n11108) );
  nnd2s1 U11301 ( .DIN1(n10808), .DIN2(n10820), .Q(n11111) );
  nnd2s1 U11302 ( .DIN1(n11112), .DIN2(n10491), .Q(n11110) );
  nnd2s1 U11303 ( .DIN1(n11113), .DIN2(n10502), .Q(n11109) );
  nor2s1 U11304 ( .DIN1(n11114), .DIN2(n11115), .Q(n10625) );
  nnd4s1 U11305 ( .DIN1(n11116), .DIN2(n11117), .DIN3(n11118), .DIN4(n11119), 
        .Q(n11115) );
  nnd2s1 U11306 ( .DIN1(n10639), .DIN2(n11120), .Q(n11119) );
  nnd2s1 U11307 ( .DIN1(n10515), .DIN2(n11121), .Q(n11118) );
  nnd2s1 U11308 ( .DIN1(n10497), .DIN2(n11122), .Q(n11117) );
  nnd2s1 U11309 ( .DIN1(n10511), .DIN2(n10628), .Q(n11116) );
  nnd4s1 U11310 ( .DIN1(n11123), .DIN2(n11124), .DIN3(n11125), .DIN4(n11126), 
        .Q(n11114) );
  nnd2s1 U11311 ( .DIN1(n10627), .DIN2(n11121), .Q(n11126) );
  nnd2s1 U11312 ( .DIN1(n10501), .DIN2(n11127), .Q(n11125) );
  nnd2s1 U11313 ( .DIN1(n10646), .DIN2(n10829), .Q(n11127) );
  nnd2s1 U11314 ( .DIN1(n10489), .DIN2(n11128), .Q(n11124) );
  nnd2s1 U11315 ( .DIN1(n11129), .DIN2(n11130), .Q(n11128) );
  nnd2s1 U11316 ( .DIN1(n11112), .DIN2(n11131), .Q(n11123) );
  nnd3s1 U11317 ( .DIN1(n11132), .DIN2(n11133), .DIN3(n10518), .Q(n11131) );
  nnd3s1 U11318 ( .DIN1(n11134), .DIN2(n11135), .DIN3(n10493), .Q(n11104) );
  nnd2s1 U11319 ( .DIN1(n10827), .DIN2(n10819), .Q(n10493) );
  nnd2s1 U11320 ( .DIN1(n10489), .DIN2(n11136), .Q(n11135) );
  nnd3s1 U11321 ( .DIN1(n11137), .DIN2(n10832), .DIN3(n10634), .Q(n11136) );
  nor2s1 U11322 ( .DIN1(n10850), .DIN2(n10491), .Q(n10634) );
  nnd2s1 U11323 ( .DIN1(n10809), .DIN2(n10519), .Q(n11134) );
  nnd3s1 U11324 ( .DIN1(n11138), .DIN2(n11139), .DIN3(n11140), .Q(n11103) );
  nnd2s1 U11325 ( .DIN1(n10840), .DIN2(n11141), .Q(n11140) );
  nnd2s1 U11326 ( .DIN1(n10817), .DIN2(n10849), .Q(n11141) );
  nnd2s1 U11327 ( .DIN1(n10499), .DIN2(n11142), .Q(n11139) );
  nnd2s1 U11328 ( .DIN1(n10829), .DIN2(n10817), .Q(n11142) );
  nnd2s1 U11329 ( .DIN1(n10639), .DIN2(n11143), .Q(n11138) );
  nnd2s1 U11330 ( .DIN1(n11096), .DIN2(n10646), .Q(n11143) );
  nnd3s1 U11331 ( .DIN1(n11144), .DIN2(n11145), .DIN3(n11146), .Q(n11074) );
  nnd2s1 U11332 ( .DIN1(n10810), .DIN2(n11122), .Q(n11146) );
  nnd2s1 U11333 ( .DIN1(n10499), .DIN2(n10841), .Q(n11145) );
  nnd2s1 U11334 ( .DIN1(n10809), .DIN2(n10842), .Q(n11144) );
  nnd4s1 U11335 ( .DIN1(n11147), .DIN2(n11148), .DIN3(n11149), .DIN4(n11150), 
        .Q(n11073) );
  nnd2s1 U11336 ( .DIN1(n10497), .DIN2(n11151), .Q(n11150) );
  nnd2s1 U11337 ( .DIN1(n10826), .DIN2(n10642), .Q(n11151) );
  nnd2s1 U11338 ( .DIN1(n10627), .DIN2(n11152), .Q(n11149) );
  nnd2s1 U11339 ( .DIN1(n11133), .DIN2(n11129), .Q(n11152) );
  nnd2s1 U11340 ( .DIN1(n10643), .DIN2(n11153), .Q(n11148) );
  nnd2s1 U11341 ( .DIN1(n10507), .DIN2(n11154), .Q(n11147) );
  nnd2s1 U11342 ( .DIN1(n11155), .DIN2(n11130), .Q(n11154) );
  or3s1 U11343 ( .DIN1(n11156), .DIN2(n11157), .DIN3(n11158), .Q(n5698) );
  nnd4s1 U11344 ( .DIN1(n10858), .DIN2(n11159), .DIN3(n10658), .DIN4(n11160), 
        .Q(n11158) );
  and3s1 U11345 ( .DIN1(n11161), .DIN2(n11162), .DIN3(n11163), .Q(n11160) );
  nor4s1 U11346 ( .DIN1(n11164), .DIN2(n11165), .DIN3(n11166), .DIN4(n11167), 
        .Q(n10658) );
  nnd4s1 U11347 ( .DIN1(n11168), .DIN2(n11169), .DIN3(n11170), .DIN4(n11171), 
        .Q(n11167) );
  nnd2s1 U11348 ( .DIN1(n10661), .DIN2(n11172), .Q(n11171) );
  nnd2s1 U11349 ( .DIN1(n10866), .DIN2(n11173), .Q(n11169) );
  nnd2s1 U11350 ( .DIN1(n10887), .DIN2(n11174), .Q(n11168) );
  nnd3s1 U11351 ( .DIN1(n11175), .DIN2(n11176), .DIN3(n11177), .Q(n11166) );
  nnd2s1 U11352 ( .DIN1(n10901), .DIN2(n11178), .Q(n11177) );
  nnd2s1 U11353 ( .DIN1(n11179), .DIN2(n11180), .Q(n11178) );
  nnd2s1 U11354 ( .DIN1(n10893), .DIN2(n11181), .Q(n11176) );
  nnd2s1 U11355 ( .DIN1(n11182), .DIN2(n10912), .Q(n11181) );
  nnd2s1 U11356 ( .DIN1(n10877), .DIN2(n11183), .Q(n11175) );
  nnd2s1 U11357 ( .DIN1(n11184), .DIN2(n10917), .Q(n11183) );
  nor2s1 U11358 ( .DIN1(n11185), .DIN2(n11186), .Q(n11165) );
  and2s1 U11359 ( .DIN1(n10663), .DIN2(n11187), .Q(n11164) );
  nnd3s1 U11360 ( .DIN1(n11188), .DIN2(n10683), .DIN3(n10680), .Q(n11187) );
  nor3s1 U11361 ( .DIN1(n11189), .DIN2(n11190), .DIN3(n11191), .Q(n10858) );
  nnd4s1 U11362 ( .DIN1(n11192), .DIN2(n11193), .DIN3(n10659), .DIN4(n11194), 
        .Q(n11191) );
  and3s1 U11363 ( .DIN1(n11195), .DIN2(n11196), .DIN3(n11197), .Q(n11194) );
  nnd2s1 U11364 ( .DIN1(n10877), .DIN2(n10879), .Q(n11197) );
  nnd2s1 U11365 ( .DIN1(n11198), .DIN2(n10685), .Q(n11196) );
  nnd2s1 U11366 ( .DIN1(n11199), .DIN2(n10878), .Q(n11195) );
  nor2s1 U11367 ( .DIN1(n11200), .DIN2(n11201), .Q(n10659) );
  nnd4s1 U11368 ( .DIN1(n11202), .DIN2(n11203), .DIN3(n11204), .DIN4(n11205), 
        .Q(n11201) );
  nnd2s1 U11369 ( .DIN1(n10677), .DIN2(n11206), .Q(n11205) );
  nnd2s1 U11370 ( .DIN1(n10672), .DIN2(n11207), .Q(n11204) );
  nnd2s1 U11371 ( .DIN1(n11172), .DIN2(n11208), .Q(n11203) );
  nnd2s1 U11372 ( .DIN1(n10893), .DIN2(n10664), .Q(n11202) );
  nnd4s1 U11373 ( .DIN1(n11209), .DIN2(n11210), .DIN3(n11211), .DIN4(n11212), 
        .Q(n11200) );
  nnd2s1 U11374 ( .DIN1(n10661), .DIN2(n11207), .Q(n11212) );
  nnd2s1 U11375 ( .DIN1(n10884), .DIN2(n11213), .Q(n11211) );
  nnd2s1 U11376 ( .DIN1(n10684), .DIN2(n10889), .Q(n11213) );
  nnd2s1 U11377 ( .DIN1(n10904), .DIN2(n11214), .Q(n11210) );
  nnd2s1 U11378 ( .DIN1(n11215), .DIN2(n11216), .Q(n11214) );
  nnd2s1 U11379 ( .DIN1(n11198), .DIN2(n11217), .Q(n11209) );
  nnd3s1 U11380 ( .DIN1(n11218), .DIN2(n11219), .DIN3(n11220), .Q(n11217) );
  nnd3s1 U11381 ( .DIN1(n11221), .DIN2(n11222), .DIN3(n11223), .Q(n11190) );
  nnd2s1 U11382 ( .DIN1(n10904), .DIN2(n11224), .Q(n11222) );
  nnd3s1 U11383 ( .DIN1(n11225), .DIN2(n10892), .DIN3(n10671), .Q(n11224) );
  nor2s1 U11384 ( .DIN1(n10913), .DIN2(n10685), .Q(n10671) );
  nnd2s1 U11385 ( .DIN1(n10865), .DIN2(n10910), .Q(n11221) );
  nnd3s1 U11386 ( .DIN1(n11226), .DIN2(n11227), .DIN3(n11228), .Q(n11189) );
  nnd2s1 U11387 ( .DIN1(n10901), .DIN2(n11229), .Q(n11228) );
  nnd2s1 U11388 ( .DIN1(n10874), .DIN2(n10912), .Q(n11229) );
  nnd2s1 U11389 ( .DIN1(n10662), .DIN2(n11230), .Q(n11227) );
  nnd2s1 U11390 ( .DIN1(n10889), .DIN2(n10874), .Q(n11230) );
  nnd2s1 U11391 ( .DIN1(n10677), .DIN2(n11231), .Q(n11226) );
  nnd2s1 U11392 ( .DIN1(n11182), .DIN2(n10684), .Q(n11231) );
  nnd3s1 U11393 ( .DIN1(n11232), .DIN2(n11233), .DIN3(n11234), .Q(n11157) );
  nnd2s1 U11394 ( .DIN1(n10866), .DIN2(n11208), .Q(n11234) );
  nnd2s1 U11395 ( .DIN1(n10662), .DIN2(n10902), .Q(n11233) );
  nnd2s1 U11396 ( .DIN1(n10865), .DIN2(n10903), .Q(n11232) );
  nnd4s1 U11397 ( .DIN1(n11235), .DIN2(n11236), .DIN3(n11237), .DIN4(n11238), 
        .Q(n11156) );
  nnd2s1 U11398 ( .DIN1(n11172), .DIN2(n11239), .Q(n11238) );
  nnd2s1 U11399 ( .DIN1(n10886), .DIN2(n10680), .Q(n11239) );
  nnd2s1 U11400 ( .DIN1(n10661), .DIN2(n11240), .Q(n11237) );
  nnd2s1 U11401 ( .DIN1(n11219), .DIN2(n11215), .Q(n11240) );
  nnd2s1 U11402 ( .DIN1(n10681), .DIN2(n11241), .Q(n11236) );
  nnd2s1 U11403 ( .DIN1(n11242), .DIN2(n11243), .Q(n11235) );
  nnd2s1 U11404 ( .DIN1(n11244), .DIN2(n11216), .Q(n11243) );
  xor2s1 U11405 ( .DIN1(n10420), .DIN2(n11245), .Q(n11069) );
  xor2s1 U11406 ( .DIN1(n1496), .DIN2(n5025), .Q(n11245) );
  or3s1 U11407 ( .DIN1(n11246), .DIN2(n11247), .DIN3(n11248), .Q(n5025) );
  nnd4s1 U11408 ( .DIN1(n11249), .DIN2(n11250), .DIN3(n10527), .DIN4(n11251), 
        .Q(n11248) );
  and3s1 U11409 ( .DIN1(n10695), .DIN2(n10970), .DIN3(n10942), .Q(n11251) );
  nor4s1 U11410 ( .DIN1(n11252), .DIN2(n11253), .DIN3(n11254), .DIN4(n11255), 
        .Q(n10942) );
  nnd4s1 U11411 ( .DIN1(n11256), .DIN2(n11257), .DIN3(n11258), .DIN4(n11259), 
        .Q(n11255) );
  nor2s1 U11412 ( .DIN1(n11260), .DIN2(n11261), .Q(n11259) );
  nor2s1 U11413 ( .DIN1(n10964), .DIN2(n10754), .Q(n11261) );
  nor2s1 U11414 ( .DIN1(n10740), .DIN2(n10933), .Q(n11260) );
  or2s1 U11415 ( .DIN1(n10957), .DIN2(n11262), .Q(n11258) );
  nnd2s1 U11416 ( .DIN1(n10996), .DIN2(n11263), .Q(n11257) );
  nnd3s1 U11417 ( .DIN1(n10958), .DIN2(n10539), .DIN3(n10549), .Q(n11263) );
  nnd2s1 U11418 ( .DIN1(n11264), .DIN2(n11265), .Q(n11256) );
  nnd3s1 U11419 ( .DIN1(n11266), .DIN2(n10724), .DIN3(n10739), .Q(n11265) );
  nnd3s1 U11420 ( .DIN1(n11267), .DIN2(n11268), .DIN3(n11269), .Q(n11254) );
  nnd2s1 U11421 ( .DIN1(n10744), .DIN2(n10701), .Q(n11269) );
  nnd2s1 U11422 ( .DIN1(n10758), .DIN2(n10715), .Q(n11268) );
  nnd2s1 U11423 ( .DIN1(n10934), .DIN2(n10722), .Q(n11267) );
  nor2s1 U11424 ( .DIN1(n11270), .DIN2(n10537), .Q(n11253) );
  nor2s1 U11425 ( .DIN1(n10932), .DIN2(n11271), .Q(n11252) );
  nor4s1 U11426 ( .DIN1(n11272), .DIN2(n11273), .DIN3(n11274), .DIN4(n11275), 
        .Q(n10970) );
  nnd4s1 U11427 ( .DIN1(n11276), .DIN2(n11277), .DIN3(n11278), .DIN4(n11279), 
        .Q(n11275) );
  nnd2s1 U11428 ( .DIN1(n10716), .DIN2(n10952), .Q(n11279) );
  nor2s1 U11429 ( .DIN1(n11280), .DIN2(n11281), .Q(n11278) );
  nor2s1 U11430 ( .DIN1(n11266), .DIN2(n10957), .Q(n11281) );
  nor2s1 U11431 ( .DIN1(n10734), .DIN2(n10964), .Q(n11280) );
  nnd2s1 U11432 ( .DIN1(n10752), .DIN2(n10722), .Q(n11277) );
  nnd2s1 U11433 ( .DIN1(n10533), .DIN2(n10702), .Q(n11276) );
  nnd3s1 U11434 ( .DIN1(n11282), .DIN2(n11283), .DIN3(n11284), .Q(n11274) );
  nnd2s1 U11435 ( .DIN1(n10532), .DIN2(n11285), .Q(n11284) );
  nnd2s1 U11436 ( .DIN1(n10939), .DIN2(n10724), .Q(n11285) );
  nnd2s1 U11437 ( .DIN1(n10701), .DIN2(n11286), .Q(n11283) );
  nnd2s1 U11438 ( .DIN1(n11287), .DIN2(n10958), .Q(n11286) );
  nnd2s1 U11439 ( .DIN1(n10744), .DIN2(n11288), .Q(n11282) );
  nnd2s1 U11440 ( .DIN1(n10998), .DIN2(n10757), .Q(n11288) );
  nor2s1 U11441 ( .DIN1(n11289), .DIN2(n10756), .Q(n11273) );
  nor2s1 U11442 ( .DIN1(n10951), .DIN2(n10937), .Q(n11289) );
  nor2s1 U11443 ( .DIN1(n11290), .DIN2(n10548), .Q(n11272) );
  nor2s1 U11444 ( .DIN1(n10996), .DIN2(n10749), .Q(n11290) );
  nor4s1 U11445 ( .DIN1(n11291), .DIN2(n11292), .DIN3(n11293), .DIN4(n11294), 
        .Q(n10695) );
  nnd4s1 U11446 ( .DIN1(n11295), .DIN2(n11296), .DIN3(n11297), .DIN4(n11298), 
        .Q(n11294) );
  nor2s1 U11447 ( .DIN1(n11299), .DIN2(n11300), .Q(n11297) );
  nor2s1 U11448 ( .DIN1(n10940), .DIN2(n10558), .Q(n11300) );
  nor2s1 U11449 ( .DIN1(n10712), .DIN2(n10964), .Q(n11299) );
  nnd2s1 U11450 ( .DIN1(n10934), .DIN2(n10952), .Q(n11296) );
  nnd2s1 U11451 ( .DIN1(n10703), .DIN2(n10729), .Q(n11295) );
  nnd3s1 U11452 ( .DIN1(n11301), .DIN2(n11302), .DIN3(n11303), .Q(n11293) );
  nnd2s1 U11453 ( .DIN1(n10533), .DIN2(n11304), .Q(n11303) );
  nnd2s1 U11454 ( .DIN1(n10541), .DIN2(n11305), .Q(n11302) );
  nnd2s1 U11455 ( .DIN1(n10724), .DIN2(n10940), .Q(n11305) );
  nnd2s1 U11456 ( .DIN1(n10996), .DIN2(n11306), .Q(n11301) );
  nnd3s1 U11457 ( .DIN1(n10966), .DIN2(n10957), .DIN3(n11307), .Q(n11306) );
  nor2s1 U11458 ( .DIN1(n10725), .DIN2(n10557), .Q(n11292) );
  nor2s1 U11459 ( .DIN1(n10552), .DIN2(n10756), .Q(n11291) );
  nor3s1 U11460 ( .DIN1(n11308), .DIN2(n11309), .DIN3(n11310), .Q(n10527) );
  nnd4s1 U11461 ( .DIN1(n10971), .DIN2(n10697), .DIN3(n11008), .DIN4(n11311), 
        .Q(n11310) );
  and3s1 U11462 ( .DIN1(n11312), .DIN2(n11313), .DIN3(n11314), .Q(n11311) );
  nnd2s1 U11463 ( .DIN1(n10533), .DIN2(n10937), .Q(n11314) );
  nnd2s1 U11464 ( .DIN1(n10714), .DIN2(n10952), .Q(n11313) );
  nnd2s1 U11465 ( .DIN1(n10742), .DIN2(n10555), .Q(n11312) );
  nor4s1 U11466 ( .DIN1(n11315), .DIN2(n11316), .DIN3(n11317), .DIN4(n11318), 
        .Q(n11008) );
  nnd4s1 U11467 ( .DIN1(n11319), .DIN2(n11320), .DIN3(n11321), .DIN4(n11322), 
        .Q(n11318) );
  nnd2s1 U11468 ( .DIN1(n10555), .DIN2(n11323), .Q(n11322) );
  nor2s1 U11469 ( .DIN1(n11324), .DIN2(n11325), .Q(n11321) );
  nor2s1 U11470 ( .DIN1(n11326), .DIN2(n10966), .Q(n11325) );
  nor2s1 U11471 ( .DIN1(n10714), .DIN2(n10934), .Q(n11326) );
  nor2s1 U11472 ( .DIN1(n11327), .DIN2(n10757), .Q(n11324) );
  nor2s1 U11473 ( .DIN1(n10742), .DIN2(n10554), .Q(n11327) );
  nnd2s1 U11474 ( .DIN1(n10937), .DIN2(n11328), .Q(n11320) );
  nnd3s1 U11475 ( .DIN1(n10725), .DIN2(n10932), .DIN3(n10992), .Q(n11328) );
  nnd2s1 U11476 ( .DIN1(n10749), .DIN2(n11329), .Q(n11319) );
  nnd3s1 U11477 ( .DIN1(n11330), .DIN2(n11331), .DIN3(n11332), .Q(n11317) );
  nnd2s1 U11478 ( .DIN1(n10996), .DIN2(n10951), .Q(n11332) );
  nnd2s1 U11479 ( .DIN1(n10744), .DIN2(n10758), .Q(n11330) );
  nor2s1 U11480 ( .DIN1(n10939), .DIN2(n10957), .Q(n11316) );
  nor2s1 U11481 ( .DIN1(n10756), .DIN2(n10754), .Q(n11315) );
  nor4s1 U11482 ( .DIN1(n11333), .DIN2(n11334), .DIN3(n11335), .DIN4(n11336), 
        .Q(n10697) );
  nnd4s1 U11483 ( .DIN1(n11337), .DIN2(n11338), .DIN3(n11339), .DIN4(n11340), 
        .Q(n11336) );
  nnd2s1 U11484 ( .DIN1(n10937), .DIN2(n10758), .Q(n11340) );
  nnd2s1 U11485 ( .DIN1(n10749), .DIN2(n11264), .Q(n11339) );
  nnd2s1 U11486 ( .DIN1(n10752), .DIN2(n10952), .Q(n11338) );
  nnd2s1 U11487 ( .DIN1(n10555), .DIN2(n10715), .Q(n11337) );
  nnd3s1 U11488 ( .DIN1(n11341), .DIN2(n11342), .DIN3(n11343), .Q(n11335) );
  nnd2s1 U11489 ( .DIN1(n10550), .DIN2(n11344), .Q(n11343) );
  nnd2s1 U11490 ( .DIN1(n11003), .DIN2(n10731), .Q(n11344) );
  nor2s1 U11491 ( .DIN1(n10744), .DIN2(n10951), .Q(n11003) );
  nnd2s1 U11492 ( .DIN1(n10743), .DIN2(n11345), .Q(n11342) );
  nnd2s1 U11493 ( .DIN1(n11287), .DIN2(n10731), .Q(n11345) );
  nor2s1 U11494 ( .DIN1(n10951), .DIN2(n11329), .Q(n11287) );
  nnd2s1 U11495 ( .DIN1(n10990), .DIN2(n11346), .Q(n11341) );
  nnd2s1 U11496 ( .DIN1(n10939), .DIN2(n10964), .Q(n11346) );
  nor2s1 U11497 ( .DIN1(n10964), .DIN2(n10957), .Q(n11334) );
  nor2s1 U11498 ( .DIN1(n10713), .DIN2(n10940), .Q(n11333) );
  hi1s1 U11499 ( .DIN(n11347), .Q(n10713) );
  nor2s1 U11500 ( .DIN1(n11348), .DIN2(n11349), .Q(n10971) );
  nnd4s1 U11501 ( .DIN1(n11350), .DIN2(n11351), .DIN3(n11352), .DIN4(n11353), 
        .Q(n11349) );
  nnd2s1 U11502 ( .DIN1(n10952), .DIN2(n11354), .Q(n11353) );
  nnd3s1 U11503 ( .DIN1(n11266), .DIN2(n10940), .DIN3(n10725), .Q(n11354) );
  nnd2s1 U11504 ( .DIN1(n10934), .DIN2(n10702), .Q(n11350) );
  nnd4s1 U11505 ( .DIN1(n11355), .DIN2(n11356), .DIN3(n11357), .DIN4(n11358), 
        .Q(n11348) );
  nnd2s1 U11506 ( .DIN1(n10716), .DIN2(n11359), .Q(n11358) );
  nnd2s1 U11507 ( .DIN1(n10990), .DIN2(n11360), .Q(n11357) );
  nnd2s1 U11508 ( .DIN1(n10538), .DIN2(n10932), .Q(n11360) );
  nnd2s1 U11509 ( .DIN1(n10752), .DIN2(n11361), .Q(n11356) );
  nnd2s1 U11510 ( .DIN1(n11362), .DIN2(n10557), .Q(n11361) );
  nnd2s1 U11511 ( .DIN1(n10541), .DIN2(n11363), .Q(n11355) );
  nnd2s1 U11512 ( .DIN1(n10933), .DIN2(n10725), .Q(n11363) );
  nnd3s1 U11513 ( .DIN1(n11364), .DIN2(n11365), .DIN3(n11366), .Q(n11309) );
  nnd2s1 U11514 ( .DIN1(n10710), .DIN2(n11329), .Q(n11366) );
  nnd2s1 U11515 ( .DIN1(n10951), .DIN2(n11367), .Q(n11365) );
  nnd3s1 U11516 ( .DIN1(n10992), .DIN2(n11266), .DIN3(n11368), .Q(n11367) );
  or2s1 U11517 ( .DIN1(n10731), .DIN2(n11369), .Q(n11364) );
  nnd3s1 U11518 ( .DIN1(n11370), .DIN2(n11371), .DIN3(n11372), .Q(n11308) );
  nnd2s1 U11519 ( .DIN1(n10541), .DIN2(n11373), .Q(n11372) );
  nnd2s1 U11520 ( .DIN1(n10739), .DIN2(n10998), .Q(n11373) );
  nnd2s1 U11521 ( .DIN1(n10749), .DIN2(n11374), .Q(n11371) );
  nnd2s1 U11522 ( .DIN1(n10961), .DIN2(n10958), .Q(n11374) );
  nnd2s1 U11523 ( .DIN1(n10729), .DIN2(n11375), .Q(n11370) );
  nnd2s1 U11524 ( .DIN1(n10740), .DIN2(n10966), .Q(n11375) );
  nor2s1 U11525 ( .DIN1(n10717), .DIN2(n10744), .Q(n10740) );
  nnd2s1 U11526 ( .DIN1(n10703), .DIN2(n10710), .Q(n11250) );
  nnd3s1 U11527 ( .DIN1(n11376), .DIN2(n11377), .DIN3(n11378), .Q(n11247) );
  nnd2s1 U11528 ( .DIN1(n10555), .DIN2(n10722), .Q(n11378) );
  nnd2s1 U11529 ( .DIN1(n11379), .DIN2(n11380), .Q(n11377) );
  nnd2s1 U11530 ( .DIN1(n11329), .DIN2(n10752), .Q(n11376) );
  nnd4s1 U11531 ( .DIN1(n11381), .DIN2(n11382), .DIN3(n11383), .DIN4(n11384), 
        .Q(n11246) );
  nnd2s1 U11532 ( .DIN1(n10743), .DIN2(n11385), .Q(n11384) );
  nnd2s1 U11533 ( .DIN1(n10552), .DIN2(n10754), .Q(n11385) );
  nor2s1 U11534 ( .DIN1(n10715), .DIN2(n10702), .Q(n10552) );
  nnd2s1 U11535 ( .DIN1(n10744), .DIN2(n11386), .Q(n11383) );
  nnd2s1 U11536 ( .DIN1(n10992), .DIN2(n10728), .Q(n11386) );
  nnd2s1 U11537 ( .DIN1(n10715), .DIN2(n11387), .Q(n11382) );
  nnd2s1 U11538 ( .DIN1(n10727), .DIN2(n10739), .Q(n11387) );
  nnd2s1 U11539 ( .DIN1(n10937), .DIN2(n10983), .Q(n11381) );
  or3s1 U11540 ( .DIN1(n11388), .DIN2(n11389), .DIN3(n11390), .Q(n10420) );
  nnd4s1 U11541 ( .DIN1(n11012), .DIN2(n11391), .DIN3(n10767), .DIN4(n11392), 
        .Q(n11390) );
  and3s1 U11542 ( .DIN1(n11393), .DIN2(n11394), .DIN3(n11395), .Q(n11392) );
  nor4s1 U11543 ( .DIN1(n11396), .DIN2(n11397), .DIN3(n11398), .DIN4(n11399), 
        .Q(n10767) );
  nnd4s1 U11544 ( .DIN1(n11400), .DIN2(n11401), .DIN3(n11402), .DIN4(n11403), 
        .Q(n11399) );
  nnd2s1 U11545 ( .DIN1(n10770), .DIN2(n10578), .Q(n11403) );
  nnd2s1 U11546 ( .DIN1(n11020), .DIN2(n11404), .Q(n11401) );
  nnd2s1 U11547 ( .DIN1(n11037), .DIN2(n10579), .Q(n11400) );
  nnd3s1 U11548 ( .DIN1(n11405), .DIN2(n11406), .DIN3(n11407), .Q(n11398) );
  nnd2s1 U11549 ( .DIN1(n11050), .DIN2(n11408), .Q(n11407) );
  nnd2s1 U11550 ( .DIN1(n11409), .DIN2(n10594), .Q(n11408) );
  nnd2s1 U11551 ( .DIN1(n10592), .DIN2(n11410), .Q(n11406) );
  nnd2s1 U11552 ( .DIN1(n11411), .DIN2(n11059), .Q(n11410) );
  nnd2s1 U11553 ( .DIN1(n11018), .DIN2(n11412), .Q(n11405) );
  nnd2s1 U11554 ( .DIN1(n11413), .DIN2(n10591), .Q(n11412) );
  nor2s1 U11555 ( .DIN1(n11414), .DIN2(n11415), .Q(n11397) );
  and2s1 U11556 ( .DIN1(n10571), .DIN2(n11416), .Q(n11396) );
  nnd3s1 U11557 ( .DIN1(n11417), .DIN2(n10788), .DIN3(n10785), .Q(n11416) );
  nor3s1 U11558 ( .DIN1(n11418), .DIN2(n11419), .DIN3(n11420), .Q(n11012) );
  nnd4s1 U11559 ( .DIN1(n11421), .DIN2(n11422), .DIN3(n10768), .DIN4(n11423), 
        .Q(n11420) );
  and3s1 U11560 ( .DIN1(n11424), .DIN2(n11425), .DIN3(n11426), .Q(n11423) );
  nnd2s1 U11561 ( .DIN1(n11018), .DIN2(n11030), .Q(n11426) );
  nnd2s1 U11562 ( .DIN1(n11427), .DIN2(n10572), .Q(n11425) );
  nnd2s1 U11563 ( .DIN1(n11428), .DIN2(n10583), .Q(n11424) );
  nor2s1 U11564 ( .DIN1(n11429), .DIN2(n11430), .Q(n10768) );
  nnd4s1 U11565 ( .DIN1(n11431), .DIN2(n11432), .DIN3(n11433), .DIN4(n11434), 
        .Q(n11430) );
  nnd2s1 U11566 ( .DIN1(n10782), .DIN2(n11435), .Q(n11434) );
  nnd2s1 U11567 ( .DIN1(n10596), .DIN2(n11436), .Q(n11433) );
  nnd2s1 U11568 ( .DIN1(n10578), .DIN2(n11437), .Q(n11432) );
  nnd2s1 U11569 ( .DIN1(n10592), .DIN2(n10771), .Q(n11431) );
  nnd4s1 U11570 ( .DIN1(n11438), .DIN2(n11439), .DIN3(n11440), .DIN4(n11441), 
        .Q(n11429) );
  nnd2s1 U11571 ( .DIN1(n10770), .DIN2(n11436), .Q(n11441) );
  nnd2s1 U11572 ( .DIN1(n10582), .DIN2(n11442), .Q(n11440) );
  nnd2s1 U11573 ( .DIN1(n10789), .DIN2(n11039), .Q(n11442) );
  nnd2s1 U11574 ( .DIN1(n10570), .DIN2(n11443), .Q(n11439) );
  nnd2s1 U11575 ( .DIN1(n11444), .DIN2(n11445), .Q(n11443) );
  nnd2s1 U11576 ( .DIN1(n11427), .DIN2(n11446), .Q(n11438) );
  nnd3s1 U11577 ( .DIN1(n11447), .DIN2(n11448), .DIN3(n10599), .Q(n11446) );
  nnd3s1 U11578 ( .DIN1(n11449), .DIN2(n11450), .DIN3(n10574), .Q(n11419) );
  nnd2s1 U11579 ( .DIN1(n11037), .DIN2(n11029), .Q(n10574) );
  nnd2s1 U11580 ( .DIN1(n10570), .DIN2(n11451), .Q(n11450) );
  nnd3s1 U11581 ( .DIN1(n11452), .DIN2(n11042), .DIN3(n10777), .Q(n11451) );
  nor2s1 U11582 ( .DIN1(n11060), .DIN2(n10572), .Q(n10777) );
  nnd2s1 U11583 ( .DIN1(n11019), .DIN2(n10600), .Q(n11449) );
  nnd3s1 U11584 ( .DIN1(n11453), .DIN2(n11454), .DIN3(n11455), .Q(n11418) );
  nnd2s1 U11585 ( .DIN1(n11050), .DIN2(n11456), .Q(n11455) );
  nnd2s1 U11586 ( .DIN1(n11027), .DIN2(n11059), .Q(n11456) );
  nnd2s1 U11587 ( .DIN1(n10580), .DIN2(n11457), .Q(n11454) );
  nnd2s1 U11588 ( .DIN1(n11039), .DIN2(n11027), .Q(n11457) );
  nnd2s1 U11589 ( .DIN1(n10782), .DIN2(n11458), .Q(n11453) );
  nnd2s1 U11590 ( .DIN1(n11411), .DIN2(n10789), .Q(n11458) );
  nnd3s1 U11591 ( .DIN1(n11459), .DIN2(n11460), .DIN3(n11461), .Q(n11389) );
  nnd2s1 U11592 ( .DIN1(n11020), .DIN2(n11437), .Q(n11461) );
  nnd2s1 U11593 ( .DIN1(n10580), .DIN2(n11051), .Q(n11460) );
  nnd2s1 U11594 ( .DIN1(n11019), .DIN2(n11052), .Q(n11459) );
  nnd4s1 U11595 ( .DIN1(n11462), .DIN2(n11463), .DIN3(n11464), .DIN4(n11465), 
        .Q(n11388) );
  nnd2s1 U11596 ( .DIN1(n10578), .DIN2(n11466), .Q(n11465) );
  nnd2s1 U11597 ( .DIN1(n11036), .DIN2(n10785), .Q(n11466) );
  nnd2s1 U11598 ( .DIN1(n10770), .DIN2(n11467), .Q(n11464) );
  nnd2s1 U11599 ( .DIN1(n11448), .DIN2(n11444), .Q(n11467) );
  nnd2s1 U11600 ( .DIN1(n10786), .DIN2(n11468), .Q(n11463) );
  nnd2s1 U11601 ( .DIN1(n10588), .DIN2(n11469), .Q(n11462) );
  nnd2s1 U11602 ( .DIN1(n11470), .DIN2(n11445), .Q(n11469) );
  nnd2s1 U11603 ( .DIN1(n11471), .DIN2(n1600), .Q(n11066) );
  xor2s1 U11604 ( .DIN1(w1[4]), .DIN2(text_in_r[68]), .Q(n11471) );
  nnd2s1 U11605 ( .DIN1(n11472), .DIN2(n11473), .Q(N165) );
  nnd2s1 U11606 ( .DIN1(n11474), .DIN2(n1632), .Q(n11473) );
  xor2s1 U11607 ( .DIN1(n11475), .DIN2(n11476), .Q(n11474) );
  xor2s1 U11608 ( .DIN1(n11477), .DIN2(n11478), .Q(n11476) );
  xor2s1 U11609 ( .DIN1(n5424), .DIN2(n10442), .Q(n11478) );
  xnr2s1 U11610 ( .DIN1(n5425), .DIN2(n11479), .Q(n10442) );
  hi1s1 U11611 ( .DIN(n5072), .Q(n11479) );
  or3s1 U11612 ( .DIN1(n11480), .DIN2(n11481), .DIN3(n11482), .Q(n5072) );
  nnd4s1 U11613 ( .DIN1(n11483), .DIN2(n11484), .DIN3(n10622), .DIN4(n11485), 
        .Q(n11482) );
  and3s1 U11614 ( .DIN1(n10803), .DIN2(n11106), .DIN3(n11076), .Q(n11485) );
  nor4s1 U11615 ( .DIN1(n11486), .DIN2(n11487), .DIN3(n11488), .DIN4(n11489), 
        .Q(n11076) );
  nnd4s1 U11616 ( .DIN1(n11490), .DIN2(n11491), .DIN3(n11492), .DIN4(n11493), 
        .Q(n11489) );
  nnd2s1 U11617 ( .DIN1(n10502), .DIN2(n10643), .Q(n11493) );
  nor2s1 U11618 ( .DIN1(n11494), .DIN2(n11495), .Q(n11492) );
  nor2s1 U11619 ( .DIN1(n10642), .DIN2(n11496), .Q(n11495) );
  nor2s1 U11620 ( .DIN1(n11497), .DIN2(n10849), .Q(n11494) );
  nnd2s1 U11621 ( .DIN1(n10492), .DIN2(n10820), .Q(n11491) );
  nnd2s1 U11622 ( .DIN1(n10827), .DIN2(n10515), .Q(n11490) );
  nnd3s1 U11623 ( .DIN1(n11498), .DIN2(n11499), .DIN3(n11500), .Q(n11488) );
  nnd2s1 U11624 ( .DIN1(n10850), .DIN2(n10854), .Q(n11500) );
  nnd2s1 U11625 ( .DIN1(n10500), .DIN2(n11501), .Q(n11499) );
  nnd3s1 U11626 ( .DIN1(n11098), .DIN2(n11496), .DIN3(n11132), .Q(n11501) );
  nnd2s1 U11627 ( .DIN1(n11113), .DIN2(n11502), .Q(n11498) );
  nnd3s1 U11628 ( .DIN1(n10817), .DIN2(n10514), .DIN3(n10641), .Q(n11502) );
  nor2s1 U11629 ( .DIN1(n10817), .DIN2(n10518), .Q(n11487) );
  nor2s1 U11630 ( .DIN1(n11503), .DIN2(n11504), .Q(n11486) );
  nor4s1 U11631 ( .DIN1(n11505), .DIN2(n11506), .DIN3(n11507), .DIN4(n11508), 
        .Q(n11106) );
  nnd4s1 U11632 ( .DIN1(n11509), .DIN2(n11510), .DIN3(n11511), .DIN4(n11512), 
        .Q(n11508) );
  nor2s1 U11633 ( .DIN1(n11513), .DIN2(n11514), .Q(n11512) );
  nor2s1 U11634 ( .DIN1(n11496), .DIN2(n11504), .Q(n11514) );
  nor2s1 U11635 ( .DIN1(n10853), .DIN2(n10514), .Q(n11513) );
  nnd2s1 U11636 ( .DIN1(n10628), .DIN2(n10519), .Q(n11510) );
  nnd2s1 U11637 ( .DIN1(n10809), .DIN2(n10499), .Q(n11509) );
  nnd3s1 U11638 ( .DIN1(n11515), .DIN2(n11516), .DIN3(n11517), .Q(n11507) );
  nnd2s1 U11639 ( .DIN1(n10819), .DIN2(n11518), .Q(n11517) );
  nnd2s1 U11640 ( .DIN1(n11133), .DIN2(n10832), .Q(n11518) );
  nnd2s1 U11641 ( .DIN1(n10627), .DIN2(n11519), .Q(n11516) );
  nnd2s1 U11642 ( .DIN1(n11155), .DIN2(n11098), .Q(n11519) );
  nnd2s1 U11643 ( .DIN1(n10501), .DIN2(n10851), .Q(n11515) );
  nnd2s1 U11644 ( .DIN1(n10834), .DIN2(n11099), .Q(n10851) );
  nor2s1 U11645 ( .DIN1(n11520), .DIN2(n10646), .Q(n11506) );
  nor2s1 U11646 ( .DIN1(n10490), .DIN2(n10511), .Q(n11520) );
  nor2s1 U11647 ( .DIN1(n11521), .DIN2(n11130), .Q(n11505) );
  and2s1 U11648 ( .DIN1(n10817), .DIN2(n11522), .Q(n11521) );
  nor4s1 U11649 ( .DIN1(n11523), .DIN2(n11524), .DIN3(n11525), .DIN4(n11526), 
        .Q(n10803) );
  nnd4s1 U11650 ( .DIN1(n11527), .DIN2(n11528), .DIN3(n11529), .DIN4(n11530), 
        .Q(n11526) );
  nnd2s1 U11651 ( .DIN1(n11112), .DIN2(n10820), .Q(n11530) );
  nor2s1 U11652 ( .DIN1(n11531), .DIN2(n11532), .Q(n11529) );
  nor2s1 U11653 ( .DIN1(n11533), .DIN2(n10646), .Q(n11531) );
  nnd2s1 U11654 ( .DIN1(n10808), .DIN2(n10827), .Q(n11528) );
  nnd2s1 U11655 ( .DIN1(n10810), .DIN2(n10507), .Q(n11527) );
  nnd3s1 U11656 ( .DIN1(n11534), .DIN2(n11535), .DIN3(n11536), .Q(n11525) );
  nnd2s1 U11657 ( .DIN1(n10499), .DIN2(n11537), .Q(n11536) );
  nnd2s1 U11658 ( .DIN1(n10515), .DIN2(n11538), .Q(n11535) );
  nnd2s1 U11659 ( .DIN1(n11130), .DIN2(n11098), .Q(n11538) );
  nnd2s1 U11660 ( .DIN1(n11113), .DIN2(n11539), .Q(n11534) );
  nnd3s1 U11661 ( .DIN1(n11102), .DIN2(n11504), .DIN3(n11540), .Q(n11539) );
  nor2s1 U11662 ( .DIN1(n10514), .DIN2(n10518), .Q(n11524) );
  nor2s1 U11663 ( .DIN1(n10648), .DIN2(n10510), .Q(n11523) );
  nor3s1 U11664 ( .DIN1(n11541), .DIN2(n11542), .DIN3(n11543), .Q(n10622) );
  nnd4s1 U11665 ( .DIN1(n11107), .DIN2(n10805), .DIN3(n11080), .DIN4(n11544), 
        .Q(n11543) );
  and3s1 U11666 ( .DIN1(n11545), .DIN2(n11546), .DIN3(n11547), .Q(n11544) );
  nnd2s1 U11667 ( .DIN1(n10810), .DIN2(n10498), .Q(n11547) );
  nnd2s1 U11668 ( .DIN1(n10489), .DIN2(n10643), .Q(n11545) );
  nor4s1 U11669 ( .DIN1(n11548), .DIN2(n11549), .DIN3(n11550), .DIN4(n11551), 
        .Q(n11080) );
  nnd4s1 U11670 ( .DIN1(n11552), .DIN2(n11553), .DIN3(n11554), .DIN4(n11555), 
        .Q(n11551) );
  nnd2s1 U11671 ( .DIN1(n10810), .DIN2(n11556), .Q(n11555) );
  nnd2s1 U11672 ( .DIN1(n11557), .DIN2(n11102), .Q(n11556) );
  nor2s1 U11673 ( .DIN1(n11558), .DIN2(n11559), .Q(n11554) );
  nor2s1 U11674 ( .DIN1(n11560), .DIN2(n10853), .Q(n11559) );
  nor2s1 U11675 ( .DIN1(n10489), .DIN2(n10650), .Q(n11560) );
  nor2s1 U11676 ( .DIN1(n11561), .DIN2(n10517), .Q(n11558) );
  nor2s1 U11677 ( .DIN1(n11562), .DIN2(n10809), .Q(n11561) );
  nnd2s1 U11678 ( .DIN1(n10507), .DIN2(n11563), .Q(n11553) );
  nnd3s1 U11679 ( .DIN1(n11533), .DIN2(n11129), .DIN3(n10518), .Q(n11563) );
  nnd2s1 U11680 ( .DIN1(n11113), .DIN2(n11562), .Q(n11552) );
  nnd3s1 U11681 ( .DIN1(n11564), .DIN2(n11565), .DIN3(n11566), .Q(n11550) );
  nnd2s1 U11682 ( .DIN1(n10850), .DIN2(n11567), .Q(n11566) );
  nnd2s1 U11683 ( .DIN1(n10497), .DIN2(n10500), .Q(n11565) );
  nnd2s1 U11684 ( .DIN1(n10627), .DIN2(n10501), .Q(n11564) );
  nor2s1 U11685 ( .DIN1(n11496), .DIN2(n10646), .Q(n11549) );
  nor2s1 U11686 ( .DIN1(n11155), .DIN2(n11504), .Q(n11548) );
  nor4s1 U11687 ( .DIN1(n11568), .DIN2(n11569), .DIN3(n11570), .DIN4(n11571), 
        .Q(n10805) );
  nnd4s1 U11688 ( .DIN1(n11572), .DIN2(n11573), .DIN3(n11574), .DIN4(n11575), 
        .Q(n11571) );
  nnd2s1 U11689 ( .DIN1(n10498), .DIN2(n10519), .Q(n11575) );
  nnd2s1 U11690 ( .DIN1(n10643), .DIN2(n10819), .Q(n11574) );
  nnd2s1 U11691 ( .DIN1(n10840), .DIN2(n10507), .Q(n11573) );
  nnd2s1 U11692 ( .DIN1(n10808), .DIN2(n10810), .Q(n11572) );
  nnd3s1 U11693 ( .DIN1(n11576), .DIN2(n11577), .DIN3(n11578), .Q(n11570) );
  nnd2s1 U11694 ( .DIN1(n10491), .DIN2(n11579), .Q(n11578) );
  nnd3s1 U11695 ( .DIN1(n10829), .DIN2(n11099), .DIN3(n10646), .Q(n11579) );
  nnd2s1 U11696 ( .DIN1(n10843), .DIN2(n11580), .Q(n11577) );
  nnd2s1 U11697 ( .DIN1(n11522), .DIN2(n10829), .Q(n11580) );
  nor2s1 U11698 ( .DIN1(n11567), .DIN2(n11562), .Q(n11522) );
  nnd2s1 U11699 ( .DIN1(n11112), .DIN2(n11581), .Q(n11576) );
  nnd2s1 U11700 ( .DIN1(n11497), .DIN2(n11155), .Q(n11581) );
  nor2s1 U11701 ( .DIN1(n11102), .DIN2(n11133), .Q(n11569) );
  nor2s1 U11702 ( .DIN1(n10835), .DIN2(n11130), .Q(n11568) );
  hi1s1 U11703 ( .DIN(n10520), .Q(n10835) );
  nor2s1 U11704 ( .DIN1(n11582), .DIN2(n11583), .Q(n11107) );
  nnd4s1 U11705 ( .DIN1(n11584), .DIN2(n11585), .DIN3(n11586), .DIN4(n11587), 
        .Q(n11583) );
  nnd2s1 U11706 ( .DIN1(n10498), .DIN2(n11588), .Q(n11587) );
  nnd3s1 U11707 ( .DIN1(n11130), .DIN2(n11496), .DIN3(n11533), .Q(n11588) );
  nnd2s1 U11708 ( .DIN1(n10497), .DIN2(n10809), .Q(n11585) );
  nnd4s1 U11709 ( .DIN1(n11589), .DIN2(n11590), .DIN3(n11591), .DIN4(n11592), 
        .Q(n11582) );
  nnd2s1 U11710 ( .DIN1(n10519), .DIN2(n11593), .Q(n11592) );
  nnd2s1 U11711 ( .DIN1(n11594), .DIN2(n10646), .Q(n11593) );
  nnd2s1 U11712 ( .DIN1(n10490), .DIN2(n11595), .Q(n11591) );
  nnd2s1 U11713 ( .DIN1(n10515), .DIN2(n11596), .Q(n11590) );
  nnd2s1 U11714 ( .DIN1(n11133), .DIN2(n11533), .Q(n11596) );
  nnd2s1 U11715 ( .DIN1(n11112), .DIN2(n11597), .Q(n11589) );
  nnd2s1 U11716 ( .DIN1(n10633), .DIN2(n11129), .Q(n11597) );
  nnd3s1 U11717 ( .DIN1(n11598), .DIN2(n11599), .DIN3(n11600), .Q(n11542) );
  nnd2s1 U11718 ( .DIN1(n10499), .DIN2(n10507), .Q(n11600) );
  nnd2s1 U11719 ( .DIN1(n11562), .DIN2(n11601), .Q(n11599) );
  nnd3s1 U11720 ( .DIN1(n10518), .DIN2(n11496), .DIN3(n11602), .Q(n11601) );
  or2s1 U11721 ( .DIN1(n10829), .DIN2(n11603), .Q(n11598) );
  nnd3s1 U11722 ( .DIN1(n11604), .DIN2(n11605), .DIN3(n11606), .Q(n11541) );
  nnd2s1 U11723 ( .DIN1(n10515), .DIN2(n11607), .Q(n11606) );
  nnd2s1 U11724 ( .DIN1(n11137), .DIN2(n11132), .Q(n11607) );
  nnd2s1 U11725 ( .DIN1(n10827), .DIN2(n11608), .Q(n11605) );
  or2s1 U11726 ( .DIN1(n10854), .DIN2(n10500), .Q(n11608) );
  nnd2s1 U11727 ( .DIN1(n10646), .DIN2(n10632), .Q(n10854) );
  nnd2s1 U11728 ( .DIN1(n10850), .DIN2(n11609), .Q(n11604) );
  nnd2s1 U11729 ( .DIN1(n10513), .DIN2(n10817), .Q(n11609) );
  nnd2s1 U11730 ( .DIN1(n10643), .DIN2(n10628), .Q(n11484) );
  nnd2s1 U11731 ( .DIN1(n10808), .DIN2(n10511), .Q(n11483) );
  nnd3s1 U11732 ( .DIN1(n11610), .DIN2(n11611), .DIN3(n11612), .Q(n11481) );
  nnd2s1 U11733 ( .DIN1(n11567), .DIN2(n10519), .Q(n11612) );
  nnd2s1 U11734 ( .DIN1(n11089), .DIN2(n11613), .Q(n11611) );
  nnd4s1 U11735 ( .DIN1(n11614), .DIN2(n11615), .DIN3(n11616), .DIN4(n11617), 
        .Q(n11480) );
  nnd2s1 U11736 ( .DIN1(n10843), .DIN2(n11618), .Q(n11617) );
  nnd2s1 U11737 ( .DIN1(n10648), .DIN2(n10849), .Q(n11618) );
  nor2s1 U11738 ( .DIN1(n10809), .DIN2(n10819), .Q(n10648) );
  nnd2s1 U11739 ( .DIN1(n10819), .DIN2(n11619), .Q(n11616) );
  nnd2s1 U11740 ( .DIN1(n10831), .DIN2(n11132), .Q(n11619) );
  nnd2s1 U11741 ( .DIN1(n10492), .DIN2(n11620), .Q(n11615) );
  nnd2s1 U11742 ( .DIN1(n10832), .DIN2(n10518), .Q(n11620) );
  nnd2s1 U11743 ( .DIN1(n10507), .DIN2(n11121), .Q(n11614) );
  or3s1 U11744 ( .DIN1(n11621), .DIN2(n11622), .DIN3(n11623), .Q(n5425) );
  nnd4s1 U11745 ( .DIN1(n11624), .DIN2(n11625), .DIN3(n10656), .DIN4(n11626), 
        .Q(n11623) );
  and3s1 U11746 ( .DIN1(n10859), .DIN2(n11192), .DIN3(n11159), .Q(n11626) );
  nor4s1 U11747 ( .DIN1(n11627), .DIN2(n11628), .DIN3(n11629), .DIN4(n11630), 
        .Q(n11159) );
  nnd4s1 U11748 ( .DIN1(n11631), .DIN2(n11632), .DIN3(n11633), .DIN4(n11634), 
        .Q(n11630) );
  nnd2s1 U11749 ( .DIN1(n10878), .DIN2(n10681), .Q(n11634) );
  nor2s1 U11750 ( .DIN1(n11635), .DIN2(n11636), .Q(n11633) );
  nor2s1 U11751 ( .DIN1(n10680), .DIN2(n11637), .Q(n11636) );
  nor2s1 U11752 ( .DIN1(n11638), .DIN2(n10912), .Q(n11635) );
  nnd2s1 U11753 ( .DIN1(n10867), .DIN2(n10879), .Q(n11632) );
  nnd2s1 U11754 ( .DIN1(n10887), .DIN2(n10672), .Q(n11631) );
  nnd3s1 U11755 ( .DIN1(n11639), .DIN2(n11640), .DIN3(n11641), .Q(n11629) );
  nnd2s1 U11756 ( .DIN1(n10913), .DIN2(n10918), .Q(n11641) );
  nnd2s1 U11757 ( .DIN1(n11642), .DIN2(n11643), .Q(n11640) );
  nnd3s1 U11758 ( .DIN1(n11184), .DIN2(n11637), .DIN3(n11218), .Q(n11643) );
  nnd2s1 U11759 ( .DIN1(n11199), .DIN2(n11644), .Q(n11639) );
  nnd3s1 U11760 ( .DIN1(n10874), .DIN2(n10670), .DIN3(n10679), .Q(n11644) );
  nor2s1 U11761 ( .DIN1(n10874), .DIN2(n11220), .Q(n11628) );
  nor2s1 U11762 ( .DIN1(n11645), .DIN2(n11646), .Q(n11627) );
  nor4s1 U11763 ( .DIN1(n11647), .DIN2(n11648), .DIN3(n11649), .DIN4(n11650), 
        .Q(n11192) );
  nnd4s1 U11764 ( .DIN1(n11651), .DIN2(n11652), .DIN3(n11653), .DIN4(n11654), 
        .Q(n11650) );
  nor2s1 U11765 ( .DIN1(n11655), .DIN2(n11656), .Q(n11654) );
  nor2s1 U11766 ( .DIN1(n11637), .DIN2(n11646), .Q(n11656) );
  nor2s1 U11767 ( .DIN1(n10916), .DIN2(n10670), .Q(n11655) );
  nnd2s1 U11768 ( .DIN1(n10664), .DIN2(n10910), .Q(n11652) );
  nnd2s1 U11769 ( .DIN1(n10865), .DIN2(n10662), .Q(n11651) );
  nnd3s1 U11770 ( .DIN1(n11657), .DIN2(n11658), .DIN3(n11659), .Q(n11649) );
  nnd2s1 U11771 ( .DIN1(n10876), .DIN2(n11660), .Q(n11659) );
  nnd2s1 U11772 ( .DIN1(n11219), .DIN2(n10892), .Q(n11660) );
  nnd2s1 U11773 ( .DIN1(n10661), .DIN2(n11661), .Q(n11658) );
  nnd2s1 U11774 ( .DIN1(n11244), .DIN2(n11184), .Q(n11661) );
  nnd2s1 U11775 ( .DIN1(n10884), .DIN2(n10914), .Q(n11657) );
  nnd2s1 U11776 ( .DIN1(n10895), .DIN2(n11185), .Q(n10914) );
  nor2s1 U11777 ( .DIN1(n11662), .DIN2(n10684), .Q(n11648) );
  nor2s1 U11778 ( .DIN1(n10663), .DIN2(n10893), .Q(n11662) );
  nor2s1 U11779 ( .DIN1(n11663), .DIN2(n11216), .Q(n11647) );
  and2s1 U11780 ( .DIN1(n10874), .DIN2(n11664), .Q(n11663) );
  nor4s1 U11781 ( .DIN1(n11665), .DIN2(n11666), .DIN3(n11667), .DIN4(n11668), 
        .Q(n10859) );
  nnd4s1 U11782 ( .DIN1(n11669), .DIN2(n11670), .DIN3(n11671), .DIN4(n11672), 
        .Q(n11668) );
  nnd2s1 U11783 ( .DIN1(n11198), .DIN2(n10879), .Q(n11672) );
  nor2s1 U11784 ( .DIN1(n11673), .DIN2(n11674), .Q(n11671) );
  nor2s1 U11785 ( .DIN1(n11675), .DIN2(n10684), .Q(n11673) );
  nnd2s1 U11786 ( .DIN1(n10877), .DIN2(n10887), .Q(n11670) );
  nnd2s1 U11787 ( .DIN1(n10866), .DIN2(n11242), .Q(n11669) );
  nnd3s1 U11788 ( .DIN1(n11676), .DIN2(n11677), .DIN3(n11678), .Q(n11667) );
  nnd2s1 U11789 ( .DIN1(n10662), .DIN2(n11679), .Q(n11678) );
  nnd2s1 U11790 ( .DIN1(n10672), .DIN2(n11680), .Q(n11677) );
  nnd2s1 U11791 ( .DIN1(n11216), .DIN2(n11184), .Q(n11680) );
  nnd2s1 U11792 ( .DIN1(n11199), .DIN2(n11681), .Q(n11676) );
  nnd3s1 U11793 ( .DIN1(n11188), .DIN2(n11646), .DIN3(n11682), .Q(n11681) );
  nor2s1 U11794 ( .DIN1(n10670), .DIN2(n11220), .Q(n11666) );
  nor2s1 U11795 ( .DIN1(n10687), .DIN2(n10917), .Q(n11665) );
  nor3s1 U11796 ( .DIN1(n11683), .DIN2(n11684), .DIN3(n11685), .Q(n10656) );
  nnd4s1 U11797 ( .DIN1(n11193), .DIN2(n10861), .DIN3(n11163), .DIN4(n11686), 
        .Q(n11685) );
  and3s1 U11798 ( .DIN1(n11687), .DIN2(n11688), .DIN3(n11689), .Q(n11686) );
  nnd2s1 U11799 ( .DIN1(n10866), .DIN2(n11174), .Q(n11689) );
  nnd2s1 U11800 ( .DIN1(n10904), .DIN2(n10681), .Q(n11687) );
  nor4s1 U11801 ( .DIN1(n11690), .DIN2(n11691), .DIN3(n11692), .DIN4(n11693), 
        .Q(n11163) );
  nnd4s1 U11802 ( .DIN1(n11694), .DIN2(n11695), .DIN3(n11696), .DIN4(n11697), 
        .Q(n11693) );
  nnd2s1 U11803 ( .DIN1(n10866), .DIN2(n11698), .Q(n11697) );
  nnd2s1 U11804 ( .DIN1(n11699), .DIN2(n11188), .Q(n11698) );
  nor2s1 U11805 ( .DIN1(n11700), .DIN2(n11701), .Q(n11696) );
  nor2s1 U11806 ( .DIN1(n11702), .DIN2(n10916), .Q(n11701) );
  nor2s1 U11807 ( .DIN1(n10904), .DIN2(n10689), .Q(n11702) );
  nor2s1 U11808 ( .DIN1(n11703), .DIN2(n11704), .Q(n11700) );
  nor2s1 U11809 ( .DIN1(n11705), .DIN2(n10865), .Q(n11703) );
  nnd2s1 U11810 ( .DIN1(n11242), .DIN2(n11706), .Q(n11695) );
  nnd3s1 U11811 ( .DIN1(n11675), .DIN2(n11215), .DIN3(n11220), .Q(n11706) );
  nnd2s1 U11812 ( .DIN1(n11199), .DIN2(n11705), .Q(n11694) );
  nnd3s1 U11813 ( .DIN1(n11707), .DIN2(n11708), .DIN3(n11709), .Q(n11692) );
  nnd2s1 U11814 ( .DIN1(n10913), .DIN2(n11710), .Q(n11709) );
  nnd2s1 U11815 ( .DIN1(n11172), .DIN2(n11642), .Q(n11708) );
  nnd2s1 U11816 ( .DIN1(n10661), .DIN2(n10884), .Q(n11707) );
  nor2s1 U11817 ( .DIN1(n11637), .DIN2(n10684), .Q(n11691) );
  nor2s1 U11818 ( .DIN1(n11244), .DIN2(n11646), .Q(n11690) );
  nor4s1 U11819 ( .DIN1(n11711), .DIN2(n11712), .DIN3(n11713), .DIN4(n11714), 
        .Q(n10861) );
  nnd4s1 U11820 ( .DIN1(n11715), .DIN2(n11716), .DIN3(n11717), .DIN4(n11718), 
        .Q(n11714) );
  nnd2s1 U11821 ( .DIN1(n11174), .DIN2(n10910), .Q(n11718) );
  nnd2s1 U11822 ( .DIN1(n10681), .DIN2(n10876), .Q(n11717) );
  nnd2s1 U11823 ( .DIN1(n10901), .DIN2(n11242), .Q(n11716) );
  nnd2s1 U11824 ( .DIN1(n10877), .DIN2(n10866), .Q(n11715) );
  nnd3s1 U11825 ( .DIN1(n11719), .DIN2(n11720), .DIN3(n11721), .Q(n11713) );
  nnd2s1 U11826 ( .DIN1(n10685), .DIN2(n11722), .Q(n11721) );
  nnd3s1 U11827 ( .DIN1(n10889), .DIN2(n11185), .DIN3(n10684), .Q(n11722) );
  nnd2s1 U11828 ( .DIN1(n10905), .DIN2(n11723), .Q(n11720) );
  nnd2s1 U11829 ( .DIN1(n11664), .DIN2(n10889), .Q(n11723) );
  nor2s1 U11830 ( .DIN1(n11710), .DIN2(n11705), .Q(n11664) );
  nnd2s1 U11831 ( .DIN1(n11198), .DIN2(n11724), .Q(n11719) );
  nnd2s1 U11832 ( .DIN1(n11638), .DIN2(n11244), .Q(n11724) );
  nor2s1 U11833 ( .DIN1(n11188), .DIN2(n11219), .Q(n11712) );
  nor2s1 U11834 ( .DIN1(n10896), .DIN2(n11216), .Q(n11711) );
  hi1s1 U11835 ( .DIN(n11725), .Q(n10896) );
  nor2s1 U11836 ( .DIN1(n11726), .DIN2(n11727), .Q(n11193) );
  nnd4s1 U11837 ( .DIN1(n11728), .DIN2(n11729), .DIN3(n11730), .DIN4(n11731), 
        .Q(n11727) );
  nnd2s1 U11838 ( .DIN1(n11174), .DIN2(n11732), .Q(n11731) );
  nnd3s1 U11839 ( .DIN1(n11216), .DIN2(n11637), .DIN3(n11675), .Q(n11732) );
  nnd2s1 U11840 ( .DIN1(n11172), .DIN2(n10865), .Q(n11729) );
  nnd4s1 U11841 ( .DIN1(n11733), .DIN2(n11734), .DIN3(n11735), .DIN4(n11736), 
        .Q(n11726) );
  nnd2s1 U11842 ( .DIN1(n10910), .DIN2(n11737), .Q(n11736) );
  nnd2s1 U11843 ( .DIN1(n11738), .DIN2(n10684), .Q(n11737) );
  nnd2s1 U11844 ( .DIN1(n10663), .DIN2(n11739), .Q(n11735) );
  nnd2s1 U11845 ( .DIN1(n10672), .DIN2(n11740), .Q(n11734) );
  nnd2s1 U11846 ( .DIN1(n11219), .DIN2(n11675), .Q(n11740) );
  nnd2s1 U11847 ( .DIN1(n11198), .DIN2(n11741), .Q(n11733) );
  nnd2s1 U11848 ( .DIN1(n10669), .DIN2(n11215), .Q(n11741) );
  nnd3s1 U11849 ( .DIN1(n11742), .DIN2(n11743), .DIN3(n11744), .Q(n11684) );
  nnd2s1 U11850 ( .DIN1(n10662), .DIN2(n11242), .Q(n11744) );
  nnd2s1 U11851 ( .DIN1(n11705), .DIN2(n11745), .Q(n11743) );
  nnd3s1 U11852 ( .DIN1(n11220), .DIN2(n11637), .DIN3(n11746), .Q(n11745) );
  or2s1 U11853 ( .DIN1(n10889), .DIN2(n11747), .Q(n11742) );
  nnd3s1 U11854 ( .DIN1(n11748), .DIN2(n11749), .DIN3(n11750), .Q(n11683) );
  nnd2s1 U11855 ( .DIN1(n10672), .DIN2(n11751), .Q(n11750) );
  nnd2s1 U11856 ( .DIN1(n11225), .DIN2(n11218), .Q(n11751) );
  nnd2s1 U11857 ( .DIN1(n10887), .DIN2(n11752), .Q(n11749) );
  or2s1 U11858 ( .DIN1(n10918), .DIN2(n11642), .Q(n11752) );
  nnd2s1 U11859 ( .DIN1(n10684), .DIN2(n10668), .Q(n10918) );
  nnd2s1 U11860 ( .DIN1(n10913), .DIN2(n11753), .Q(n11748) );
  nnd2s1 U11861 ( .DIN1(n11180), .DIN2(n10874), .Q(n11753) );
  nnd2s1 U11862 ( .DIN1(n10681), .DIN2(n10664), .Q(n11625) );
  nnd2s1 U11863 ( .DIN1(n10877), .DIN2(n10893), .Q(n11624) );
  nnd3s1 U11864 ( .DIN1(n11754), .DIN2(n11755), .DIN3(n11756), .Q(n11622) );
  nnd2s1 U11865 ( .DIN1(n11710), .DIN2(n10910), .Q(n11756) );
  nnd2s1 U11866 ( .DIN1(n11173), .DIN2(n11757), .Q(n11755) );
  nnd4s1 U11867 ( .DIN1(n11758), .DIN2(n11759), .DIN3(n11760), .DIN4(n11761), 
        .Q(n11621) );
  nnd2s1 U11868 ( .DIN1(n10905), .DIN2(n11762), .Q(n11761) );
  nnd2s1 U11869 ( .DIN1(n10687), .DIN2(n10912), .Q(n11762) );
  nor2s1 U11870 ( .DIN1(n10865), .DIN2(n10876), .Q(n10687) );
  nnd2s1 U11871 ( .DIN1(n10876), .DIN2(n11763), .Q(n11760) );
  nnd2s1 U11872 ( .DIN1(n10891), .DIN2(n11218), .Q(n11763) );
  nnd2s1 U11873 ( .DIN1(n10867), .DIN2(n11764), .Q(n11759) );
  nnd2s1 U11874 ( .DIN1(n10892), .DIN2(n11220), .Q(n11764) );
  nnd2s1 U11875 ( .DIN1(n11242), .DIN2(n11207), .Q(n11758) );
  xor2s1 U11876 ( .DIN1(n5048), .DIN2(n11765), .Q(n11475) );
  xor2s1 U11877 ( .DIN1(w1[3]), .DIN2(n10443), .Q(n11765) );
  hi1s1 U11878 ( .DIN(n5024), .Q(n10443) );
  or3s1 U11879 ( .DIN1(n11766), .DIN2(n11767), .DIN3(n11768), .Q(n5024) );
  nnd4s1 U11880 ( .DIN1(n11769), .DIN2(n11770), .DIN3(n11771), .DIN4(n11772), 
        .Q(n11768) );
  and3s1 U11881 ( .DIN1(n11773), .DIN2(n11774), .DIN3(n11775), .Q(n11772) );
  nnd2s1 U11882 ( .DIN1(n10710), .DIN2(n10717), .Q(n11774) );
  nnd2s1 U11883 ( .DIN1(n10703), .DIN2(n10533), .Q(n11773) );
  nnd3s1 U11884 ( .DIN1(n11776), .DIN2(n11777), .DIN3(n11778), .Q(n11767) );
  nnd2s1 U11885 ( .DIN1(n10937), .DIN2(n10701), .Q(n11778) );
  or2s1 U11886 ( .DIN1(n10961), .DIN2(n11779), .Q(n11777) );
  nnd2s1 U11887 ( .DIN1(n10990), .DIN2(n10752), .Q(n11776) );
  nnd4s1 U11888 ( .DIN1(n11780), .DIN2(n11781), .DIN3(n11782), .DIN4(n11783), 
        .Q(n11766) );
  nnd2s1 U11889 ( .DIN1(n11329), .DIN2(n11784), .Q(n11783) );
  nnd2s1 U11890 ( .DIN1(n11369), .DIN2(n10932), .Q(n11784) );
  nnd2s1 U11891 ( .DIN1(n10716), .DIN2(n11785), .Q(n11782) );
  nnd2s1 U11892 ( .DIN1(n10963), .DIN2(n10548), .Q(n11785) );
  nor2s1 U11893 ( .DIN1(n10952), .DIN2(n10951), .Q(n10963) );
  nnd2s1 U11894 ( .DIN1(n10744), .DIN2(n11786), .Q(n11781) );
  nnd2s1 U11895 ( .DIN1(n10756), .DIN2(n10933), .Q(n11786) );
  nnd2s1 U11896 ( .DIN1(n10550), .DIN2(n11787), .Q(n11780) );
  or3s1 U11897 ( .DIN1(n11788), .DIN2(n11789), .DIN3(n11790), .Q(n5048) );
  nnd4s1 U11898 ( .DIN1(n11791), .DIN2(n11792), .DIN3(n10765), .DIN4(n11793), 
        .Q(n11790) );
  and3s1 U11899 ( .DIN1(n11013), .DIN2(n11421), .DIN3(n11391), .Q(n11793) );
  nor4s1 U11900 ( .DIN1(n11794), .DIN2(n11795), .DIN3(n11796), .DIN4(n11797), 
        .Q(n11391) );
  nnd4s1 U11901 ( .DIN1(n11798), .DIN2(n11799), .DIN3(n11800), .DIN4(n11801), 
        .Q(n11797) );
  nnd2s1 U11902 ( .DIN1(n10583), .DIN2(n10786), .Q(n11801) );
  nor2s1 U11903 ( .DIN1(n11802), .DIN2(n11803), .Q(n11800) );
  nor2s1 U11904 ( .DIN1(n10785), .DIN2(n11804), .Q(n11803) );
  nor2s1 U11905 ( .DIN1(n11805), .DIN2(n11059), .Q(n11802) );
  nnd2s1 U11906 ( .DIN1(n10573), .DIN2(n11030), .Q(n11799) );
  nnd2s1 U11907 ( .DIN1(n11037), .DIN2(n10596), .Q(n11798) );
  nnd3s1 U11908 ( .DIN1(n11806), .DIN2(n11807), .DIN3(n11808), .Q(n11796) );
  nnd2s1 U11909 ( .DIN1(n11060), .DIN2(n11064), .Q(n11808) );
  nnd2s1 U11910 ( .DIN1(n10581), .DIN2(n11809), .Q(n11807) );
  nnd3s1 U11911 ( .DIN1(n11413), .DIN2(n11804), .DIN3(n11447), .Q(n11809) );
  nnd2s1 U11912 ( .DIN1(n11428), .DIN2(n11810), .Q(n11806) );
  nnd3s1 U11913 ( .DIN1(n11027), .DIN2(n10595), .DIN3(n10784), .Q(n11810) );
  nor2s1 U11914 ( .DIN1(n11027), .DIN2(n10599), .Q(n11795) );
  nor2s1 U11915 ( .DIN1(n11811), .DIN2(n11812), .Q(n11794) );
  nor4s1 U11916 ( .DIN1(n11813), .DIN2(n11814), .DIN3(n11815), .DIN4(n11816), 
        .Q(n11421) );
  nnd4s1 U11917 ( .DIN1(n11817), .DIN2(n11818), .DIN3(n11819), .DIN4(n11820), 
        .Q(n11816) );
  nor2s1 U11918 ( .DIN1(n11821), .DIN2(n11822), .Q(n11820) );
  nor2s1 U11919 ( .DIN1(n11804), .DIN2(n11812), .Q(n11822) );
  nor2s1 U11920 ( .DIN1(n11063), .DIN2(n10595), .Q(n11821) );
  nnd2s1 U11921 ( .DIN1(n10771), .DIN2(n10600), .Q(n11818) );
  nnd2s1 U11922 ( .DIN1(n11019), .DIN2(n10580), .Q(n11817) );
  nnd3s1 U11923 ( .DIN1(n11823), .DIN2(n11824), .DIN3(n11825), .Q(n11815) );
  nnd2s1 U11924 ( .DIN1(n11029), .DIN2(n11826), .Q(n11825) );
  nnd2s1 U11925 ( .DIN1(n11448), .DIN2(n11042), .Q(n11826) );
  nnd2s1 U11926 ( .DIN1(n10770), .DIN2(n11827), .Q(n11824) );
  nnd2s1 U11927 ( .DIN1(n11470), .DIN2(n11413), .Q(n11827) );
  nnd2s1 U11928 ( .DIN1(n10582), .DIN2(n11061), .Q(n11823) );
  nnd2s1 U11929 ( .DIN1(n11044), .DIN2(n11414), .Q(n11061) );
  nor2s1 U11930 ( .DIN1(n11828), .DIN2(n10789), .Q(n11814) );
  nor2s1 U11931 ( .DIN1(n10571), .DIN2(n10592), .Q(n11828) );
  nor2s1 U11932 ( .DIN1(n11829), .DIN2(n11445), .Q(n11813) );
  and2s1 U11933 ( .DIN1(n11027), .DIN2(n11830), .Q(n11829) );
  nor4s1 U11934 ( .DIN1(n11831), .DIN2(n11832), .DIN3(n11833), .DIN4(n11834), 
        .Q(n11013) );
  nnd4s1 U11935 ( .DIN1(n11835), .DIN2(n11836), .DIN3(n11837), .DIN4(n11838), 
        .Q(n11834) );
  nnd2s1 U11936 ( .DIN1(n11427), .DIN2(n11030), .Q(n11838) );
  nor2s1 U11937 ( .DIN1(n11839), .DIN2(n11840), .Q(n11837) );
  nor2s1 U11938 ( .DIN1(n11841), .DIN2(n10789), .Q(n11839) );
  nnd2s1 U11939 ( .DIN1(n11018), .DIN2(n11037), .Q(n11836) );
  nnd2s1 U11940 ( .DIN1(n11020), .DIN2(n10588), .Q(n11835) );
  nnd3s1 U11941 ( .DIN1(n11842), .DIN2(n11843), .DIN3(n11844), .Q(n11833) );
  nnd2s1 U11942 ( .DIN1(n10580), .DIN2(n11845), .Q(n11844) );
  nnd2s1 U11943 ( .DIN1(n10596), .DIN2(n11846), .Q(n11843) );
  nnd2s1 U11944 ( .DIN1(n11445), .DIN2(n11413), .Q(n11846) );
  nnd2s1 U11945 ( .DIN1(n11428), .DIN2(n11847), .Q(n11842) );
  nnd3s1 U11946 ( .DIN1(n11417), .DIN2(n11812), .DIN3(n11848), .Q(n11847) );
  nor2s1 U11947 ( .DIN1(n10595), .DIN2(n10599), .Q(n11832) );
  nor2s1 U11948 ( .DIN1(n10791), .DIN2(n10591), .Q(n11831) );
  nor3s1 U11949 ( .DIN1(n11849), .DIN2(n11850), .DIN3(n11851), .Q(n10765) );
  nnd4s1 U11950 ( .DIN1(n11422), .DIN2(n11015), .DIN3(n11395), .DIN4(n11852), 
        .Q(n11851) );
  and3s1 U11951 ( .DIN1(n11853), .DIN2(n11854), .DIN3(n11855), .Q(n11852) );
  nnd2s1 U11952 ( .DIN1(n11020), .DIN2(n10579), .Q(n11855) );
  nnd2s1 U11953 ( .DIN1(n10570), .DIN2(n10786), .Q(n11853) );
  nor4s1 U11954 ( .DIN1(n11856), .DIN2(n11857), .DIN3(n11858), .DIN4(n11859), 
        .Q(n11395) );
  nnd4s1 U11955 ( .DIN1(n11860), .DIN2(n11861), .DIN3(n11862), .DIN4(n11863), 
        .Q(n11859) );
  nnd2s1 U11956 ( .DIN1(n11020), .DIN2(n11864), .Q(n11863) );
  nnd2s1 U11957 ( .DIN1(n11865), .DIN2(n11417), .Q(n11864) );
  nor2s1 U11958 ( .DIN1(n11866), .DIN2(n11867), .Q(n11862) );
  nor2s1 U11959 ( .DIN1(n11868), .DIN2(n11063), .Q(n11867) );
  nor2s1 U11960 ( .DIN1(n10570), .DIN2(n10793), .Q(n11868) );
  nor2s1 U11961 ( .DIN1(n11869), .DIN2(n10598), .Q(n11866) );
  nor2s1 U11962 ( .DIN1(n11870), .DIN2(n11019), .Q(n11869) );
  nnd2s1 U11963 ( .DIN1(n10588), .DIN2(n11871), .Q(n11861) );
  nnd3s1 U11964 ( .DIN1(n11841), .DIN2(n11444), .DIN3(n10599), .Q(n11871) );
  nnd2s1 U11965 ( .DIN1(n11428), .DIN2(n11870), .Q(n11860) );
  nnd3s1 U11966 ( .DIN1(n11872), .DIN2(n11873), .DIN3(n11874), .Q(n11858) );
  nnd2s1 U11967 ( .DIN1(n11060), .DIN2(n11875), .Q(n11874) );
  nnd2s1 U11968 ( .DIN1(n10578), .DIN2(n10581), .Q(n11873) );
  nnd2s1 U11969 ( .DIN1(n10770), .DIN2(n10582), .Q(n11872) );
  nor2s1 U11970 ( .DIN1(n11804), .DIN2(n10789), .Q(n11857) );
  nor2s1 U11971 ( .DIN1(n11470), .DIN2(n11812), .Q(n11856) );
  nor4s1 U11972 ( .DIN1(n11876), .DIN2(n11877), .DIN3(n11878), .DIN4(n11879), 
        .Q(n11015) );
  nnd4s1 U11973 ( .DIN1(n11880), .DIN2(n11881), .DIN3(n11882), .DIN4(n11883), 
        .Q(n11879) );
  nnd2s1 U11974 ( .DIN1(n10579), .DIN2(n10600), .Q(n11883) );
  nnd2s1 U11975 ( .DIN1(n10786), .DIN2(n11029), .Q(n11882) );
  nnd2s1 U11976 ( .DIN1(n11050), .DIN2(n10588), .Q(n11881) );
  nnd2s1 U11977 ( .DIN1(n11018), .DIN2(n11020), .Q(n11880) );
  nnd3s1 U11978 ( .DIN1(n11884), .DIN2(n11885), .DIN3(n11886), .Q(n11878) );
  nnd2s1 U11979 ( .DIN1(n10572), .DIN2(n11887), .Q(n11886) );
  nnd3s1 U11980 ( .DIN1(n11039), .DIN2(n11414), .DIN3(n10789), .Q(n11887) );
  nnd2s1 U11981 ( .DIN1(n11053), .DIN2(n11888), .Q(n11885) );
  nnd2s1 U11982 ( .DIN1(n11830), .DIN2(n11039), .Q(n11888) );
  nor2s1 U11983 ( .DIN1(n11875), .DIN2(n11870), .Q(n11830) );
  nnd2s1 U11984 ( .DIN1(n11427), .DIN2(n11889), .Q(n11884) );
  nnd2s1 U11985 ( .DIN1(n11805), .DIN2(n11470), .Q(n11889) );
  nor2s1 U11986 ( .DIN1(n11417), .DIN2(n11448), .Q(n11877) );
  nor2s1 U11987 ( .DIN1(n11045), .DIN2(n11445), .Q(n11876) );
  hi1s1 U11988 ( .DIN(n10601), .Q(n11045) );
  nor2s1 U11989 ( .DIN1(n11890), .DIN2(n11891), .Q(n11422) );
  nnd4s1 U11990 ( .DIN1(n11892), .DIN2(n11893), .DIN3(n11894), .DIN4(n11895), 
        .Q(n11891) );
  nnd2s1 U11991 ( .DIN1(n10579), .DIN2(n11896), .Q(n11895) );
  nnd3s1 U11992 ( .DIN1(n11445), .DIN2(n11804), .DIN3(n11841), .Q(n11896) );
  nnd2s1 U11993 ( .DIN1(n10578), .DIN2(n11019), .Q(n11893) );
  nnd4s1 U11994 ( .DIN1(n11897), .DIN2(n11898), .DIN3(n11899), .DIN4(n11900), 
        .Q(n11890) );
  nnd2s1 U11995 ( .DIN1(n10600), .DIN2(n11901), .Q(n11900) );
  nnd2s1 U11996 ( .DIN1(n11902), .DIN2(n10789), .Q(n11901) );
  nnd2s1 U11997 ( .DIN1(n10571), .DIN2(n11903), .Q(n11899) );
  nnd2s1 U11998 ( .DIN1(n10596), .DIN2(n11904), .Q(n11898) );
  nnd2s1 U11999 ( .DIN1(n11448), .DIN2(n11841), .Q(n11904) );
  nnd2s1 U12000 ( .DIN1(n11427), .DIN2(n11905), .Q(n11897) );
  nnd2s1 U12001 ( .DIN1(n10776), .DIN2(n11444), .Q(n11905) );
  nnd3s1 U12002 ( .DIN1(n11906), .DIN2(n11907), .DIN3(n11908), .Q(n11850) );
  nnd2s1 U12003 ( .DIN1(n10580), .DIN2(n10588), .Q(n11908) );
  nnd2s1 U12004 ( .DIN1(n11870), .DIN2(n11909), .Q(n11907) );
  nnd3s1 U12005 ( .DIN1(n10599), .DIN2(n11804), .DIN3(n11910), .Q(n11909) );
  or2s1 U12006 ( .DIN1(n11039), .DIN2(n11911), .Q(n11906) );
  nnd3s1 U12007 ( .DIN1(n11912), .DIN2(n11913), .DIN3(n11914), .Q(n11849) );
  nnd2s1 U12008 ( .DIN1(n10596), .DIN2(n11915), .Q(n11914) );
  nnd2s1 U12009 ( .DIN1(n11452), .DIN2(n11447), .Q(n11915) );
  nnd2s1 U12010 ( .DIN1(n11037), .DIN2(n11916), .Q(n11913) );
  or2s1 U12011 ( .DIN1(n11064), .DIN2(n10581), .Q(n11916) );
  nnd2s1 U12012 ( .DIN1(n10789), .DIN2(n10775), .Q(n11064) );
  nnd2s1 U12013 ( .DIN1(n11060), .DIN2(n11917), .Q(n11912) );
  nnd2s1 U12014 ( .DIN1(n10594), .DIN2(n11027), .Q(n11917) );
  nnd2s1 U12015 ( .DIN1(n10786), .DIN2(n10771), .Q(n11792) );
  nnd2s1 U12016 ( .DIN1(n11018), .DIN2(n10592), .Q(n11791) );
  nnd3s1 U12017 ( .DIN1(n11918), .DIN2(n11919), .DIN3(n11920), .Q(n11789) );
  nnd2s1 U12018 ( .DIN1(n11875), .DIN2(n10600), .Q(n11920) );
  nnd2s1 U12019 ( .DIN1(n11404), .DIN2(n11921), .Q(n11919) );
  nnd4s1 U12020 ( .DIN1(n11922), .DIN2(n11923), .DIN3(n11924), .DIN4(n11925), 
        .Q(n11788) );
  nnd2s1 U12021 ( .DIN1(n11053), .DIN2(n11926), .Q(n11925) );
  nnd2s1 U12022 ( .DIN1(n10791), .DIN2(n11059), .Q(n11926) );
  nor2s1 U12023 ( .DIN1(n11019), .DIN2(n11029), .Q(n10791) );
  nnd2s1 U12024 ( .DIN1(n11029), .DIN2(n11927), .Q(n11924) );
  nnd2s1 U12025 ( .DIN1(n11041), .DIN2(n11447), .Q(n11927) );
  nnd2s1 U12026 ( .DIN1(n10573), .DIN2(n11928), .Q(n11923) );
  nnd2s1 U12027 ( .DIN1(n11042), .DIN2(n10599), .Q(n11928) );
  nnd2s1 U12028 ( .DIN1(n10588), .DIN2(n11436), .Q(n11922) );
  nnd2s1 U12029 ( .DIN1(n11929), .DIN2(n1600), .Q(n11472) );
  xor2s1 U12030 ( .DIN1(w1[3]), .DIN2(text_in_r[67]), .Q(n11929) );
  nnd3s1 U12031 ( .DIN1(n11930), .DIN2(n11931), .DIN3(n11932), .Q(N164) );
  nnd2s1 U12032 ( .DIN1(n1598), .DIN2(n11933), .Q(n11932) );
  xor2s1 U12033 ( .DIN1(w1[2]), .DIN2(text_in_r[66]), .Q(n11933) );
  nnd2s1 U12034 ( .DIN1(n11934), .DIN2(n5423), .Q(n11931) );
  nnd2s1 U12035 ( .DIN1(n11935), .DIN2(n11936), .Q(n11934) );
  nnd2s1 U12036 ( .DIN1(n10285), .DIN2(n11937), .Q(n11936) );
  nnd2s1 U12037 ( .DIN1(n11938), .DIN2(n10287), .Q(n11935) );
  nnd2s1 U12038 ( .DIN1(n11939), .DIN2(n11940), .Q(n11930) );
  nnd2s1 U12039 ( .DIN1(n11941), .DIN2(n11942), .Q(n11940) );
  nnd2s1 U12040 ( .DIN1(n10287), .DIN2(n11937), .Q(n11942) );
  nor2s1 U12041 ( .DIN1(n10450), .DIN2(n1595), .Q(n10287) );
  nnd2s1 U12042 ( .DIN1(n11938), .DIN2(n10285), .Q(n11941) );
  nor2s1 U12043 ( .DIN1(n11943), .DIN2(n1596), .Q(n10285) );
  hi1s1 U12044 ( .DIN(n10450), .Q(n11943) );
  xor2s1 U12045 ( .DIN1(n5424), .DIN2(n5071), .Q(n10450) );
  hi1s1 U12046 ( .DIN(n10301), .Q(n5071) );
  or3s1 U12047 ( .DIN1(n11944), .DIN2(n11945), .DIN3(n11946), .Q(n10301) );
  nnd4s1 U12048 ( .DIN1(n11947), .DIN2(n11948), .DIN3(n10483), .DIN4(n11949), 
        .Q(n11946) );
  and3s1 U12049 ( .DIN1(n11950), .DIN2(n11951), .DIN3(n11952), .Q(n11949) );
  nnd2s1 U12050 ( .DIN1(n10511), .DIN2(n10502), .Q(n11951) );
  nnd2s1 U12051 ( .DIN1(n10507), .DIN2(n10820), .Q(n11950) );
  nor3s1 U12052 ( .DIN1(n11953), .DIN2(n11954), .DIN3(n11955), .Q(n10483) );
  nnd4s1 U12053 ( .DIN1(n11956), .DIN2(n11957), .DIN3(n11958), .DIN4(n11959), 
        .Q(n11955) );
  and3s1 U12054 ( .DIN1(n11960), .DIN2(n11961), .DIN3(n11962), .Q(n11959) );
  nnd2s1 U12055 ( .DIN1(n10639), .DIN2(n10492), .Q(n11962) );
  nnd2s1 U12056 ( .DIN1(n10808), .DIN2(n10497), .Q(n11961) );
  nnd2s1 U12057 ( .DIN1(n10511), .DIN2(n10819), .Q(n11960) );
  nnd3s1 U12058 ( .DIN1(n11963), .DIN2(n11964), .DIN3(n11586), .Q(n11954) );
  nnd2s1 U12059 ( .DIN1(n10810), .DIN2(n11562), .Q(n11586) );
  or2s1 U12060 ( .DIN1(n10517), .DIN2(n11594), .Q(n11964) );
  nor2s1 U12061 ( .DIN1(n10489), .DIN2(n10500), .Q(n11594) );
  nnd2s1 U12062 ( .DIN1(n10843), .DIN2(n10650), .Q(n11963) );
  nnd2s1 U12063 ( .DIN1(n10834), .DIN2(n10641), .Q(n10650) );
  nnd4s1 U12064 ( .DIN1(n11965), .DIN2(n11966), .DIN3(n11967), .DIN4(n11968), 
        .Q(n11953) );
  nnd2s1 U12065 ( .DIN1(n11089), .DIN2(n11969), .Q(n11968) );
  nnd2s1 U12066 ( .DIN1(n10491), .DIN2(n11970), .Q(n11967) );
  nnd2s1 U12067 ( .DIN1(n10641), .DIN2(n10849), .Q(n11970) );
  nnd2s1 U12068 ( .DIN1(n10809), .DIN2(n11971), .Q(n11966) );
  nnd2s1 U12069 ( .DIN1(n10832), .DIN2(n10510), .Q(n11971) );
  nnd2s1 U12070 ( .DIN1(n10515), .DIN2(n11972), .Q(n11965) );
  nnd2s1 U12071 ( .DIN1(n11602), .DIN2(n11496), .Q(n11972) );
  hi1s1 U12072 ( .DIN(n10842), .Q(n11602) );
  nnd2s1 U12073 ( .DIN1(n11129), .DIN2(n10853), .Q(n10842) );
  nnd3s1 U12074 ( .DIN1(n11973), .DIN2(n11974), .DIN3(n11975), .Q(n11945) );
  nnd2s1 U12075 ( .DIN1(n10808), .DIN2(n10499), .Q(n11975) );
  or2s1 U12076 ( .DIN1(n10513), .DIN2(n10509), .Q(n11974) );
  nor2s1 U12077 ( .DIN1(n10639), .DIN2(n10643), .Q(n10509) );
  nnd2s1 U12078 ( .DIN1(n11112), .DIN2(n10519), .Q(n11973) );
  nnd4s1 U12079 ( .DIN1(n11976), .DIN2(n11977), .DIN3(n11978), .DIN4(n11979), 
        .Q(n11944) );
  nnd2s1 U12080 ( .DIN1(n11567), .DIN2(n11980), .Q(n11979) );
  nnd2s1 U12081 ( .DIN1(n11603), .DIN2(n11129), .Q(n11980) );
  nnd2s1 U12082 ( .DIN1(n10490), .DIN2(n11981), .Q(n11978) );
  nnd2s1 U12083 ( .DIN1(n11096), .DIN2(n10642), .Q(n11981) );
  nor2s1 U12084 ( .DIN1(n10498), .DIN2(n11562), .Q(n11096) );
  nnd2s1 U12085 ( .DIN1(n10491), .DIN2(n11982), .Q(n11977) );
  nnd2s1 U12086 ( .DIN1(n10492), .DIN2(n11969), .Q(n11976) );
  nnd2s1 U12087 ( .DIN1(n11133), .DIN2(n10510), .Q(n11969) );
  or3s1 U12088 ( .DIN1(n11983), .DIN2(n11984), .DIN3(n11985), .Q(n5424) );
  nnd4s1 U12089 ( .DIN1(n11986), .DIN2(n11987), .DIN3(n11988), .DIN4(n11989), 
        .Q(n11985) );
  and3s1 U12090 ( .DIN1(n11990), .DIN2(n11991), .DIN3(n11992), .Q(n11989) );
  nnd2s1 U12091 ( .DIN1(n10893), .DIN2(n10878), .Q(n11991) );
  nnd2s1 U12092 ( .DIN1(n11242), .DIN2(n10879), .Q(n11990) );
  nnd3s1 U12093 ( .DIN1(n11993), .DIN2(n11994), .DIN3(n11995), .Q(n11984) );
  nnd2s1 U12094 ( .DIN1(n10877), .DIN2(n10662), .Q(n11995) );
  or2s1 U12095 ( .DIN1(n11180), .DIN2(n11996), .Q(n11994) );
  nnd2s1 U12096 ( .DIN1(n11198), .DIN2(n10910), .Q(n11993) );
  nnd4s1 U12097 ( .DIN1(n11997), .DIN2(n11998), .DIN3(n11999), .DIN4(n12000), 
        .Q(n11983) );
  nnd2s1 U12098 ( .DIN1(n11710), .DIN2(n12001), .Q(n12000) );
  nnd2s1 U12099 ( .DIN1(n11747), .DIN2(n11215), .Q(n12001) );
  nnd2s1 U12100 ( .DIN1(n10663), .DIN2(n12002), .Q(n11999) );
  nnd2s1 U12101 ( .DIN1(n11182), .DIN2(n10680), .Q(n12002) );
  nor2s1 U12102 ( .DIN1(n11174), .DIN2(n11705), .Q(n11182) );
  nnd2s1 U12103 ( .DIN1(n10685), .DIN2(n12003), .Q(n11998) );
  nnd2s1 U12104 ( .DIN1(n10867), .DIN2(n12004), .Q(n11997) );
  hi1s1 U12105 ( .DIN(n11937), .Q(n11938) );
  xor2s1 U12106 ( .DIN1(n5047), .DIN2(n12005), .Q(n11937) );
  xnr2s1 U12107 ( .DIN1(n5023), .DIN2(w1[2]), .Q(n12005) );
  or3s1 U12108 ( .DIN1(n12006), .DIN2(n12007), .DIN3(n12008), .Q(n5023) );
  nnd4s1 U12109 ( .DIN1(n11006), .DIN2(n12009), .DIN3(n12010), .DIN4(n12011), 
        .Q(n12008) );
  and4s1 U12110 ( .DIN1(n12012), .DIN2(n12013), .DIN3(n12014), .DIN4(n12015), 
        .Q(n12011) );
  nnd2s1 U12111 ( .DIN1(n10546), .DIN2(n12016), .Q(n12015) );
  nnd2s1 U12112 ( .DIN1(n10957), .DIN2(n10548), .Q(n12016) );
  nnd2s1 U12113 ( .DIN1(n10937), .DIN2(n12017), .Q(n12014) );
  nnd2s1 U12114 ( .DIN1(n10933), .DIN2(n10964), .Q(n12017) );
  nnd2s1 U12115 ( .DIN1(n10702), .DIN2(n12018), .Q(n12013) );
  nnd3s1 U12116 ( .DIN1(n10739), .DIN2(n10940), .DIN3(n10538), .Q(n12018) );
  nnd2s1 U12117 ( .DIN1(n10550), .DIN2(n12019), .Q(n12012) );
  nnd2s1 U12118 ( .DIN1(n10729), .DIN2(n10951), .Q(n12010) );
  nnd2s1 U12119 ( .DIN1(n10703), .DIN2(n10743), .Q(n12009) );
  nnd2s1 U12120 ( .DIN1(n10717), .DIN2(n10758), .Q(n11006) );
  nnd3s1 U12121 ( .DIN1(n12020), .DIN2(n12021), .DIN3(n11769), .Q(n12007) );
  nor4s1 U12122 ( .DIN1(n12022), .DIN2(n12023), .DIN3(n12024), .DIN4(n12025), 
        .Q(n11769) );
  nnd4s1 U12123 ( .DIN1(n12026), .DIN2(n12027), .DIN3(n11352), .DIN4(n12028), 
        .Q(n12025) );
  nnd2s1 U12124 ( .DIN1(n10758), .DIN2(n11347), .Q(n12028) );
  nnd2s1 U12125 ( .DIN1(n10732), .DIN2(n11329), .Q(n11352) );
  nnd2s1 U12126 ( .DIN1(n10744), .DIN2(n10743), .Q(n12027) );
  nnd2s1 U12127 ( .DIN1(n10546), .DIN2(n11379), .Q(n12026) );
  nnd3s1 U12128 ( .DIN1(n12029), .DIN2(n12030), .DIN3(n12031), .Q(n12024) );
  nnd2s1 U12129 ( .DIN1(n10934), .DIN2(n12032), .Q(n12031) );
  nnd2s1 U12130 ( .DIN1(n10548), .DIN2(n10558), .Q(n12032) );
  nnd2s1 U12131 ( .DIN1(n10714), .DIN2(n12033), .Q(n12030) );
  nnd2s1 U12132 ( .DIN1(n10957), .DIN2(n10961), .Q(n12033) );
  nnd2s1 U12133 ( .DIN1(n10722), .DIN2(n12034), .Q(n12029) );
  nnd2s1 U12134 ( .DIN1(n10538), .DIN2(n11270), .Q(n12034) );
  nor2s1 U12135 ( .DIN1(n10752), .DIN2(n10743), .Q(n10538) );
  nor2s1 U12136 ( .DIN1(n11262), .DIN2(n10734), .Q(n12023) );
  nor2s1 U12137 ( .DIN1(n10749), .DIN2(n10743), .Q(n11262) );
  nor2s1 U12138 ( .DIN1(n12035), .DIN2(n10712), .Q(n12022) );
  nor2s1 U12139 ( .DIN1(n10716), .DIN2(n10550), .Q(n12035) );
  nnd4s1 U12140 ( .DIN1(n12036), .DIN2(n12037), .DIN3(n12038), .DIN4(n12039), 
        .Q(n12006) );
  nnd2s1 U12141 ( .DIN1(n11379), .DIN2(n10716), .Q(n12039) );
  nnd2s1 U12142 ( .DIN1(n10996), .DIN2(n10541), .Q(n12038) );
  nnd2s1 U12143 ( .DIN1(n10732), .DIN2(n10952), .Q(n12037) );
  or3s1 U12144 ( .DIN1(n12040), .DIN2(n12041), .DIN3(n12042), .Q(n5047) );
  nnd4s1 U12145 ( .DIN1(n12043), .DIN2(n12044), .DIN3(n10564), .DIN4(n12045), 
        .Q(n12042) );
  and3s1 U12146 ( .DIN1(n12046), .DIN2(n12047), .DIN3(n12048), .Q(n12045) );
  nnd2s1 U12147 ( .DIN1(n10592), .DIN2(n10583), .Q(n12047) );
  nnd2s1 U12148 ( .DIN1(n10588), .DIN2(n11030), .Q(n12046) );
  nor3s1 U12149 ( .DIN1(n12049), .DIN2(n12050), .DIN3(n12051), .Q(n10564) );
  nnd4s1 U12150 ( .DIN1(n12052), .DIN2(n12053), .DIN3(n12054), .DIN4(n12055), 
        .Q(n12051) );
  and3s1 U12151 ( .DIN1(n12056), .DIN2(n12057), .DIN3(n12058), .Q(n12055) );
  nnd2s1 U12152 ( .DIN1(n10782), .DIN2(n10573), .Q(n12058) );
  nnd2s1 U12153 ( .DIN1(n11018), .DIN2(n10578), .Q(n12057) );
  nnd2s1 U12154 ( .DIN1(n10592), .DIN2(n11029), .Q(n12056) );
  nnd3s1 U12155 ( .DIN1(n12059), .DIN2(n12060), .DIN3(n11894), .Q(n12050) );
  nnd2s1 U12156 ( .DIN1(n11020), .DIN2(n11870), .Q(n11894) );
  or2s1 U12157 ( .DIN1(n10598), .DIN2(n11902), .Q(n12060) );
  nor2s1 U12158 ( .DIN1(n10570), .DIN2(n10581), .Q(n11902) );
  nnd2s1 U12159 ( .DIN1(n11053), .DIN2(n10793), .Q(n12059) );
  nnd2s1 U12160 ( .DIN1(n11044), .DIN2(n10784), .Q(n10793) );
  nnd4s1 U12161 ( .DIN1(n12061), .DIN2(n12062), .DIN3(n12063), .DIN4(n12064), 
        .Q(n12049) );
  nnd2s1 U12162 ( .DIN1(n11404), .DIN2(n12065), .Q(n12064) );
  nnd2s1 U12163 ( .DIN1(n10572), .DIN2(n12066), .Q(n12063) );
  nnd2s1 U12164 ( .DIN1(n10784), .DIN2(n11059), .Q(n12066) );
  nnd2s1 U12165 ( .DIN1(n11019), .DIN2(n12067), .Q(n12062) );
  nnd2s1 U12166 ( .DIN1(n11042), .DIN2(n10591), .Q(n12067) );
  nnd2s1 U12167 ( .DIN1(n10596), .DIN2(n12068), .Q(n12061) );
  nnd2s1 U12168 ( .DIN1(n11910), .DIN2(n11804), .Q(n12068) );
  hi1s1 U12169 ( .DIN(n11052), .Q(n11910) );
  nnd2s1 U12170 ( .DIN1(n11444), .DIN2(n11063), .Q(n11052) );
  nnd3s1 U12171 ( .DIN1(n12069), .DIN2(n12070), .DIN3(n12071), .Q(n12041) );
  nnd2s1 U12172 ( .DIN1(n11018), .DIN2(n10580), .Q(n12071) );
  or2s1 U12173 ( .DIN1(n10594), .DIN2(n10590), .Q(n12070) );
  nor2s1 U12174 ( .DIN1(n10782), .DIN2(n10786), .Q(n10590) );
  nnd2s1 U12175 ( .DIN1(n11427), .DIN2(n10600), .Q(n12069) );
  nnd4s1 U12176 ( .DIN1(n12072), .DIN2(n12073), .DIN3(n12074), .DIN4(n12075), 
        .Q(n12040) );
  nnd2s1 U12177 ( .DIN1(n11875), .DIN2(n12076), .Q(n12075) );
  nnd2s1 U12178 ( .DIN1(n11911), .DIN2(n11444), .Q(n12076) );
  nnd2s1 U12179 ( .DIN1(n10571), .DIN2(n12077), .Q(n12074) );
  nnd2s1 U12180 ( .DIN1(n11411), .DIN2(n10785), .Q(n12077) );
  nor2s1 U12181 ( .DIN1(n10579), .DIN2(n11870), .Q(n11411) );
  nnd2s1 U12182 ( .DIN1(n10572), .DIN2(n12078), .Q(n12073) );
  nnd2s1 U12183 ( .DIN1(n10573), .DIN2(n12065), .Q(n12072) );
  nnd2s1 U12184 ( .DIN1(n11448), .DIN2(n10591), .Q(n12065) );
  hi1s1 U12185 ( .DIN(n5423), .Q(n11939) );
  nnd2s1 U12186 ( .DIN1(n12079), .DIN2(n12080), .Q(N163) );
  nnd2s1 U12187 ( .DIN1(n12081), .DIN2(n1631), .Q(n12080) );
  xor2s1 U12188 ( .DIN1(n12082), .DIN2(n12083), .Q(n12081) );
  xor2s1 U12189 ( .DIN1(n11477), .DIN2(n12084), .Q(n12083) );
  xor2s1 U12190 ( .DIN1(n12085), .DIN2(n10300), .Q(n12084) );
  xor2s1 U12191 ( .DIN1(n5423), .DIN2(n5070), .Q(n10300) );
  or3s1 U12192 ( .DIN1(n12086), .DIN2(n12087), .DIN3(n12088), .Q(n5070) );
  nnd4s1 U12193 ( .DIN1(n12089), .DIN2(n11078), .DIN3(n12090), .DIN4(n12091), 
        .Q(n12088) );
  and3s1 U12194 ( .DIN1(n10481), .DIN2(n11958), .DIN3(n11947), .Q(n12091) );
  nor4s1 U12195 ( .DIN1(n12092), .DIN2(n12093), .DIN3(n12094), .DIN4(n12095), 
        .Q(n11947) );
  nnd4s1 U12196 ( .DIN1(n12096), .DIN2(n11584), .DIN3(n12097), .DIN4(n12098), 
        .Q(n12095) );
  nnd2s1 U12197 ( .DIN1(n10840), .DIN2(n10520), .Q(n12098) );
  nnd2s1 U12198 ( .DIN1(n10492), .DIN2(n10843), .Q(n12097) );
  nnd2s1 U12199 ( .DIN1(n10501), .DIN2(n11567), .Q(n11584) );
  nnd2s1 U12200 ( .DIN1(n10639), .DIN2(n11089), .Q(n12096) );
  nnd3s1 U12201 ( .DIN1(n12099), .DIN2(n12100), .DIN3(n12101), .Q(n12094) );
  nnd2s1 U12202 ( .DIN1(n10507), .DIN2(n12102), .Q(n12101) );
  nnd2s1 U12203 ( .DIN1(n10497), .DIN2(n12103), .Q(n12100) );
  nnd2s1 U12204 ( .DIN1(n10645), .DIN2(n10642), .Q(n12103) );
  nnd2s1 U12205 ( .DIN1(n10628), .DIN2(n12104), .Q(n12099) );
  nnd2s1 U12206 ( .DIN1(n10633), .DIN2(n10517), .Q(n12104) );
  nor2s1 U12207 ( .DIN1(n11503), .DIN2(n10826), .Q(n12093) );
  nor2s1 U12208 ( .DIN1(n10850), .DIN2(n10843), .Q(n11503) );
  nor2s1 U12209 ( .DIN1(n12105), .DIN2(n11497), .Q(n12092) );
  nor2s1 U12210 ( .DIN1(n10809), .DIN2(n10808), .Q(n12105) );
  nor2s1 U12211 ( .DIN1(n12106), .DIN2(n12107), .Q(n11958) );
  nnd4s1 U12212 ( .DIN1(n12108), .DIN2(n12109), .DIN3(n11610), .DIN4(n12110), 
        .Q(n12107) );
  nnd2s1 U12213 ( .DIN1(n10628), .DIN2(n10635), .Q(n12110) );
  nnd2s1 U12214 ( .DIN1(n11155), .DIN2(n10518), .Q(n10635) );
  nnd2s1 U12215 ( .DIN1(n10639), .DIN2(n10500), .Q(n11610) );
  nnd2s1 U12216 ( .DIN1(n11113), .DIN2(n11089), .Q(n12109) );
  nnd2s1 U12217 ( .DIN1(n10492), .DIN2(n10643), .Q(n12108) );
  nnd4s1 U12218 ( .DIN1(n12111), .DIN2(n12112), .DIN3(n12113), .DIN4(n12114), 
        .Q(n12106) );
  nnd2s1 U12219 ( .DIN1(n10501), .DIN2(n12115), .Q(n12114) );
  nnd2s1 U12220 ( .DIN1(n11504), .DIN2(n11099), .Q(n12115) );
  nnd2s1 U12221 ( .DIN1(n10840), .DIN2(n12116), .Q(n12113) );
  nnd2s1 U12222 ( .DIN1(n10834), .DIN2(n10849), .Q(n12116) );
  nnd2s1 U12223 ( .DIN1(n10810), .DIN2(n12117), .Q(n12112) );
  nnd3s1 U12224 ( .DIN1(n10646), .DIN2(n10642), .DIN3(n10632), .Q(n12117) );
  nnd2s1 U12225 ( .DIN1(n10827), .DIN2(n12118), .Q(n12111) );
  nnd4s1 U12226 ( .DIN1(n10817), .DIN2(n10834), .DIN3(n11102), .DIN4(n10645), 
        .Q(n12118) );
  nor2s1 U12227 ( .DIN1(n12119), .DIN2(n12120), .Q(n10481) );
  nnd4s1 U12228 ( .DIN1(n12121), .DIN2(n12122), .DIN3(n12123), .DIN4(n12124), 
        .Q(n12120) );
  nnd2s1 U12229 ( .DIN1(n10502), .DIN2(n11121), .Q(n12124) );
  nnd2s1 U12230 ( .DIN1(n10832), .DIN2(n10517), .Q(n11121) );
  nnd2s1 U12231 ( .DIN1(n10498), .DIN2(n10499), .Q(n12123) );
  nnd2s1 U12232 ( .DIN1(n10491), .DIN2(n10809), .Q(n12122) );
  nnd2s1 U12233 ( .DIN1(n10850), .DIN2(n11112), .Q(n12121) );
  nnd4s1 U12234 ( .DIN1(n12125), .DIN2(n12126), .DIN3(n12127), .DIN4(n12128), 
        .Q(n12119) );
  nnd2s1 U12235 ( .DIN1(n10627), .DIN2(n12129), .Q(n12128) );
  or2s1 U12236 ( .DIN1(n11613), .DIN2(n10501), .Q(n12129) );
  nnd2s1 U12237 ( .DIN1(n10820), .DIN2(n12130), .Q(n12127) );
  nnd2s1 U12238 ( .DIN1(n10632), .DIN2(n10829), .Q(n12130) );
  nnd2s1 U12239 ( .DIN1(n10492), .DIN2(n12131), .Q(n12126) );
  nnd2s1 U12240 ( .DIN1(n11137), .DIN2(n10518), .Q(n12131) );
  nnd2s1 U12241 ( .DIN1(n10515), .DIN2(n12132), .Q(n12125) );
  nnd3s1 U12242 ( .DIN1(n11137), .DIN2(n11133), .DIN3(n12133), .Q(n12132) );
  nnd2s1 U12243 ( .DIN1(n10502), .DIN2(n10840), .Q(n11078) );
  nnd2s1 U12244 ( .DIN1(n11113), .DIN2(n10515), .Q(n12089) );
  nnd3s1 U12245 ( .DIN1(n12134), .DIN2(n12135), .DIN3(n12136), .Q(n12087) );
  nnd2s1 U12246 ( .DIN1(n10639), .DIN2(n10819), .Q(n12136) );
  nnd2s1 U12247 ( .DIN1(n10501), .DIN2(n10498), .Q(n12135) );
  nnd2s1 U12248 ( .DIN1(n11089), .DIN2(n10490), .Q(n12134) );
  nnd4s1 U12249 ( .DIN1(n12137), .DIN2(n12138), .DIN3(n12139), .DIN4(n12140), 
        .Q(n12086) );
  nnd2s1 U12250 ( .DIN1(n11562), .DIN2(n12141), .Q(n12140) );
  nnd2s1 U12251 ( .DIN1(n11129), .DIN2(n11098), .Q(n12141) );
  nnd2s1 U12252 ( .DIN1(n10507), .DIN2(n12142), .Q(n12139) );
  nnd2s1 U12253 ( .DIN1(n11497), .DIN2(n11133), .Q(n12142) );
  nnd2s1 U12254 ( .DIN1(n10808), .DIN2(n12143), .Q(n12138) );
  nnd2s1 U12255 ( .DIN1(n10818), .DIN2(n11155), .Q(n12143) );
  nor2s1 U12256 ( .DIN1(n10491), .DIN2(n10843), .Q(n10818) );
  nnd2s1 U12257 ( .DIN1(n10809), .DIN2(n12144), .Q(n12137) );
  nnd3s1 U12258 ( .DIN1(n11132), .DIN2(n11130), .DIN3(n10633), .Q(n12144) );
  nor2s1 U12259 ( .DIN1(n10519), .DIN2(n10843), .Q(n10633) );
  or3s1 U12260 ( .DIN1(n12145), .DIN2(n12146), .DIN3(n12147), .Q(n5423) );
  nnd4s1 U12261 ( .DIN1(n12148), .DIN2(n11161), .DIN3(n12149), .DIN4(n12150), 
        .Q(n12147) );
  and3s1 U12262 ( .DIN1(n12151), .DIN2(n12152), .DIN3(n11986), .Q(n12150) );
  nor4s1 U12263 ( .DIN1(n12153), .DIN2(n12154), .DIN3(n12155), .DIN4(n12156), 
        .Q(n11986) );
  nnd4s1 U12264 ( .DIN1(n12157), .DIN2(n11728), .DIN3(n12158), .DIN4(n12159), 
        .Q(n12156) );
  nnd2s1 U12265 ( .DIN1(n10901), .DIN2(n11725), .Q(n12159) );
  nnd2s1 U12266 ( .DIN1(n10867), .DIN2(n10905), .Q(n12158) );
  nnd2s1 U12267 ( .DIN1(n10884), .DIN2(n11710), .Q(n11728) );
  nnd2s1 U12268 ( .DIN1(n10677), .DIN2(n11173), .Q(n12157) );
  nnd3s1 U12269 ( .DIN1(n12160), .DIN2(n12161), .DIN3(n12162), .Q(n12155) );
  nnd2s1 U12270 ( .DIN1(n11242), .DIN2(n12163), .Q(n12162) );
  nnd2s1 U12271 ( .DIN1(n11172), .DIN2(n12164), .Q(n12161) );
  nnd2s1 U12272 ( .DIN1(n10683), .DIN2(n10680), .Q(n12164) );
  nnd2s1 U12273 ( .DIN1(n10664), .DIN2(n12165), .Q(n12160) );
  nnd2s1 U12274 ( .DIN1(n10669), .DIN2(n11704), .Q(n12165) );
  nor2s1 U12275 ( .DIN1(n11645), .DIN2(n10886), .Q(n12154) );
  nor2s1 U12276 ( .DIN1(n10913), .DIN2(n10905), .Q(n11645) );
  nor2s1 U12277 ( .DIN1(n12166), .DIN2(n11638), .Q(n12153) );
  nor2s1 U12278 ( .DIN1(n10865), .DIN2(n10877), .Q(n12166) );
  nnd2s1 U12279 ( .DIN1(n10878), .DIN2(n10901), .Q(n11161) );
  nnd2s1 U12280 ( .DIN1(n11199), .DIN2(n10672), .Q(n12148) );
  nnd3s1 U12281 ( .DIN1(n12167), .DIN2(n12168), .DIN3(n12169), .Q(n12146) );
  nnd2s1 U12282 ( .DIN1(n10677), .DIN2(n10876), .Q(n12169) );
  nnd2s1 U12283 ( .DIN1(n10884), .DIN2(n11174), .Q(n12168) );
  nnd2s1 U12284 ( .DIN1(n11173), .DIN2(n10663), .Q(n12167) );
  nnd4s1 U12285 ( .DIN1(n12170), .DIN2(n12171), .DIN3(n12172), .DIN4(n12173), 
        .Q(n12145) );
  nnd2s1 U12286 ( .DIN1(n11705), .DIN2(n12174), .Q(n12173) );
  nnd2s1 U12287 ( .DIN1(n11215), .DIN2(n11184), .Q(n12174) );
  nnd2s1 U12288 ( .DIN1(n11242), .DIN2(n12175), .Q(n12172) );
  nnd2s1 U12289 ( .DIN1(n11638), .DIN2(n11219), .Q(n12175) );
  nnd2s1 U12290 ( .DIN1(n10877), .DIN2(n12176), .Q(n12171) );
  nnd2s1 U12291 ( .DIN1(n10875), .DIN2(n11244), .Q(n12176) );
  nor2s1 U12292 ( .DIN1(n10685), .DIN2(n10905), .Q(n10875) );
  nnd2s1 U12293 ( .DIN1(n10865), .DIN2(n12177), .Q(n12170) );
  nnd3s1 U12294 ( .DIN1(n11218), .DIN2(n11216), .DIN3(n10669), .Q(n12177) );
  nor2s1 U12295 ( .DIN1(n10910), .DIN2(n10905), .Q(n10669) );
  xor2s1 U12296 ( .DIN1(n5046), .DIN2(n12178), .Q(n12082) );
  xor2s1 U12297 ( .DIN1(w1[1]), .DIN2(n5022), .Q(n12178) );
  nor4s1 U12298 ( .DIN1(n12179), .DIN2(n12180), .DIN3(n12181), .DIN4(n12182), 
        .Q(n5022) );
  nnd4s1 U12299 ( .DIN1(n11331), .DIN2(n11007), .DIN3(n12183), .DIN4(n12184), 
        .Q(n12182) );
  nnd2s1 U12300 ( .DIN1(n10702), .DIN2(n11380), .Q(n12184) );
  nnd2s1 U12301 ( .DIN1(n10749), .DIN2(n11347), .Q(n12183) );
  nnd2s1 U12302 ( .DIN1(n10743), .DIN2(n11264), .Q(n11007) );
  nnd2s1 U12303 ( .DIN1(n10714), .DIN2(n10541), .Q(n11331) );
  nnd4s1 U12304 ( .DIN1(n12185), .DIN2(n12186), .DIN3(n12187), .DIN4(n12188), 
        .Q(n12181) );
  nnd2s1 U12305 ( .DIN1(n10550), .DIN2(n12189), .Q(n12188) );
  nnd2s1 U12306 ( .DIN1(n10548), .DIN2(n10958), .Q(n12189) );
  nnd2s1 U12307 ( .DIN1(n10703), .DIN2(n12190), .Q(n12187) );
  nnd2s1 U12308 ( .DIN1(n10932), .DIN2(n10998), .Q(n12190) );
  nnd2s1 U12309 ( .DIN1(n10996), .DIN2(n10759), .Q(n12186) );
  nnd2s1 U12310 ( .DIN1(n10734), .DIN2(n10549), .Q(n10759) );
  or2s1 U12311 ( .DIN1(n10754), .DIN2(n10727), .Q(n12185) );
  nor2s1 U12312 ( .DIN1(n10710), .DIN2(n10701), .Q(n10727) );
  nnd3s1 U12313 ( .DIN1(n11770), .DIN2(n12191), .DIN3(n12192), .Q(n12180) );
  nor4s1 U12314 ( .DIN1(n12193), .DIN2(n12194), .DIN3(n12195), .DIN4(n12196), 
        .Q(n11770) );
  nnd4s1 U12315 ( .DIN1(n12197), .DIN2(n12198), .DIN3(n12199), .DIN4(n12200), 
        .Q(n12196) );
  nor2s1 U12316 ( .DIN1(n12201), .DIN2(n12202), .Q(n12200) );
  nor2s1 U12317 ( .DIN1(n10739), .DIN2(n10557), .Q(n12202) );
  nor2s1 U12318 ( .DIN1(n10731), .DIN2(n10932), .Q(n12201) );
  nnd2s1 U12319 ( .DIN1(n10742), .DIN2(n10934), .Q(n12199) );
  or2s1 U12320 ( .DIN1(n10725), .DIN2(n10960), .Q(n12198) );
  nor2s1 U12321 ( .DIN1(n10541), .DIN2(n11379), .Q(n10960) );
  nnd2s1 U12322 ( .DIN1(n11329), .DIN2(n10701), .Q(n12197) );
  nnd3s1 U12323 ( .DIN1(n12203), .DIN2(n12204), .DIN3(n12205), .Q(n12195) );
  nnd2s1 U12324 ( .DIN1(n10952), .DIN2(n12206), .Q(n12205) );
  nnd2s1 U12325 ( .DIN1(n10724), .DIN2(n10964), .Q(n12206) );
  nnd2s1 U12326 ( .DIN1(n10716), .DIN2(n10936), .Q(n12204) );
  nnd2s1 U12327 ( .DIN1(n10966), .DIN2(n10549), .Q(n10936) );
  nnd2s1 U12328 ( .DIN1(n10722), .DIN2(n12207), .Q(n12203) );
  nnd2s1 U12329 ( .DIN1(n10728), .DIN2(n11266), .Q(n12207) );
  nor2s1 U12330 ( .DIN1(n12208), .DIN2(n10537), .Q(n12194) );
  nor2s1 U12331 ( .DIN1(n10934), .DIN2(n10546), .Q(n12208) );
  nor2s1 U12332 ( .DIN1(n12209), .DIN2(n10548), .Q(n12193) );
  nor2s1 U12333 ( .DIN1(n10743), .DIN2(n10732), .Q(n12209) );
  nnd4s1 U12334 ( .DIN1(n12036), .DIN2(n12210), .DIN3(n12211), .DIN4(n12212), 
        .Q(n12179) );
  nnd2s1 U12335 ( .DIN1(n10742), .DIN2(n10729), .Q(n12212) );
  nnd2s1 U12336 ( .DIN1(n10990), .DIN2(n10758), .Q(n12211) );
  nnd2s1 U12337 ( .DIN1(n10951), .DIN2(n10701), .Q(n12210) );
  nor3s1 U12338 ( .DIN1(n12213), .DIN2(n12214), .DIN3(n12215), .Q(n12036) );
  nnd4s1 U12339 ( .DIN1(n12216), .DIN2(n12217), .DIN3(n11775), .DIN4(n12218), 
        .Q(n12215) );
  and3s1 U12340 ( .DIN1(n12219), .DIN2(n12220), .DIN3(n12221), .Q(n12218) );
  nnd2s1 U12341 ( .DIN1(n10546), .DIN2(n10952), .Q(n12221) );
  nnd2s1 U12342 ( .DIN1(n10996), .DIN2(n10937), .Q(n12220) );
  nnd2s1 U12343 ( .DIN1(n10744), .DIN2(n10729), .Q(n12219) );
  nor2s1 U12344 ( .DIN1(n12222), .DIN2(n12223), .Q(n11775) );
  nnd4s1 U12345 ( .DIN1(n12224), .DIN2(n12225), .DIN3(n12226), .DIN4(n12227), 
        .Q(n12223) );
  nnd2s1 U12346 ( .DIN1(n10546), .DIN2(n12228), .Q(n12227) );
  nnd2s1 U12347 ( .DIN1(n11271), .DIN2(n10558), .Q(n12228) );
  nnd2s1 U12348 ( .DIN1(n10701), .DIN2(n12229), .Q(n12226) );
  nnd3s1 U12349 ( .DIN1(n10539), .DIN2(n10548), .DIN3(n10557), .Q(n12229) );
  nnd2s1 U12350 ( .DIN1(n10714), .DIN2(n10742), .Q(n12225) );
  nnd2s1 U12351 ( .DIN1(n10703), .DIN2(n10996), .Q(n12224) );
  nnd4s1 U12352 ( .DIN1(n12230), .DIN2(n12231), .DIN3(n12232), .DIN4(n12233), 
        .Q(n12222) );
  nnd2s1 U12353 ( .DIN1(n11329), .DIN2(n12234), .Q(n12233) );
  nnd2s1 U12354 ( .DIN1(n11270), .DIN2(n10933), .Q(n12234) );
  nnd2s1 U12355 ( .DIN1(n10717), .DIN2(n12235), .Q(n12232) );
  nnd2s1 U12356 ( .DIN1(n10724), .DIN2(n10757), .Q(n12235) );
  nnd2s1 U12357 ( .DIN1(n10533), .DIN2(n12236), .Q(n12231) );
  nnd2s1 U12358 ( .DIN1(n11307), .DIN2(n10712), .Q(n12236) );
  nor2s1 U12359 ( .DIN1(n11379), .DIN2(n10990), .Q(n11307) );
  nnd2s1 U12360 ( .DIN1(n10732), .DIN2(n12237), .Q(n12230) );
  nnd2s1 U12361 ( .DIN1(n10558), .DIN2(n10958), .Q(n12237) );
  nnd3s1 U12362 ( .DIN1(n12238), .DIN2(n12239), .DIN3(n12240), .Q(n12214) );
  nnd2s1 U12363 ( .DIN1(n10703), .DIN2(n10758), .Q(n12240) );
  nnd2s1 U12364 ( .DIN1(n10934), .DIN2(n11329), .Q(n12239) );
  nnd2s1 U12365 ( .DIN1(n10714), .DIN2(n10722), .Q(n12238) );
  nnd4s1 U12366 ( .DIN1(n12241), .DIN2(n12242), .DIN3(n12243), .DIN4(n12244), 
        .Q(n12213) );
  nnd2s1 U12367 ( .DIN1(n10951), .DIN2(n12245), .Q(n12244) );
  nnd2s1 U12368 ( .DIN1(n11270), .DIN2(n10998), .Q(n12245) );
  nnd2s1 U12369 ( .DIN1(n10990), .DIN2(n12246), .Q(n12243) );
  nnd4s1 U12370 ( .DIN1(n10998), .DIN2(n10725), .DIN3(n10964), .DIN4(n10940), 
        .Q(n12246) );
  nnd2s1 U12371 ( .DIN1(n10749), .DIN2(n11304), .Q(n12242) );
  nnd2s1 U12372 ( .DIN1(n10957), .DIN2(n10539), .Q(n11304) );
  nnd2s1 U12373 ( .DIN1(n10533), .DIN2(n10941), .Q(n12241) );
  nnd2s1 U12374 ( .DIN1(n10537), .DIN2(n10549), .Q(n10941) );
  or3s1 U12375 ( .DIN1(n12247), .DIN2(n12248), .DIN3(n12249), .Q(n5046) );
  nnd4s1 U12376 ( .DIN1(n12250), .DIN2(n11393), .DIN3(n12251), .DIN4(n12252), 
        .Q(n12249) );
  and3s1 U12377 ( .DIN1(n10562), .DIN2(n12054), .DIN3(n12043), .Q(n12252) );
  nor4s1 U12378 ( .DIN1(n12253), .DIN2(n12254), .DIN3(n12255), .DIN4(n12256), 
        .Q(n12043) );
  nnd4s1 U12379 ( .DIN1(n12257), .DIN2(n11892), .DIN3(n12258), .DIN4(n12259), 
        .Q(n12256) );
  nnd2s1 U12380 ( .DIN1(n11050), .DIN2(n10601), .Q(n12259) );
  nnd2s1 U12381 ( .DIN1(n10573), .DIN2(n11053), .Q(n12258) );
  nnd2s1 U12382 ( .DIN1(n10582), .DIN2(n11875), .Q(n11892) );
  nnd2s1 U12383 ( .DIN1(n10782), .DIN2(n11404), .Q(n12257) );
  nnd3s1 U12384 ( .DIN1(n12260), .DIN2(n12261), .DIN3(n12262), .Q(n12255) );
  nnd2s1 U12385 ( .DIN1(n10588), .DIN2(n12263), .Q(n12262) );
  nnd2s1 U12386 ( .DIN1(n10578), .DIN2(n12264), .Q(n12261) );
  nnd2s1 U12387 ( .DIN1(n10788), .DIN2(n10785), .Q(n12264) );
  nnd2s1 U12388 ( .DIN1(n10771), .DIN2(n12265), .Q(n12260) );
  nnd2s1 U12389 ( .DIN1(n10776), .DIN2(n10598), .Q(n12265) );
  nor2s1 U12390 ( .DIN1(n11811), .DIN2(n11036), .Q(n12254) );
  nor2s1 U12391 ( .DIN1(n11060), .DIN2(n11053), .Q(n11811) );
  nor2s1 U12392 ( .DIN1(n12266), .DIN2(n11805), .Q(n12253) );
  nor2s1 U12393 ( .DIN1(n11019), .DIN2(n11018), .Q(n12266) );
  nor2s1 U12394 ( .DIN1(n12267), .DIN2(n12268), .Q(n12054) );
  nnd4s1 U12395 ( .DIN1(n12269), .DIN2(n12270), .DIN3(n11918), .DIN4(n12271), 
        .Q(n12268) );
  nnd2s1 U12396 ( .DIN1(n10771), .DIN2(n10778), .Q(n12271) );
  nnd2s1 U12397 ( .DIN1(n11470), .DIN2(n10599), .Q(n10778) );
  nnd2s1 U12398 ( .DIN1(n10782), .DIN2(n10581), .Q(n11918) );
  nnd2s1 U12399 ( .DIN1(n11428), .DIN2(n11404), .Q(n12270) );
  nnd2s1 U12400 ( .DIN1(n10573), .DIN2(n10786), .Q(n12269) );
  nnd4s1 U12401 ( .DIN1(n12272), .DIN2(n12273), .DIN3(n12274), .DIN4(n12275), 
        .Q(n12267) );
  nnd2s1 U12402 ( .DIN1(n10582), .DIN2(n12276), .Q(n12275) );
  nnd2s1 U12403 ( .DIN1(n11812), .DIN2(n11414), .Q(n12276) );
  nnd2s1 U12404 ( .DIN1(n11050), .DIN2(n12277), .Q(n12274) );
  nnd2s1 U12405 ( .DIN1(n11044), .DIN2(n11059), .Q(n12277) );
  nnd2s1 U12406 ( .DIN1(n11020), .DIN2(n12278), .Q(n12273) );
  nnd3s1 U12407 ( .DIN1(n10789), .DIN2(n10785), .DIN3(n10775), .Q(n12278) );
  nnd2s1 U12408 ( .DIN1(n11037), .DIN2(n12279), .Q(n12272) );
  nnd4s1 U12409 ( .DIN1(n11027), .DIN2(n11044), .DIN3(n11417), .DIN4(n10788), 
        .Q(n12279) );
  nor2s1 U12410 ( .DIN1(n12280), .DIN2(n12281), .Q(n10562) );
  nnd4s1 U12411 ( .DIN1(n12282), .DIN2(n12283), .DIN3(n12284), .DIN4(n12285), 
        .Q(n12281) );
  nnd2s1 U12412 ( .DIN1(n10583), .DIN2(n11436), .Q(n12285) );
  nnd2s1 U12413 ( .DIN1(n11042), .DIN2(n10598), .Q(n11436) );
  nnd2s1 U12414 ( .DIN1(n10579), .DIN2(n10580), .Q(n12284) );
  nnd2s1 U12415 ( .DIN1(n10572), .DIN2(n11019), .Q(n12283) );
  nnd2s1 U12416 ( .DIN1(n11060), .DIN2(n11427), .Q(n12282) );
  nnd4s1 U12417 ( .DIN1(n12286), .DIN2(n12287), .DIN3(n12288), .DIN4(n12289), 
        .Q(n12280) );
  nnd2s1 U12418 ( .DIN1(n10770), .DIN2(n12290), .Q(n12289) );
  or2s1 U12419 ( .DIN1(n11921), .DIN2(n10582), .Q(n12290) );
  nnd2s1 U12420 ( .DIN1(n11030), .DIN2(n12291), .Q(n12288) );
  nnd2s1 U12421 ( .DIN1(n10775), .DIN2(n11039), .Q(n12291) );
  nnd2s1 U12422 ( .DIN1(n10573), .DIN2(n12292), .Q(n12287) );
  nnd2s1 U12423 ( .DIN1(n11452), .DIN2(n10599), .Q(n12292) );
  nnd2s1 U12424 ( .DIN1(n10596), .DIN2(n12293), .Q(n12286) );
  nnd3s1 U12425 ( .DIN1(n11452), .DIN2(n11448), .DIN3(n12294), .Q(n12293) );
  nnd2s1 U12426 ( .DIN1(n10583), .DIN2(n11050), .Q(n11393) );
  nnd2s1 U12427 ( .DIN1(n11428), .DIN2(n10596), .Q(n12250) );
  nnd3s1 U12428 ( .DIN1(n12295), .DIN2(n12296), .DIN3(n12297), .Q(n12248) );
  nnd2s1 U12429 ( .DIN1(n10782), .DIN2(n11029), .Q(n12297) );
  nnd2s1 U12430 ( .DIN1(n10582), .DIN2(n10579), .Q(n12296) );
  nnd2s1 U12431 ( .DIN1(n11404), .DIN2(n10571), .Q(n12295) );
  nnd4s1 U12432 ( .DIN1(n12298), .DIN2(n12299), .DIN3(n12300), .DIN4(n12301), 
        .Q(n12247) );
  nnd2s1 U12433 ( .DIN1(n11870), .DIN2(n12302), .Q(n12301) );
  nnd2s1 U12434 ( .DIN1(n11444), .DIN2(n11413), .Q(n12302) );
  nnd2s1 U12435 ( .DIN1(n10588), .DIN2(n12303), .Q(n12300) );
  nnd2s1 U12436 ( .DIN1(n11805), .DIN2(n11448), .Q(n12303) );
  nnd2s1 U12437 ( .DIN1(n11018), .DIN2(n12304), .Q(n12299) );
  nnd2s1 U12438 ( .DIN1(n11028), .DIN2(n11470), .Q(n12304) );
  nor2s1 U12439 ( .DIN1(n10572), .DIN2(n11053), .Q(n11028) );
  nnd2s1 U12440 ( .DIN1(n11019), .DIN2(n12305), .Q(n12298) );
  nnd3s1 U12441 ( .DIN1(n11447), .DIN2(n11445), .DIN3(n10776), .Q(n12305) );
  nor2s1 U12442 ( .DIN1(n10600), .DIN2(n11053), .Q(n10776) );
  nnd2s1 U12443 ( .DIN1(n12306), .DIN2(n1602), .Q(n12079) );
  xor2s1 U12444 ( .DIN1(w1[1]), .DIN2(text_in_r[65]), .Q(n12306) );
  nnd2s1 U12445 ( .DIN1(n12307), .DIN2(n12308), .Q(N162) );
  nnd2s1 U12446 ( .DIN1(n12309), .DIN2(n1633), .Q(n12308) );
  xor2s1 U12447 ( .DIN1(n12310), .DIN2(n12311), .Q(n12309) );
  xor2s1 U12448 ( .DIN1(n10308), .DIN2(n11071), .Q(n12311) );
  hi1s1 U12449 ( .DIN(n11477), .Q(n11071) );
  xor2s1 U12450 ( .DIN1(n5701), .DIN2(n5029), .Q(n11477) );
  nor3s1 U12451 ( .DIN1(n12312), .DIN2(n12313), .DIN3(n12314), .Q(n5029) );
  nnd4s1 U12452 ( .DIN1(n12020), .DIN2(n12192), .DIN3(n11771), .DIN4(n12315), 
        .Q(n12314) );
  and4s1 U12453 ( .DIN1(n12216), .DIN2(n12316), .DIN3(n12317), .DIN4(n10975), 
        .Q(n12315) );
  nnd2s1 U12454 ( .DIN1(n10729), .DIN2(n10715), .Q(n10975) );
  nnd2s1 U12455 ( .DIN1(n10732), .DIN2(n10717), .Q(n12317) );
  nnd2s1 U12456 ( .DIN1(n10533), .DIN2(n11264), .Q(n12316) );
  and4s1 U12457 ( .DIN1(n12318), .DIN2(n12319), .DIN3(n12320), .DIN4(n12321), 
        .Q(n12216) );
  and4s1 U12458 ( .DIN1(n12322), .DIN2(n12323), .DIN3(n12324), .DIN4(n12325), 
        .Q(n12321) );
  nnd2s1 U12459 ( .DIN1(n10742), .DIN2(n10533), .Q(n12325) );
  nnd2s1 U12460 ( .DIN1(n10532), .DIN2(n10752), .Q(n12324) );
  nnd2s1 U12461 ( .DIN1(n10550), .DIN2(n11264), .Q(n12323) );
  nnd2s1 U12462 ( .DIN1(n10934), .DIN2(n10937), .Q(n12322) );
  and3s1 U12463 ( .DIN1(n12326), .DIN2(n12327), .DIN3(n12328), .Q(n12320) );
  nnd2s1 U12464 ( .DIN1(n10703), .DIN2(n12329), .Q(n12328) );
  nnd3s1 U12465 ( .DIN1(n12330), .DIN2(n10940), .DIN3(n10757), .Q(n12329) );
  nnd2s1 U12466 ( .DIN1(n10758), .DIN2(n11323), .Q(n12327) );
  nnd2s1 U12467 ( .DIN1(n10961), .DIN2(n10751), .Q(n11323) );
  nnd2s1 U12468 ( .DIN1(n10717), .DIN2(n12331), .Q(n12326) );
  nnd2s1 U12469 ( .DIN1(n10932), .DIN2(n10725), .Q(n12331) );
  nnd2s1 U12470 ( .DIN1(n10996), .DIN2(n12332), .Q(n12319) );
  nnd4s1 U12471 ( .DIN1(n10557), .DIN2(n10548), .DIN3(n10558), .DIN4(n10754), 
        .Q(n12332) );
  nnd2s1 U12472 ( .DIN1(n10743), .DIN2(n10952), .Q(n12318) );
  nor3s1 U12473 ( .DIN1(n12333), .DIN2(n12334), .DIN3(n12335), .Q(n11771) );
  nnd4s1 U12474 ( .DIN1(n12191), .DIN2(n12217), .DIN3(n12021), .DIN4(n12336), 
        .Q(n12335) );
  and4s1 U12475 ( .DIN1(n12337), .DIN2(n12338), .DIN3(n12339), .DIN4(n12340), 
        .Q(n12336) );
  nnd2s1 U12476 ( .DIN1(n10749), .DIN2(n11379), .Q(n12340) );
  nnd2s1 U12477 ( .DIN1(n10546), .DIN2(n10744), .Q(n12339) );
  nnd2s1 U12478 ( .DIN1(n10703), .DIN2(n10934), .Q(n12338) );
  hi1s1 U12479 ( .DIN(n10957), .Q(n10703) );
  nnd2s1 U12480 ( .DIN1(n10710), .DIN2(n10715), .Q(n12337) );
  nor2s1 U12481 ( .DIN1(n12341), .DIN2(n12342), .Q(n12021) );
  nnd4s1 U12482 ( .DIN1(n11249), .DIN2(n12343), .DIN3(n12344), .DIN4(n12345), 
        .Q(n12342) );
  nnd2s1 U12483 ( .DIN1(n10732), .DIN2(n12019), .Q(n12345) );
  nnd2s1 U12484 ( .DIN1(n10957), .DIN2(n10751), .Q(n12019) );
  nnd2s1 U12485 ( .DIN1(n10996), .DIN2(n11379), .Q(n12344) );
  nnd2s1 U12486 ( .DIN1(n10744), .DIN2(n10555), .Q(n12343) );
  nnd2s1 U12487 ( .DIN1(n10546), .DIN2(n11264), .Q(n11249) );
  nnd4s1 U12488 ( .DIN1(n12346), .DIN2(n12347), .DIN3(n12348), .DIN4(n12349), 
        .Q(n12341) );
  nnd2s1 U12489 ( .DIN1(n10758), .DIN2(n12350), .Q(n12349) );
  nnd2s1 U12490 ( .DIN1(n10712), .DIN2(n10754), .Q(n12350) );
  hi1s1 U12491 ( .DIN(n11266), .Q(n10758) );
  nnd2s1 U12492 ( .DIN1(n10714), .DIN2(n12351), .Q(n12348) );
  nnd3s1 U12493 ( .DIN1(n10537), .DIN2(n10548), .DIN3(n10557), .Q(n12351) );
  nnd2s1 U12494 ( .DIN1(n10729), .DIN2(n12352), .Q(n12347) );
  nnd4s1 U12495 ( .DIN1(n10958), .DIN2(n10712), .DIN3(n10558), .DIN4(n10966), 
        .Q(n12352) );
  nnd2s1 U12496 ( .DIN1(n10722), .DIN2(n10542), .Q(n12346) );
  nnd2s1 U12497 ( .DIN1(n10939), .DIN2(n10992), .Q(n10542) );
  nor4s1 U12498 ( .DIN1(n12353), .DIN2(n12354), .DIN3(n12355), .DIN4(n12356), 
        .Q(n12217) );
  nnd4s1 U12499 ( .DIN1(n12357), .DIN2(n12358), .DIN3(n12359), .DIN4(n12360), 
        .Q(n12356) );
  and3s1 U12500 ( .DIN1(n12361), .DIN2(n12362), .DIN3(n12363), .Q(n12360) );
  nnd2s1 U12501 ( .DIN1(n10710), .DIN2(n11787), .Q(n12363) );
  nnd2s1 U12502 ( .DIN1(n10731), .DIN2(n10734), .Q(n11787) );
  nnd2s1 U12503 ( .DIN1(n11329), .DIN2(n12364), .Q(n12362) );
  nnd2s1 U12504 ( .DIN1(n11266), .DIN2(n10964), .Q(n12364) );
  hi1s1 U12505 ( .DIN(n10549), .Q(n11329) );
  nnd2s1 U12506 ( .DIN1(n10532), .DIN2(n12365), .Q(n12361) );
  nnd2s1 U12507 ( .DIN1(n10757), .DIN2(n10725), .Q(n12365) );
  nnd2s1 U12508 ( .DIN1(n10546), .DIN2(n10742), .Q(n12359) );
  nnd2s1 U12509 ( .DIN1(n10752), .DIN2(n12366), .Q(n12358) );
  nnd2s1 U12510 ( .DIN1(n10537), .DIN2(n10539), .Q(n12366) );
  nnd2s1 U12511 ( .DIN1(n11264), .DIN2(n12367), .Q(n12357) );
  nnd2s1 U12512 ( .DIN1(n10756), .DIN2(n10992), .Q(n12367) );
  nnd3s1 U12513 ( .DIN1(n12368), .DIN2(n12369), .DIN3(n12370), .Q(n12355) );
  nnd2s1 U12514 ( .DIN1(n10996), .DIN2(n10952), .Q(n12370) );
  nnd2s1 U12515 ( .DIN1(n10934), .DIN2(n10951), .Q(n12369) );
  nnd2s1 U12516 ( .DIN1(n10990), .DIN2(n10716), .Q(n12368) );
  nor2s1 U12517 ( .DIN1(n10548), .DIN2(n10933), .Q(n12354) );
  nor2s1 U12518 ( .DIN1(n10940), .DIN2(n11271), .Q(n12353) );
  nor4s1 U12519 ( .DIN1(n12371), .DIN2(n12372), .DIN3(n12373), .DIN4(n12374), 
        .Q(n12191) );
  nnd4s1 U12520 ( .DIN1(n12375), .DIN2(n12376), .DIN3(n12377), .DIN4(n12378), 
        .Q(n12374) );
  nnd2s1 U12521 ( .DIN1(n10743), .DIN2(n10951), .Q(n12378) );
  nnd2s1 U12522 ( .DIN1(n10702), .DIN2(n10716), .Q(n12377) );
  nnd2s1 U12523 ( .DIN1(n10533), .DIN2(n10722), .Q(n12376) );
  nnd2s1 U12524 ( .DIN1(n10550), .DIN2(n10541), .Q(n12375) );
  nnd3s1 U12525 ( .DIN1(n12379), .DIN2(n12380), .DIN3(n12381), .Q(n12373) );
  nnd2s1 U12526 ( .DIN1(n10744), .DIN2(n12382), .Q(n12381) );
  nnd2s1 U12527 ( .DIN1(n10757), .DIN2(n11266), .Q(n12382) );
  nnd2s1 U12528 ( .DIN1(n10714), .DIN2(n11359), .Q(n12380) );
  nnd2s1 U12529 ( .DIN1(n10754), .DIN2(n10731), .Q(n11359) );
  nnd2s1 U12530 ( .DIN1(n10742), .DIN2(n12383), .Q(n12379) );
  nnd2s1 U12531 ( .DIN1(n12384), .DIN2(n11266), .Q(n12383) );
  nor2s1 U12532 ( .DIN1(n10549), .DIN2(n10998), .Q(n12372) );
  and2s1 U12533 ( .DIN1(n10555), .DIN2(n12385), .Q(n12371) );
  nnd3s1 U12534 ( .DIN1(n10558), .DIN2(n10754), .DIN3(n10539), .Q(n12385) );
  nnd3s1 U12535 ( .DIN1(n11351), .DIN2(n12386), .DIN3(n12387), .Q(n12334) );
  nnd2s1 U12536 ( .DIN1(n10996), .DIN2(n10702), .Q(n12387) );
  hi1s1 U12537 ( .DIN(n10728), .Q(n10996) );
  nnd2s1 U12538 ( .DIN1(n10743), .DIN2(n10554), .Q(n12386) );
  nnd2s1 U12539 ( .DIN1(n10712), .DIN2(n10549), .Q(n10554) );
  hi1s1 U12540 ( .DIN(n10725), .Q(n10743) );
  nnd2s1 U12541 ( .DIN1(n12388), .DIN2(n12389), .Q(n10725) );
  nnd2s1 U12542 ( .DIN1(n10714), .DIN2(n10951), .Q(n11351) );
  hi1s1 U12543 ( .DIN(n10751), .Q(n10951) );
  hi1s1 U12544 ( .DIN(n10964), .Q(n10714) );
  nnd4s1 U12545 ( .DIN1(n12390), .DIN2(n12391), .DIN3(n12392), .DIN4(n12393), 
        .Q(n12333) );
  nnd2s1 U12546 ( .DIN1(n10550), .DIN2(n12394), .Q(n12393) );
  nnd2s1 U12547 ( .DIN1(n10754), .DIN2(n10549), .Q(n12394) );
  nnd3s1 U12548 ( .DIN1(sa30[7]), .DIN2(n1432), .DIN3(n12395), .Q(n10549) );
  nnd2s1 U12549 ( .DIN1(n10541), .DIN2(n12396), .Q(n12392) );
  nnd2s1 U12550 ( .DIN1(n11368), .DIN2(n11266), .Q(n12396) );
  hi1s1 U12551 ( .DIN(n10741), .Q(n11368) );
  nnd2s1 U12552 ( .DIN1(n10932), .DIN2(n10757), .Q(n10741) );
  nnd2s1 U12553 ( .DIN1(n10732), .DIN2(n12397), .Q(n12391) );
  nnd2s1 U12554 ( .DIN1(n10961), .DIN2(n10731), .Q(n12397) );
  or2s1 U12555 ( .DIN1(n11270), .DIN2(n11362), .Q(n12390) );
  nor2s1 U12556 ( .DIN1(n11264), .DIN2(n10742), .Q(n11362) );
  nor4s1 U12557 ( .DIN1(n12398), .DIN2(n12399), .DIN3(n12400), .DIN4(n12401), 
        .Q(n12192) );
  nnd4s1 U12558 ( .DIN1(n11298), .DIN2(n10526), .DIN3(n12402), .DIN4(n12403), 
        .Q(n12401) );
  nor2s1 U12559 ( .DIN1(n12404), .DIN2(n12405), .Q(n12403) );
  nor2s1 U12560 ( .DIN1(n10739), .DIN2(n11271), .Q(n12405) );
  nor2s1 U12561 ( .DIN1(n12330), .DIN2(n10712), .Q(n12404) );
  nnd2s1 U12562 ( .DIN1(n10729), .DIN2(n10702), .Q(n12402) );
  hi1s1 U12563 ( .DIN(n10932), .Q(n10729) );
  nnd2s1 U12564 ( .DIN1(n12406), .DIN2(n12407), .Q(n10932) );
  nnd2s1 U12565 ( .DIN1(n10722), .DIN2(n10716), .Q(n10526) );
  hi1s1 U12566 ( .DIN(n10958), .Q(n10722) );
  nnd2s1 U12567 ( .DIN1(n10555), .DIN2(n11379), .Q(n11298) );
  nnd3s1 U12568 ( .DIN1(n12408), .DIN2(n12409), .DIN3(n12410), .Q(n12400) );
  nnd2s1 U12569 ( .DIN1(n10701), .DIN2(n10982), .Q(n12410) );
  nnd2s1 U12570 ( .DIN1(n10958), .DIN2(n10734), .Q(n10982) );
  nnd3s1 U12571 ( .DIN1(n12411), .DIN2(n1383), .DIN3(sa30[6]), .Q(n10958) );
  nnd2s1 U12572 ( .DIN1(n10715), .DIN2(n12412), .Q(n12409) );
  nnd3s1 U12573 ( .DIN1(n10739), .DIN2(n11266), .DIN3(n12330), .Q(n12412) );
  hi1s1 U12574 ( .DIN(n10548), .Q(n10715) );
  nnd3s1 U12575 ( .DIN1(sa30[5]), .DIN2(n12411), .DIN3(sa30[6]), .Q(n10548) );
  nnd2s1 U12576 ( .DIN1(n11264), .DIN2(n12413), .Q(n12408) );
  nnd3s1 U12577 ( .DIN1(n10964), .DIN2(n10940), .DIN3(n10998), .Q(n12413) );
  nnd2s1 U12578 ( .DIN1(n12414), .DIN2(n12415), .Q(n10964) );
  hi1s1 U12579 ( .DIN(n10966), .Q(n11264) );
  nor2s1 U12580 ( .DIN1(n10539), .DIN2(n11266), .Q(n12399) );
  nnd2s1 U12581 ( .DIN1(n12407), .DIN2(n12389), .Q(n11266) );
  nor2s1 U12582 ( .DIN1(n11369), .DIN2(n10751), .Q(n12398) );
  nnd3s1 U12583 ( .DIN1(sa30[4]), .DIN2(n1383), .DIN3(n12416), .Q(n10751) );
  nor2s1 U12584 ( .DIN1(n10546), .DIN2(n10752), .Q(n11369) );
  nor2s1 U12585 ( .DIN1(n12417), .DIN2(n12418), .Q(n12020) );
  nnd4s1 U12586 ( .DIN1(n12419), .DIN2(n12420), .DIN3(n12421), .DIN4(n12422), 
        .Q(n12418) );
  nnd2s1 U12587 ( .DIN1(n10749), .DIN2(n10990), .Q(n12422) );
  hi1s1 U12588 ( .DIN(n10558), .Q(n10990) );
  nnd2s1 U12589 ( .DIN1(n12395), .DIN2(n12423), .Q(n10558) );
  hi1s1 U12590 ( .DIN(n10933), .Q(n10749) );
  nnd2s1 U12591 ( .DIN1(n11379), .DIN2(n10701), .Q(n12421) );
  hi1s1 U12592 ( .DIN(n10731), .Q(n11379) );
  nnd2s1 U12593 ( .DIN1(n10550), .DIN2(n10702), .Q(n12420) );
  hi1s1 U12594 ( .DIN(n10961), .Q(n10702) );
  nnd2s1 U12595 ( .DIN1(n10533), .DIN2(n10952), .Q(n12419) );
  hi1s1 U12596 ( .DIN(n10539), .Q(n10952) );
  hi1s1 U12597 ( .DIN(n10739), .Q(n10533) );
  nnd2s1 U12598 ( .DIN1(n12424), .DIN2(n12388), .Q(n10739) );
  nnd4s1 U12599 ( .DIN1(n12425), .DIN2(n12426), .DIN3(n12427), .DIN4(n12428), 
        .Q(n12417) );
  nnd2s1 U12600 ( .DIN1(n10744), .DIN2(n12429), .Q(n12428) );
  nnd2s1 U12601 ( .DIN1(n10998), .DIN2(n10992), .Q(n12429) );
  nnd2s1 U12602 ( .DIN1(n10532), .DIN2(n12430), .Q(n12427) );
  or2s1 U12603 ( .DIN1(n11380), .DIN2(n10732), .Q(n12430) );
  nnd2s1 U12604 ( .DIN1(n10992), .DIN2(n10933), .Q(n11380) );
  hi1s1 U12605 ( .DIN(n10754), .Q(n10532) );
  nnd3s1 U12606 ( .DIN1(sa30[5]), .DIN2(sa30[4]), .DIN3(n12416), .Q(n10754) );
  nnd2s1 U12607 ( .DIN1(n10717), .DIN2(n12431), .Q(n12426) );
  or2s1 U12608 ( .DIN1(n10983), .DIN2(n10701), .Q(n12431) );
  hi1s1 U12609 ( .DIN(n10940), .Q(n10701) );
  nnd2s1 U12610 ( .DIN1(n12432), .DIN2(n12389), .Q(n10940) );
  nnd2s1 U12611 ( .DIN1(n11270), .DIN2(n10728), .Q(n10983) );
  nnd2s1 U12612 ( .DIN1(n12406), .DIN2(n12432), .Q(n10728) );
  hi1s1 U12613 ( .DIN(n10537), .Q(n10717) );
  nnd3s1 U12614 ( .DIN1(sa30[5]), .DIN2(sa30[4]), .DIN3(n12423), .Q(n10537) );
  nnd2s1 U12615 ( .DIN1(n10541), .DIN2(n12433), .Q(n12425) );
  nnd3s1 U12616 ( .DIN1(n10998), .DIN2(n10933), .DIN3(n12384), .Q(n12433) );
  nor2s1 U12617 ( .DIN1(n10732), .DIN2(n10752), .Q(n12384) );
  hi1s1 U12618 ( .DIN(n10756), .Q(n10732) );
  nnd2s1 U12619 ( .DIN1(n12406), .DIN2(n12415), .Q(n10933) );
  hi1s1 U12620 ( .DIN(n11271), .Q(n10541) );
  nnd3s1 U12621 ( .DIN1(n12434), .DIN2(n12435), .DIN3(n12436), .Q(n12313) );
  nnd2s1 U12622 ( .DIN1(n10550), .DIN2(n10744), .Q(n12436) );
  hi1s1 U12623 ( .DIN(n10557), .Q(n10744) );
  nnd3s1 U12624 ( .DIN1(sa30[6]), .DIN2(sa30[7]), .DIN3(n12395), .Q(n10557) );
  hi1s1 U12625 ( .DIN(n10724), .Q(n10550) );
  nnd2s1 U12626 ( .DIN1(n12424), .DIN2(n12407), .Q(n10724) );
  nnd2s1 U12627 ( .DIN1(n10752), .DIN2(n11347), .Q(n12435) );
  nnd2s1 U12628 ( .DIN1(n10966), .DIN2(n10731), .Q(n11347) );
  nnd3s1 U12629 ( .DIN1(n12411), .DIN2(n1432), .DIN3(sa30[5]), .Q(n10731) );
  nnd3s1 U12630 ( .DIN1(sa30[6]), .DIN2(sa30[7]), .DIN3(n12437), .Q(n10966) );
  hi1s1 U12631 ( .DIN(n12330), .Q(n10752) );
  nnd2s1 U12632 ( .DIN1(n12415), .DIN2(n12389), .Q(n12330) );
  and2s1 U12633 ( .DIN1(sa30[0]), .DIN2(n1538), .Q(n12389) );
  nnd2s1 U12634 ( .DIN1(n10742), .DIN2(n10716), .Q(n12434) );
  hi1s1 U12635 ( .DIN(n10757), .Q(n10716) );
  nnd2s1 U12636 ( .DIN1(n12414), .DIN2(n12407), .Q(n10757) );
  and2s1 U12637 ( .DIN1(sa30[3]), .DIN2(n1533), .Q(n12407) );
  hi1s1 U12638 ( .DIN(n10734), .Q(n10742) );
  nnd2s1 U12639 ( .DIN1(n12423), .DIN2(n12437), .Q(n10734) );
  nnd4s1 U12640 ( .DIN1(n12438), .DIN2(n12439), .DIN3(n12440), .DIN4(n12441), 
        .Q(n12312) );
  nnd2s1 U12641 ( .DIN1(n10934), .DIN2(n12442), .Q(n12441) );
  nnd2s1 U12642 ( .DIN1(n11271), .DIN2(n10539), .Q(n12442) );
  hi1s1 U12643 ( .DIN(n10992), .Q(n10934) );
  nnd2s1 U12644 ( .DIN1(n12414), .DIN2(n12432), .Q(n10992) );
  nnd2s1 U12645 ( .DIN1(n10710), .DIN2(n12443), .Q(n12440) );
  nnd2s1 U12646 ( .DIN1(n10539), .DIN2(n10961), .Q(n12443) );
  nnd3s1 U12647 ( .DIN1(sa30[7]), .DIN2(n1432), .DIN3(n12437), .Q(n10961) );
  nnd2s1 U12648 ( .DIN1(n12416), .DIN2(n12437), .Q(n10539) );
  nor2s1 U12649 ( .DIN1(n1383), .DIN2(sa30[4]), .Q(n12437) );
  hi1s1 U12650 ( .DIN(n10998), .Q(n10710) );
  nnd2s1 U12651 ( .DIN1(n12415), .DIN2(n12424), .Q(n10998) );
  nor2s1 U12652 ( .DIN1(sa30[3]), .DIN2(sa30[1]), .Q(n12415) );
  nnd2s1 U12653 ( .DIN1(n10555), .DIN2(n12444), .Q(n12439) );
  nnd2s1 U12654 ( .DIN1(n11271), .DIN2(n10957), .Q(n12444) );
  nnd2s1 U12655 ( .DIN1(n12395), .DIN2(n12416), .Q(n10957) );
  nor2s1 U12656 ( .DIN1(n1432), .DIN2(sa30[7]), .Q(n12416) );
  nor2s1 U12657 ( .DIN1(sa30[5]), .DIN2(sa30[4]), .Q(n12395) );
  nnd3s1 U12658 ( .DIN1(sa30[4]), .DIN2(n1383), .DIN3(n12423), .Q(n11271) );
  nor2s1 U12659 ( .DIN1(sa30[7]), .DIN2(sa30[6]), .Q(n12423) );
  nnd2s1 U12660 ( .DIN1(n10937), .DIN2(n12445), .Q(n12438) );
  nnd2s1 U12661 ( .DIN1(n11779), .DIN2(n10756), .Q(n12445) );
  nnd2s1 U12662 ( .DIN1(n12432), .DIN2(n12424), .Q(n10756) );
  nor2s1 U12663 ( .DIN1(sa30[2]), .DIN2(sa30[0]), .Q(n12424) );
  and2s1 U12664 ( .DIN1(sa30[1]), .DIN2(sa30[3]), .Q(n12432) );
  nor2s1 U12665 ( .DIN1(n10546), .DIN2(n10555), .Q(n11779) );
  hi1s1 U12666 ( .DIN(n11270), .Q(n10555) );
  nnd2s1 U12667 ( .DIN1(n12414), .DIN2(n12388), .Q(n11270) );
  and2s1 U12668 ( .DIN1(sa30[2]), .DIN2(sa30[0]), .Q(n12414) );
  hi1s1 U12669 ( .DIN(n10939), .Q(n10546) );
  nnd2s1 U12670 ( .DIN1(n12406), .DIN2(n12388), .Q(n10939) );
  nor2s1 U12671 ( .DIN1(n1533), .DIN2(sa30[3]), .Q(n12388) );
  nor2s1 U12672 ( .DIN1(n1538), .DIN2(sa30[0]), .Q(n12406) );
  hi1s1 U12673 ( .DIN(n10712), .Q(n10937) );
  nnd3s1 U12674 ( .DIN1(n1383), .DIN2(n1432), .DIN3(n12411), .Q(n10712) );
  and2s1 U12675 ( .DIN1(sa30[7]), .DIN2(sa30[4]), .Q(n12411) );
  or3s1 U12676 ( .DIN1(n12446), .DIN2(n12447), .DIN3(n12448), .Q(n5701) );
  nnd4s1 U12677 ( .DIN1(n12151), .DIN2(n12449), .DIN3(n11988), .DIN4(n12450), 
        .Q(n12448) );
  and4s1 U12678 ( .DIN1(n12451), .DIN2(n12452), .DIN3(n12453), .DIN4(n10864), 
        .Q(n12450) );
  nnd2s1 U12679 ( .DIN1(n10877), .DIN2(n10681), .Q(n10864) );
  nnd2s1 U12680 ( .DIN1(n10904), .DIN2(n10663), .Q(n12453) );
  nnd2s1 U12681 ( .DIN1(n10685), .DIN2(n10867), .Q(n12452) );
  nor3s1 U12682 ( .DIN1(n12454), .DIN2(n12455), .DIN3(n12456), .Q(n11988) );
  nnd4s1 U12683 ( .DIN1(n12457), .DIN2(n12458), .DIN3(n12152), .DIN4(n12459), 
        .Q(n12456) );
  and3s1 U12684 ( .DIN1(n12460), .DIN2(n12461), .DIN3(n12462), .Q(n12459) );
  nnd2s1 U12685 ( .DIN1(n10677), .DIN2(n10867), .Q(n12462) );
  nnd2s1 U12686 ( .DIN1(n10877), .DIN2(n11172), .Q(n12461) );
  nnd2s1 U12687 ( .DIN1(n10893), .DIN2(n10876), .Q(n12460) );
  nor2s1 U12688 ( .DIN1(n12463), .DIN2(n12464), .Q(n12152) );
  nnd4s1 U12689 ( .DIN1(n12465), .DIN2(n12466), .DIN3(n11754), .DIN4(n12467), 
        .Q(n12464) );
  nnd2s1 U12690 ( .DIN1(n10664), .DIN2(n10673), .Q(n12467) );
  nnd2s1 U12691 ( .DIN1(n11244), .DIN2(n11220), .Q(n10673) );
  nnd2s1 U12692 ( .DIN1(n10677), .DIN2(n11642), .Q(n11754) );
  nnd2s1 U12693 ( .DIN1(n11199), .DIN2(n11173), .Q(n12466) );
  nnd2s1 U12694 ( .DIN1(n10867), .DIN2(n10681), .Q(n12465) );
  nnd4s1 U12695 ( .DIN1(n12468), .DIN2(n12469), .DIN3(n12470), .DIN4(n12471), 
        .Q(n12463) );
  nnd2s1 U12696 ( .DIN1(n10884), .DIN2(n12472), .Q(n12471) );
  nnd2s1 U12697 ( .DIN1(n11646), .DIN2(n11185), .Q(n12472) );
  nnd2s1 U12698 ( .DIN1(n10901), .DIN2(n12473), .Q(n12470) );
  nnd2s1 U12699 ( .DIN1(n10895), .DIN2(n10912), .Q(n12473) );
  nnd2s1 U12700 ( .DIN1(n10866), .DIN2(n12474), .Q(n12469) );
  nnd3s1 U12701 ( .DIN1(n10684), .DIN2(n10680), .DIN3(n10668), .Q(n12474) );
  nnd2s1 U12702 ( .DIN1(n10887), .DIN2(n12475), .Q(n12468) );
  nnd4s1 U12703 ( .DIN1(n10874), .DIN2(n10895), .DIN3(n11188), .DIN4(n10683), 
        .Q(n12475) );
  nnd3s1 U12704 ( .DIN1(n12476), .DIN2(n12477), .DIN3(n11730), .Q(n12455) );
  nnd2s1 U12705 ( .DIN1(n10866), .DIN2(n11705), .Q(n11730) );
  or2s1 U12706 ( .DIN1(n11704), .DIN2(n11738), .Q(n12477) );
  nor2s1 U12707 ( .DIN1(n10904), .DIN2(n11642), .Q(n11738) );
  nnd2s1 U12708 ( .DIN1(n10905), .DIN2(n10689), .Q(n12476) );
  nnd2s1 U12709 ( .DIN1(n10895), .DIN2(n10679), .Q(n10689) );
  nnd4s1 U12710 ( .DIN1(n12478), .DIN2(n12479), .DIN3(n12480), .DIN4(n12481), 
        .Q(n12454) );
  nnd2s1 U12711 ( .DIN1(n11173), .DIN2(n12004), .Q(n12481) );
  nnd2s1 U12712 ( .DIN1(n11219), .DIN2(n10917), .Q(n12004) );
  nnd2s1 U12713 ( .DIN1(n10685), .DIN2(n12482), .Q(n12480) );
  nnd2s1 U12714 ( .DIN1(n10679), .DIN2(n10912), .Q(n12482) );
  nnd2s1 U12715 ( .DIN1(n10865), .DIN2(n12483), .Q(n12479) );
  nnd2s1 U12716 ( .DIN1(n10892), .DIN2(n10917), .Q(n12483) );
  nnd2s1 U12717 ( .DIN1(n10672), .DIN2(n12484), .Q(n12478) );
  nnd2s1 U12718 ( .DIN1(n11746), .DIN2(n11637), .Q(n12484) );
  hi1s1 U12719 ( .DIN(n10903), .Q(n11746) );
  nnd2s1 U12720 ( .DIN1(n11215), .DIN2(n10916), .Q(n10903) );
  nor2s1 U12721 ( .DIN1(n12485), .DIN2(n12486), .Q(n12151) );
  nnd4s1 U12722 ( .DIN1(n12487), .DIN2(n12488), .DIN3(n12489), .DIN4(n12490), 
        .Q(n12486) );
  nnd2s1 U12723 ( .DIN1(n10878), .DIN2(n11207), .Q(n12490) );
  nnd2s1 U12724 ( .DIN1(n10892), .DIN2(n11704), .Q(n11207) );
  nnd2s1 U12725 ( .DIN1(n11174), .DIN2(n10662), .Q(n12489) );
  nnd2s1 U12726 ( .DIN1(n10685), .DIN2(n10865), .Q(n12488) );
  nnd2s1 U12727 ( .DIN1(n10913), .DIN2(n11198), .Q(n12487) );
  nnd4s1 U12728 ( .DIN1(n12491), .DIN2(n12492), .DIN3(n12493), .DIN4(n12494), 
        .Q(n12485) );
  nnd2s1 U12729 ( .DIN1(n10661), .DIN2(n12495), .Q(n12494) );
  or2s1 U12730 ( .DIN1(n11757), .DIN2(n10884), .Q(n12495) );
  nnd2s1 U12731 ( .DIN1(n10879), .DIN2(n12496), .Q(n12493) );
  nnd2s1 U12732 ( .DIN1(n10668), .DIN2(n10889), .Q(n12496) );
  nnd2s1 U12733 ( .DIN1(n10867), .DIN2(n12497), .Q(n12492) );
  nnd2s1 U12734 ( .DIN1(n11225), .DIN2(n11220), .Q(n12497) );
  nnd2s1 U12735 ( .DIN1(n10672), .DIN2(n12498), .Q(n12491) );
  nnd3s1 U12736 ( .DIN1(n11225), .DIN2(n11219), .DIN3(n12499), .Q(n12498) );
  nnd4s1 U12737 ( .DIN1(n11223), .DIN2(n12500), .DIN3(n12501), .DIN4(n12502), 
        .Q(n12447) );
  nnd2s1 U12738 ( .DIN1(n11172), .DIN2(n11174), .Q(n12502) );
  nnd2s1 U12739 ( .DIN1(n10662), .DIN2(n11642), .Q(n12501) );
  nnd2s1 U12740 ( .DIN1(n10884), .DIN2(n10878), .Q(n12500) );
  nnd2s1 U12741 ( .DIN1(n10887), .DIN2(n10876), .Q(n11223) );
  nnd4s1 U12742 ( .DIN1(n12503), .DIN2(n12504), .DIN3(n12505), .DIN4(n12506), 
        .Q(n12446) );
  nnd2s1 U12743 ( .DIN1(n11242), .DIN2(n12507), .Q(n12506) );
  nnd2s1 U12744 ( .DIN1(n11996), .DIN2(n10917), .Q(n12507) );
  nor2s1 U12745 ( .DIN1(n10677), .DIN2(n10681), .Q(n11996) );
  nnd2s1 U12746 ( .DIN1(n10893), .DIN2(n12508), .Q(n12505) );
  nnd2s1 U12747 ( .DIN1(n11180), .DIN2(n10670), .Q(n12508) );
  nnd2s1 U12748 ( .DIN1(n10672), .DIN2(n12509), .Q(n12504) );
  nnd2s1 U12749 ( .DIN1(n11704), .DIN2(n11220), .Q(n12509) );
  nnd2s1 U12750 ( .DIN1(n10910), .DIN2(n11725), .Q(n12503) );
  xor2s1 U12751 ( .DIN1(n5422), .DIN2(n5069), .Q(n10308) );
  nor4s1 U12752 ( .DIN1(n12510), .DIN2(n12511), .DIN3(n12512), .DIN4(n12513), 
        .Q(n5069) );
  nnd4s1 U12753 ( .DIN1(n11079), .DIN2(n12514), .DIN3(n12515), .DIN4(n12516), 
        .Q(n12513) );
  nnd2s1 U12754 ( .DIN1(n10809), .DIN2(n11613), .Q(n12516) );
  nnd2s1 U12755 ( .DIN1(n11133), .DIN2(n10518), .Q(n11613) );
  nnd2s1 U12756 ( .DIN1(n10850), .DIN2(n10520), .Q(n12515) );
  nnd2s1 U12757 ( .DIN1(n10829), .DIN2(n11102), .Q(n10520) );
  nnd2s1 U12758 ( .DIN1(n11562), .DIN2(n10820), .Q(n12514) );
  nnd2s1 U12759 ( .DIN1(n10843), .DIN2(n10500), .Q(n11079) );
  nnd4s1 U12760 ( .DIN1(n12517), .DIN2(n12518), .DIN3(n12519), .DIN4(n12520), 
        .Q(n12512) );
  nnd2s1 U12761 ( .DIN1(n10491), .DIN2(n12521), .Q(n12520) );
  nnd2s1 U12762 ( .DIN1(n10642), .DIN2(n10817), .Q(n12521) );
  nnd2s1 U12763 ( .DIN1(n10808), .DIN2(n12522), .Q(n12519) );
  nnd2s1 U12764 ( .DIN1(n11137), .DIN2(n11129), .Q(n12522) );
  or2s1 U12765 ( .DIN1(n10849), .DIN2(n10831), .Q(n12518) );
  nor2s1 U12766 ( .DIN1(n10511), .DIN2(n10820), .Q(n10831) );
  nnd2s1 U12767 ( .DIN1(n11113), .DIN2(n10841), .Q(n12517) );
  nnd2s1 U12768 ( .DIN1(n10826), .DIN2(n10641), .Q(n10841) );
  nnd3s1 U12769 ( .DIN1(n11948), .DIN2(n11956), .DIN3(n10482), .Q(n12511) );
  nor4s1 U12770 ( .DIN1(n12523), .DIN2(n12524), .DIN3(n12525), .DIN4(n12526), 
        .Q(n10482) );
  nnd4s1 U12771 ( .DIN1(n12527), .DIN2(n12528), .DIN3(n12529), .DIN4(n12530), 
        .Q(n12526) );
  nnd2s1 U12772 ( .DIN1(n10515), .DIN2(n10499), .Q(n12530) );
  nor2s1 U12773 ( .DIN1(n12531), .DIN2(n11532), .Q(n12529) );
  nor2s1 U12774 ( .DIN1(n10829), .DIN2(n10517), .Q(n11532) );
  nor2s1 U12775 ( .DIN1(n10817), .DIN2(n10853), .Q(n12531) );
  nnd2s1 U12776 ( .DIN1(n10840), .DIN2(n10498), .Q(n12528) );
  nnd2s1 U12777 ( .DIN1(n10809), .DIN2(n10827), .Q(n12527) );
  hi1s1 U12778 ( .DIN(n10513), .Q(n10809) );
  nnd3s1 U12779 ( .DIN1(n12532), .DIN2(n12533), .DIN3(n12534), .Q(n12525) );
  nnd2s1 U12780 ( .DIN1(n10820), .DIN2(n11120), .Q(n12534) );
  nnd2s1 U12781 ( .DIN1(n10826), .DIN2(n10817), .Q(n11120) );
  nnd2s1 U12782 ( .DIN1(n10500), .DIN2(n12535), .Q(n12533) );
  nnd3s1 U12783 ( .DIN1(n11130), .DIN2(n11497), .DIN3(n11137), .Q(n12535) );
  nnd2s1 U12784 ( .DIN1(n10819), .DIN2(n12536), .Q(n12532) );
  nnd3s1 U12785 ( .DIN1(n11132), .DIN2(n11496), .DIN3(n11100), .Q(n12536) );
  nor2s1 U12786 ( .DIN1(n11100), .DIN2(n10834), .Q(n12524) );
  nor2s1 U12787 ( .DIN1(n11603), .DIN2(n11099), .Q(n12523) );
  nor2s1 U12788 ( .DIN1(n10639), .DIN2(n10519), .Q(n11603) );
  and4s1 U12789 ( .DIN1(n12537), .DIN2(n12538), .DIN3(n12539), .DIN4(n12540), 
        .Q(n11956) );
  and4s1 U12790 ( .DIN1(n12541), .DIN2(n11546), .DIN3(n12542), .DIN4(n12543), 
        .Q(n12540) );
  nnd2s1 U12791 ( .DIN1(n10843), .DIN2(n11562), .Q(n12543) );
  nnd2s1 U12792 ( .DIN1(n10499), .DIN2(n10628), .Q(n12542) );
  nnd2s1 U12793 ( .DIN1(n10511), .DIN2(n11567), .Q(n11546) );
  nnd2s1 U12794 ( .DIN1(n10491), .DIN2(n10515), .Q(n12541) );
  and3s1 U12795 ( .DIN1(n12544), .DIN2(n12545), .DIN3(n12546), .Q(n12539) );
  nnd2s1 U12796 ( .DIN1(n10840), .DIN2(n12547), .Q(n12546) );
  nnd2s1 U12797 ( .DIN1(n10646), .DIN2(n10826), .Q(n12547) );
  nnd2s1 U12798 ( .DIN1(n10490), .DIN2(n12548), .Q(n12545) );
  nnd2s1 U12799 ( .DIN1(n10513), .DIN2(n10646), .Q(n12548) );
  nnd2s1 U12800 ( .DIN1(n10810), .DIN2(n11595), .Q(n12544) );
  nnd2s1 U12801 ( .DIN1(n10829), .DIN2(n10849), .Q(n11595) );
  nnd2s1 U12802 ( .DIN1(n10643), .DIN2(n12549), .Q(n12538) );
  nnd3s1 U12803 ( .DIN1(n10849), .DIN2(n10645), .DIN3(n10514), .Q(n12549) );
  hi1s1 U12804 ( .DIN(n10517), .Q(n10643) );
  or2s1 U12805 ( .DIN1(n10826), .DIN2(n12133), .Q(n12537) );
  nor2s1 U12806 ( .DIN1(n10501), .DIN2(n10519), .Q(n12133) );
  nor4s1 U12807 ( .DIN1(n12550), .DIN2(n12551), .DIN3(n12552), .DIN4(n12553), 
        .Q(n11948) );
  nnd4s1 U12808 ( .DIN1(n12554), .DIN2(n12555), .DIN3(n12556), .DIN4(n12557), 
        .Q(n12553) );
  nor2s1 U12809 ( .DIN1(n12558), .DIN2(n12559), .Q(n12557) );
  nor2s1 U12810 ( .DIN1(n11130), .DIN2(n10641), .Q(n12559) );
  nor2s1 U12811 ( .DIN1(n11132), .DIN2(n10646), .Q(n12558) );
  nnd2s1 U12812 ( .DIN1(n10827), .DIN2(n11089), .Q(n12556) );
  or2s1 U12813 ( .DIN1(n11533), .DIN2(n11094), .Q(n12555) );
  nor2s1 U12814 ( .DIN1(n10515), .DIN2(n11089), .Q(n11094) );
  nnd2s1 U12815 ( .DIN1(n10489), .DIN2(n10497), .Q(n12554) );
  nnd3s1 U12816 ( .DIN1(n12560), .DIN2(n12561), .DIN3(n12562), .Q(n12552) );
  nnd2s1 U12817 ( .DIN1(n10490), .DIN2(n11153), .Q(n12562) );
  nnd2s1 U12818 ( .DIN1(n10641), .DIN2(n11102), .Q(n11153) );
  hi1s1 U12819 ( .DIN(n10853), .Q(n10490) );
  nnd2s1 U12820 ( .DIN1(n10628), .DIN2(n12563), .Q(n12561) );
  nnd2s1 U12821 ( .DIN1(n11496), .DIN2(n10832), .Q(n12563) );
  nnd2s1 U12822 ( .DIN1(n10819), .DIN2(n12564), .Q(n12560) );
  nnd2s1 U12823 ( .DIN1(n10510), .DIN2(n11533), .Q(n12564) );
  nor2s1 U12824 ( .DIN1(n12565), .DIN2(n10514), .Q(n12551) );
  nor2s1 U12825 ( .DIN1(n10491), .DIN2(n10810), .Q(n12565) );
  nor2s1 U12826 ( .DIN1(n12566), .DIN2(n10632), .Q(n12550) );
  nor2s1 U12827 ( .DIN1(n10497), .DIN2(n10639), .Q(n12566) );
  nnd4s1 U12828 ( .DIN1(n12090), .DIN2(n12567), .DIN3(n12568), .DIN4(n12569), 
        .Q(n12510) );
  nnd2s1 U12829 ( .DIN1(n10489), .DIN2(n10827), .Q(n12569) );
  nnd2s1 U12830 ( .DIN1(n10810), .DIN2(n10515), .Q(n12568) );
  nnd2s1 U12831 ( .DIN1(n11112), .DIN2(n10840), .Q(n12567) );
  nor3s1 U12832 ( .DIN1(n12570), .DIN2(n12571), .DIN3(n12572), .Q(n12090) );
  nnd4s1 U12833 ( .DIN1(n10485), .DIN2(n11957), .DIN3(n11952), .DIN4(n12573), 
        .Q(n12572) );
  and3s1 U12834 ( .DIN1(n12574), .DIN2(n12575), .DIN3(n12576), .Q(n12573) );
  nnd2s1 U12835 ( .DIN1(n10808), .DIN2(n10840), .Q(n12576) );
  nnd2s1 U12836 ( .DIN1(n10492), .DIN2(n10827), .Q(n12575) );
  hi1s1 U12837 ( .DIN(n11129), .Q(n10827) );
  hi1s1 U12838 ( .DIN(n10646), .Q(n10492) );
  nnd2s1 U12839 ( .DIN1(n11113), .DIN2(n10507), .Q(n12574) );
  hi1s1 U12840 ( .DIN(n10834), .Q(n10507) );
  and4s1 U12841 ( .DIN1(n12577), .DIN2(n12578), .DIN3(n12579), .DIN4(n12580), 
        .Q(n11952) );
  and4s1 U12842 ( .DIN1(n12581), .DIN2(n12582), .DIN3(n11511), .DIN4(n11087), 
        .Q(n12580) );
  nnd2s1 U12843 ( .DIN1(n10501), .DIN2(n10628), .Q(n11087) );
  nnd2s1 U12844 ( .DIN1(n10810), .DIN2(n10489), .Q(n11511) );
  nnd2s1 U12845 ( .DIN1(n10639), .DIN2(n10515), .Q(n12582) );
  nnd2s1 U12846 ( .DIN1(n10808), .DIN2(n11113), .Q(n12581) );
  and3s1 U12847 ( .DIN1(n12583), .DIN2(n12584), .DIN3(n12585), .Q(n12579) );
  nnd2s1 U12848 ( .DIN1(n10502), .DIN2(n12102), .Q(n12585) );
  nnd2s1 U12849 ( .DIN1(n11098), .DIN2(n10853), .Q(n12102) );
  nnd2s1 U12850 ( .DIN1(n10499), .DIN2(n12586), .Q(n12584) );
  nnd2s1 U12851 ( .DIN1(n11540), .DIN2(n10834), .Q(n12586) );
  nor2s1 U12852 ( .DIN1(n11112), .DIN2(n11089), .Q(n11540) );
  hi1s1 U12853 ( .DIN(n10829), .Q(n11089) );
  nnd2s1 U12854 ( .DIN1(n11567), .DIN2(n12587), .Q(n12583) );
  nnd2s1 U12855 ( .DIN1(n11133), .DIN2(n10517), .Q(n12587) );
  nnd2s1 U12856 ( .DIN1(n11112), .DIN2(n12588), .Q(n12578) );
  nnd2s1 U12857 ( .DIN1(n11155), .DIN2(n10510), .Q(n12588) );
  nnd2s1 U12858 ( .DIN1(n10820), .DIN2(n12589), .Q(n12577) );
  nnd3s1 U12859 ( .DIN1(n10642), .DIN2(n10514), .DIN3(n10646), .Q(n12589) );
  and4s1 U12860 ( .DIN1(n12590), .DIN2(n12591), .DIN3(n12592), .DIN4(n12593), 
        .Q(n11957) );
  nor4s1 U12861 ( .DIN1(n12594), .DIN2(n12595), .DIN3(n12596), .DIN4(n12597), 
        .Q(n12593) );
  nor2s1 U12862 ( .DIN1(n12598), .DIN2(n10641), .Q(n12597) );
  nor2s1 U12863 ( .DIN1(n10810), .DIN2(n10840), .Q(n12598) );
  nor2s1 U12864 ( .DIN1(n12599), .DIN2(n11102), .Q(n12596) );
  nor2s1 U12865 ( .DIN1(n10497), .DIN2(n10501), .Q(n12599) );
  hi1s1 U12866 ( .DIN(n10510), .Q(n10501) );
  nnd3s1 U12867 ( .DIN1(n12600), .DIN2(n1365), .DIN3(sa12[1]), .Q(n10510) );
  nor2s1 U12868 ( .DIN1(n12601), .DIN2(n10853), .Q(n12595) );
  nor2s1 U12869 ( .DIN1(n10627), .DIN2(n11112), .Q(n12601) );
  nnd3s1 U12870 ( .DIN1(n12602), .DIN2(n12603), .DIN3(n12604), .Q(n12594) );
  nnd2s1 U12871 ( .DIN1(n10497), .DIN2(n11562), .Q(n12604) );
  nnd2s1 U12872 ( .DIN1(n10498), .DIN2(n12605), .Q(n12603) );
  nnd2s1 U12873 ( .DIN1(n10832), .DIN2(n11100), .Q(n12605) );
  nnd2s1 U12874 ( .DIN1(n10511), .DIN2(n11982), .Q(n12602) );
  nnd2s1 U12875 ( .DIN1(n10826), .DIN2(n10829), .Q(n11982) );
  nnd2s1 U12876 ( .DIN1(n12606), .DIN2(n12607), .Q(n10829) );
  hi1s1 U12877 ( .DIN(n11137), .Q(n10511) );
  and3s1 U12878 ( .DIN1(n12608), .DIN2(n12609), .DIN3(n12610), .Q(n12592) );
  nnd2s1 U12879 ( .DIN1(n10850), .DIN2(n10819), .Q(n12610) );
  hi1s1 U12880 ( .DIN(n10642), .Q(n10819) );
  nnd2s1 U12881 ( .DIN1(n10627), .DIN2(n10843), .Q(n12609) );
  nnd2s1 U12882 ( .DIN1(n10502), .DIN2(n10519), .Q(n12608) );
  nnd2s1 U12883 ( .DIN1(n10639), .DIN2(n10489), .Q(n12591) );
  nnd2s1 U12884 ( .DIN1(n10515), .DIN2(n10820), .Q(n12590) );
  hi1s1 U12885 ( .DIN(n11130), .Q(n10820) );
  hi1s1 U12886 ( .DIN(n11557), .Q(n10515) );
  nnd2s1 U12887 ( .DIN1(n12606), .DIN2(n12611), .Q(n11557) );
  nor4s1 U12888 ( .DIN1(n12612), .DIN2(n12613), .DIN3(n12614), .DIN4(n12615), 
        .Q(n10485) );
  nnd4s1 U12889 ( .DIN1(n12616), .DIN2(n12617), .DIN3(n12618), .DIN4(n12619), 
        .Q(n12615) );
  nnd2s1 U12890 ( .DIN1(n10843), .DIN2(n10498), .Q(n12619) );
  hi1s1 U12891 ( .DIN(n11533), .Q(n10843) );
  nnd2s1 U12892 ( .DIN1(n10491), .DIN2(n10500), .Q(n12618) );
  hi1s1 U12893 ( .DIN(n11102), .Q(n10500) );
  nnd2s1 U12894 ( .DIN1(n12620), .DIN2(n12607), .Q(n11102) );
  hi1s1 U12895 ( .DIN(n11098), .Q(n10491) );
  nnd3s1 U12896 ( .DIN1(n1365), .DIN2(n1433), .DIN3(n12600), .Q(n11098) );
  nnd2s1 U12897 ( .DIN1(n10627), .DIN2(n10519), .Q(n12617) );
  hi1s1 U12898 ( .DIN(n11100), .Q(n10519) );
  hi1s1 U12899 ( .DIN(n10849), .Q(n10627) );
  nnd2s1 U12900 ( .DIN1(n10489), .DIN2(n10499), .Q(n12616) );
  hi1s1 U12901 ( .DIN(n10826), .Q(n10489) );
  nnd2s1 U12902 ( .DIN1(n12621), .DIN2(n12622), .Q(n10826) );
  nnd3s1 U12903 ( .DIN1(n12623), .DIN2(n12624), .DIN3(n12625), .Q(n12614) );
  nnd2s1 U12904 ( .DIN1(n10808), .DIN2(n12626), .Q(n12625) );
  nnd3s1 U12905 ( .DIN1(n10853), .DIN2(n11130), .DIN3(n11100), .Q(n12626) );
  nnd3s1 U12906 ( .DIN1(n12627), .DIN2(n1446), .DIN3(sa12[0]), .Q(n11100) );
  nnd3s1 U12907 ( .DIN1(sa12[0]), .DIN2(n1433), .DIN3(n12628), .Q(n10853) );
  hi1s1 U12908 ( .DIN(n11504), .Q(n10808) );
  nnd2s1 U12909 ( .DIN1(n10502), .DIN2(n12629), .Q(n12624) );
  nnd2s1 U12910 ( .DIN1(n11129), .DIN2(n11533), .Q(n12629) );
  nnd3s1 U12911 ( .DIN1(n1365), .DIN2(n1433), .DIN3(n12628), .Q(n11129) );
  hi1s1 U12912 ( .DIN(n10632), .Q(n10502) );
  nnd2s1 U12913 ( .DIN1(n10840), .DIN2(n12630), .Q(n12623) );
  nnd2s1 U12914 ( .DIN1(n10513), .DIN2(n11099), .Q(n12630) );
  nnd2s1 U12915 ( .DIN1(n12621), .DIN2(n12607), .Q(n10513) );
  hi1s1 U12916 ( .DIN(n11496), .Q(n10840) );
  nnd3s1 U12917 ( .DIN1(sa12[0]), .DIN2(n1433), .DIN3(n12600), .Q(n11496) );
  nor2s1 U12918 ( .DIN1(n10834), .DIN2(n10518), .Q(n12613) );
  nnd2s1 U12919 ( .DIN1(n12606), .DIN2(n12631), .Q(n10834) );
  and2s1 U12920 ( .DIN1(n11113), .DIN2(n12632), .Q(n12612) );
  nnd4s1 U12921 ( .DIN1(n10646), .DIN2(n10642), .DIN3(n10849), .DIN4(n10645), 
        .Q(n12632) );
  nnd2s1 U12922 ( .DIN1(n12622), .DIN2(n12633), .Q(n10849) );
  nnd2s1 U12923 ( .DIN1(n12633), .DIN2(n12607), .Q(n10642) );
  nor2s1 U12924 ( .DIN1(n1521), .DIN2(n1403), .Q(n12607) );
  nnd2s1 U12925 ( .DIN1(n12631), .DIN2(n12620), .Q(n10646) );
  hi1s1 U12926 ( .DIN(n10832), .Q(n11113) );
  nnd3s1 U12927 ( .DIN1(sa12[1]), .DIN2(n1365), .DIN3(n12628), .Q(n10832) );
  nnd3s1 U12928 ( .DIN1(n12634), .DIN2(n12635), .DIN3(n12636), .Q(n12571) );
  nnd2s1 U12929 ( .DIN1(n10639), .DIN2(n10498), .Q(n12636) );
  hi1s1 U12930 ( .DIN(n10514), .Q(n10498) );
  hi1s1 U12931 ( .DIN(n11155), .Q(n10639) );
  nnd3s1 U12932 ( .DIN1(sa12[2]), .DIN2(n1365), .DIN3(n12637), .Q(n11155) );
  nnd2s1 U12933 ( .DIN1(n11567), .DIN2(n10497), .Q(n12635) );
  hi1s1 U12934 ( .DIN(n10518), .Q(n10497) );
  nnd3s1 U12935 ( .DIN1(sa12[1]), .DIN2(sa12[0]), .DIN3(n12628), .Q(n10518) );
  and2s1 U12936 ( .DIN1(sa12[3]), .DIN2(sa12[2]), .Q(n12628) );
  hi1s1 U12937 ( .DIN(n10641), .Q(n11567) );
  nnd2s1 U12938 ( .DIN1(n10810), .DIN2(n10628), .Q(n12634) );
  hi1s1 U12939 ( .DIN(n10817), .Q(n10628) );
  nnd2s1 U12940 ( .DIN1(n12631), .DIN2(n12633), .Q(n10817) );
  hi1s1 U12941 ( .DIN(n11497), .Q(n10810) );
  nnd4s1 U12942 ( .DIN1(n12638), .DIN2(n12639), .DIN3(n12640), .DIN4(n12641), 
        .Q(n12570) );
  nnd2s1 U12943 ( .DIN1(n11562), .DIN2(n12642), .Q(n12641) );
  nnd2s1 U12944 ( .DIN1(n11137), .DIN2(n10517), .Q(n12642) );
  nnd3s1 U12945 ( .DIN1(sa12[2]), .DIN2(sa12[0]), .DIN3(n12637), .Q(n10517) );
  hi1s1 U12946 ( .DIN(n11099), .Q(n11562) );
  nnd2s1 U12947 ( .DIN1(n12611), .DIN2(n12633), .Q(n11099) );
  and2s1 U12948 ( .DIN1(sa12[4]), .DIN2(sa12[6]), .Q(n12633) );
  nnd2s1 U12949 ( .DIN1(n11112), .DIN2(n12643), .Q(n12640) );
  nnd4s1 U12950 ( .DIN1(n11137), .DIN2(n11533), .DIN3(n11130), .DIN4(n11497), 
        .Q(n12643) );
  nnd3s1 U12951 ( .DIN1(sa12[0]), .DIN2(n12627), .DIN3(sa12[2]), .Q(n11497) );
  nnd3s1 U12952 ( .DIN1(n12600), .DIN2(sa12[0]), .DIN3(sa12[1]), .Q(n11130) );
  and2s1 U12953 ( .DIN1(sa12[3]), .DIN2(n1446), .Q(n12600) );
  nnd3s1 U12954 ( .DIN1(sa12[0]), .DIN2(n1446), .DIN3(n12637), .Q(n11533) );
  nnd3s1 U12955 ( .DIN1(n1365), .DIN2(n1446), .DIN3(n12627), .Q(n11137) );
  hi1s1 U12956 ( .DIN(n10645), .Q(n11112) );
  nnd2s1 U12957 ( .DIN1(n12611), .DIN2(n12621), .Q(n10645) );
  nnd2s1 U12958 ( .DIN1(n10850), .DIN2(n11537), .Q(n12639) );
  nnd2s1 U12959 ( .DIN1(n11504), .DIN2(n10514), .Q(n11537) );
  nnd2s1 U12960 ( .DIN1(n12622), .DIN2(n12620), .Q(n10514) );
  nnd2s1 U12961 ( .DIN1(n12611), .DIN2(n12620), .Q(n11504) );
  and2s1 U12962 ( .DIN1(sa12[6]), .DIN2(n1534), .Q(n12620) );
  nor2s1 U12963 ( .DIN1(sa12[7]), .DIN2(sa12[5]), .Q(n12611) );
  hi1s1 U12964 ( .DIN(n11133), .Q(n10850) );
  nnd3s1 U12965 ( .DIN1(n12627), .DIN2(n1365), .DIN3(sa12[2]), .Q(n11133) );
  nor2s1 U12966 ( .DIN1(sa12[3]), .DIN2(sa12[1]), .Q(n12627) );
  nnd2s1 U12967 ( .DIN1(n10499), .DIN2(n11122), .Q(n12638) );
  nnd2s1 U12968 ( .DIN1(n10632), .DIN2(n10641), .Q(n11122) );
  nnd2s1 U12969 ( .DIN1(n12621), .DIN2(n12631), .Q(n10641) );
  nor2s1 U12970 ( .DIN1(n1521), .DIN2(sa12[5]), .Q(n12631) );
  nor2s1 U12971 ( .DIN1(sa12[6]), .DIN2(sa12[4]), .Q(n12621) );
  nnd2s1 U12972 ( .DIN1(n12606), .DIN2(n12622), .Q(n10632) );
  nor2s1 U12973 ( .DIN1(n1403), .DIN2(sa12[7]), .Q(n12622) );
  nor2s1 U12974 ( .DIN1(n1534), .DIN2(sa12[6]), .Q(n12606) );
  hi1s1 U12975 ( .DIN(n11132), .Q(n10499) );
  nnd3s1 U12976 ( .DIN1(n1365), .DIN2(n1446), .DIN3(n12637), .Q(n11132) );
  nor2s1 U12977 ( .DIN1(n1433), .DIN2(sa12[3]), .Q(n12637) );
  hi1s1 U12978 ( .DIN(n12085), .Q(n5422) );
  or4s1 U12979 ( .DIN1(n12644), .DIN2(n12645), .DIN3(n12646), .DIN4(n12647), 
        .Q(n12085) );
  nnd4s1 U12980 ( .DIN1(n11162), .DIN2(n12648), .DIN3(n12649), .DIN4(n12650), 
        .Q(n12647) );
  nnd2s1 U12981 ( .DIN1(n10865), .DIN2(n11757), .Q(n12650) );
  nnd2s1 U12982 ( .DIN1(n11219), .DIN2(n11220), .Q(n11757) );
  nnd2s1 U12983 ( .DIN1(n10913), .DIN2(n11725), .Q(n12649) );
  nnd2s1 U12984 ( .DIN1(n10889), .DIN2(n11188), .Q(n11725) );
  nnd2s1 U12985 ( .DIN1(n11705), .DIN2(n10879), .Q(n12648) );
  nnd2s1 U12986 ( .DIN1(n10905), .DIN2(n11642), .Q(n11162) );
  nnd4s1 U12987 ( .DIN1(n12651), .DIN2(n12652), .DIN3(n12653), .DIN4(n12654), 
        .Q(n12646) );
  nnd2s1 U12988 ( .DIN1(n10685), .DIN2(n12655), .Q(n12654) );
  nnd2s1 U12989 ( .DIN1(n10680), .DIN2(n10874), .Q(n12655) );
  nnd2s1 U12990 ( .DIN1(n10877), .DIN2(n12656), .Q(n12653) );
  nnd2s1 U12991 ( .DIN1(n11225), .DIN2(n11215), .Q(n12656) );
  or2s1 U12992 ( .DIN1(n10912), .DIN2(n10891), .Q(n12652) );
  nor2s1 U12993 ( .DIN1(n10893), .DIN2(n10879), .Q(n10891) );
  nnd2s1 U12994 ( .DIN1(n11199), .DIN2(n10902), .Q(n12651) );
  nnd2s1 U12995 ( .DIN1(n10886), .DIN2(n10679), .Q(n10902) );
  nnd3s1 U12996 ( .DIN1(n11987), .DIN2(n12457), .DIN3(n12449), .Q(n12645) );
  nor4s1 U12997 ( .DIN1(n12657), .DIN2(n12658), .DIN3(n12659), .DIN4(n12660), 
        .Q(n12449) );
  nnd4s1 U12998 ( .DIN1(n12661), .DIN2(n12662), .DIN3(n12663), .DIN4(n12664), 
        .Q(n12660) );
  nnd2s1 U12999 ( .DIN1(n10672), .DIN2(n10662), .Q(n12664) );
  nor2s1 U13000 ( .DIN1(n12665), .DIN2(n11674), .Q(n12663) );
  nor2s1 U13001 ( .DIN1(n10889), .DIN2(n11704), .Q(n11674) );
  nor2s1 U13002 ( .DIN1(n10874), .DIN2(n10916), .Q(n12665) );
  nnd2s1 U13003 ( .DIN1(n10901), .DIN2(n11174), .Q(n12662) );
  nnd2s1 U13004 ( .DIN1(n10865), .DIN2(n10887), .Q(n12661) );
  hi1s1 U13005 ( .DIN(n11180), .Q(n10865) );
  nnd3s1 U13006 ( .DIN1(n12666), .DIN2(n12667), .DIN3(n12668), .Q(n12659) );
  nnd2s1 U13007 ( .DIN1(n10879), .DIN2(n11206), .Q(n12668) );
  nnd2s1 U13008 ( .DIN1(n10886), .DIN2(n10874), .Q(n11206) );
  nnd2s1 U13009 ( .DIN1(n11642), .DIN2(n12669), .Q(n12667) );
  nnd3s1 U13010 ( .DIN1(n11216), .DIN2(n11638), .DIN3(n11225), .Q(n12669) );
  nnd2s1 U13011 ( .DIN1(n10876), .DIN2(n12670), .Q(n12666) );
  nnd3s1 U13012 ( .DIN1(n11218), .DIN2(n11637), .DIN3(n11186), .Q(n12670) );
  nor2s1 U13013 ( .DIN1(n11186), .DIN2(n10895), .Q(n12658) );
  nor2s1 U13014 ( .DIN1(n11747), .DIN2(n11185), .Q(n12657) );
  nor2s1 U13015 ( .DIN1(n10677), .DIN2(n10910), .Q(n11747) );
  and4s1 U13016 ( .DIN1(n12671), .DIN2(n12672), .DIN3(n12673), .DIN4(n12674), 
        .Q(n12457) );
  and4s1 U13017 ( .DIN1(n12675), .DIN2(n11688), .DIN3(n12676), .DIN4(n12677), 
        .Q(n12674) );
  nnd2s1 U13018 ( .DIN1(n10905), .DIN2(n11705), .Q(n12677) );
  nnd2s1 U13019 ( .DIN1(n10662), .DIN2(n10664), .Q(n12676) );
  nnd2s1 U13020 ( .DIN1(n10893), .DIN2(n11710), .Q(n11688) );
  nnd2s1 U13021 ( .DIN1(n10685), .DIN2(n10672), .Q(n12675) );
  and3s1 U13022 ( .DIN1(n12678), .DIN2(n12679), .DIN3(n12680), .Q(n12673) );
  nnd2s1 U13023 ( .DIN1(n10901), .DIN2(n12681), .Q(n12680) );
  nnd2s1 U13024 ( .DIN1(n10684), .DIN2(n10886), .Q(n12681) );
  nnd2s1 U13025 ( .DIN1(n10663), .DIN2(n12682), .Q(n12679) );
  nnd2s1 U13026 ( .DIN1(n11180), .DIN2(n10684), .Q(n12682) );
  nnd2s1 U13027 ( .DIN1(n10866), .DIN2(n11739), .Q(n12678) );
  nnd2s1 U13028 ( .DIN1(n10889), .DIN2(n10912), .Q(n11739) );
  nnd2s1 U13029 ( .DIN1(n10681), .DIN2(n12683), .Q(n12672) );
  nnd3s1 U13030 ( .DIN1(n10912), .DIN2(n10683), .DIN3(n10670), .Q(n12683) );
  hi1s1 U13031 ( .DIN(n11704), .Q(n10681) );
  or2s1 U13032 ( .DIN1(n10886), .DIN2(n12499), .Q(n12671) );
  nor2s1 U13033 ( .DIN1(n10884), .DIN2(n10910), .Q(n12499) );
  nor4s1 U13034 ( .DIN1(n12684), .DIN2(n12685), .DIN3(n12686), .DIN4(n12687), 
        .Q(n11987) );
  nnd4s1 U13035 ( .DIN1(n12688), .DIN2(n12689), .DIN3(n12690), .DIN4(n12691), 
        .Q(n12687) );
  nor2s1 U13036 ( .DIN1(n12692), .DIN2(n12693), .Q(n12691) );
  nor2s1 U13037 ( .DIN1(n11216), .DIN2(n10679), .Q(n12693) );
  nor2s1 U13038 ( .DIN1(n11218), .DIN2(n10684), .Q(n12692) );
  nnd2s1 U13039 ( .DIN1(n10887), .DIN2(n11173), .Q(n12690) );
  or2s1 U13040 ( .DIN1(n11675), .DIN2(n11179), .Q(n12689) );
  nor2s1 U13041 ( .DIN1(n10672), .DIN2(n11173), .Q(n11179) );
  nnd2s1 U13042 ( .DIN1(n10904), .DIN2(n11172), .Q(n12688) );
  nnd3s1 U13043 ( .DIN1(n12694), .DIN2(n12695), .DIN3(n12696), .Q(n12686) );
  nnd2s1 U13044 ( .DIN1(n10663), .DIN2(n11241), .Q(n12696) );
  nnd2s1 U13045 ( .DIN1(n10679), .DIN2(n11188), .Q(n11241) );
  hi1s1 U13046 ( .DIN(n10916), .Q(n10663) );
  nnd2s1 U13047 ( .DIN1(n10664), .DIN2(n12697), .Q(n12695) );
  nnd2s1 U13048 ( .DIN1(n11637), .DIN2(n10892), .Q(n12697) );
  nnd2s1 U13049 ( .DIN1(n10876), .DIN2(n12698), .Q(n12694) );
  nnd2s1 U13050 ( .DIN1(n10917), .DIN2(n11675), .Q(n12698) );
  nor2s1 U13051 ( .DIN1(n12699), .DIN2(n10670), .Q(n12685) );
  nor2s1 U13052 ( .DIN1(n10685), .DIN2(n10866), .Q(n12699) );
  nor2s1 U13053 ( .DIN1(n12700), .DIN2(n10668), .Q(n12684) );
  nor2s1 U13054 ( .DIN1(n11172), .DIN2(n10677), .Q(n12700) );
  nnd4s1 U13055 ( .DIN1(n12149), .DIN2(n12701), .DIN3(n12702), .DIN4(n12703), 
        .Q(n12644) );
  nnd2s1 U13056 ( .DIN1(n10904), .DIN2(n10887), .Q(n12703) );
  nnd2s1 U13057 ( .DIN1(n10866), .DIN2(n10672), .Q(n12702) );
  nnd2s1 U13058 ( .DIN1(n11198), .DIN2(n10901), .Q(n12701) );
  nor3s1 U13059 ( .DIN1(n12704), .DIN2(n12705), .DIN3(n12706), .Q(n12149) );
  nnd4s1 U13060 ( .DIN1(n12451), .DIN2(n12458), .DIN3(n11992), .DIN4(n12707), 
        .Q(n12706) );
  and3s1 U13061 ( .DIN1(n12708), .DIN2(n12709), .DIN3(n12710), .Q(n12707) );
  nnd2s1 U13062 ( .DIN1(n10877), .DIN2(n10901), .Q(n12710) );
  nnd2s1 U13063 ( .DIN1(n10867), .DIN2(n10887), .Q(n12709) );
  hi1s1 U13064 ( .DIN(n11215), .Q(n10887) );
  hi1s1 U13065 ( .DIN(n10684), .Q(n10867) );
  nnd2s1 U13066 ( .DIN1(n11199), .DIN2(n11242), .Q(n12708) );
  hi1s1 U13067 ( .DIN(n10895), .Q(n11242) );
  and4s1 U13068 ( .DIN1(n12711), .DIN2(n12712), .DIN3(n12713), .DIN4(n12714), 
        .Q(n11992) );
  and4s1 U13069 ( .DIN1(n12715), .DIN2(n12716), .DIN3(n11653), .DIN4(n11170), 
        .Q(n12714) );
  nnd2s1 U13070 ( .DIN1(n10884), .DIN2(n10664), .Q(n11170) );
  nnd2s1 U13071 ( .DIN1(n10866), .DIN2(n10904), .Q(n11653) );
  nnd2s1 U13072 ( .DIN1(n10677), .DIN2(n10672), .Q(n12716) );
  nnd2s1 U13073 ( .DIN1(n10877), .DIN2(n11199), .Q(n12715) );
  and3s1 U13074 ( .DIN1(n12717), .DIN2(n12718), .DIN3(n12719), .Q(n12713) );
  nnd2s1 U13075 ( .DIN1(n10878), .DIN2(n12163), .Q(n12719) );
  nnd2s1 U13076 ( .DIN1(n11184), .DIN2(n10916), .Q(n12163) );
  nnd2s1 U13077 ( .DIN1(n10662), .DIN2(n12720), .Q(n12718) );
  nnd2s1 U13078 ( .DIN1(n11682), .DIN2(n10895), .Q(n12720) );
  nor2s1 U13079 ( .DIN1(n11198), .DIN2(n11173), .Q(n11682) );
  hi1s1 U13080 ( .DIN(n10889), .Q(n11173) );
  nnd2s1 U13081 ( .DIN1(n11710), .DIN2(n12721), .Q(n12717) );
  nnd2s1 U13082 ( .DIN1(n11219), .DIN2(n11704), .Q(n12721) );
  nnd2s1 U13083 ( .DIN1(n11198), .DIN2(n12722), .Q(n12712) );
  nnd2s1 U13084 ( .DIN1(n11244), .DIN2(n10917), .Q(n12722) );
  nnd2s1 U13085 ( .DIN1(n10879), .DIN2(n12723), .Q(n12711) );
  nnd3s1 U13086 ( .DIN1(n10680), .DIN2(n10670), .DIN3(n10684), .Q(n12723) );
  and4s1 U13087 ( .DIN1(n12724), .DIN2(n12725), .DIN3(n12726), .DIN4(n12727), 
        .Q(n12458) );
  nor4s1 U13088 ( .DIN1(n12728), .DIN2(n12729), .DIN3(n12730), .DIN4(n12731), 
        .Q(n12727) );
  nor2s1 U13089 ( .DIN1(n12732), .DIN2(n10679), .Q(n12731) );
  nor2s1 U13090 ( .DIN1(n10866), .DIN2(n10901), .Q(n12732) );
  nor2s1 U13091 ( .DIN1(n12733), .DIN2(n11188), .Q(n12730) );
  nor2s1 U13092 ( .DIN1(n11172), .DIN2(n10884), .Q(n12733) );
  hi1s1 U13093 ( .DIN(n10917), .Q(n10884) );
  nnd3s1 U13094 ( .DIN1(n12734), .DIN2(n1366), .DIN3(sa01[1]), .Q(n10917) );
  nor2s1 U13095 ( .DIN1(n12735), .DIN2(n10916), .Q(n12729) );
  nor2s1 U13096 ( .DIN1(n10661), .DIN2(n11198), .Q(n12735) );
  nnd3s1 U13097 ( .DIN1(n12736), .DIN2(n12737), .DIN3(n12738), .Q(n12728) );
  nnd2s1 U13098 ( .DIN1(n11172), .DIN2(n11705), .Q(n12738) );
  nnd2s1 U13099 ( .DIN1(n11174), .DIN2(n12739), .Q(n12737) );
  nnd2s1 U13100 ( .DIN1(n10892), .DIN2(n11186), .Q(n12739) );
  nnd2s1 U13101 ( .DIN1(n10893), .DIN2(n12003), .Q(n12736) );
  nnd2s1 U13102 ( .DIN1(n10886), .DIN2(n10889), .Q(n12003) );
  nnd2s1 U13103 ( .DIN1(n12740), .DIN2(n12741), .Q(n10889) );
  hi1s1 U13104 ( .DIN(n11225), .Q(n10893) );
  and3s1 U13105 ( .DIN1(n12742), .DIN2(n12743), .DIN3(n12744), .Q(n12726) );
  nnd2s1 U13106 ( .DIN1(n10913), .DIN2(n10876), .Q(n12744) );
  hi1s1 U13107 ( .DIN(n10680), .Q(n10876) );
  nnd2s1 U13108 ( .DIN1(n10661), .DIN2(n10905), .Q(n12743) );
  nnd2s1 U13109 ( .DIN1(n10878), .DIN2(n10910), .Q(n12742) );
  nnd2s1 U13110 ( .DIN1(n10677), .DIN2(n10904), .Q(n12725) );
  nnd2s1 U13111 ( .DIN1(n10672), .DIN2(n10879), .Q(n12724) );
  hi1s1 U13112 ( .DIN(n11216), .Q(n10879) );
  hi1s1 U13113 ( .DIN(n11699), .Q(n10672) );
  nnd2s1 U13114 ( .DIN1(n12740), .DIN2(n12745), .Q(n11699) );
  nor4s1 U13115 ( .DIN1(n12746), .DIN2(n12747), .DIN3(n12748), .DIN4(n12749), 
        .Q(n12451) );
  nnd4s1 U13116 ( .DIN1(n12750), .DIN2(n12751), .DIN3(n12752), .DIN4(n12753), 
        .Q(n12749) );
  nnd2s1 U13117 ( .DIN1(n10905), .DIN2(n11174), .Q(n12753) );
  hi1s1 U13118 ( .DIN(n11675), .Q(n10905) );
  nnd2s1 U13119 ( .DIN1(n10685), .DIN2(n11642), .Q(n12752) );
  hi1s1 U13120 ( .DIN(n11188), .Q(n11642) );
  nnd2s1 U13121 ( .DIN1(n12754), .DIN2(n12741), .Q(n11188) );
  hi1s1 U13122 ( .DIN(n11184), .Q(n10685) );
  nnd3s1 U13123 ( .DIN1(n1366), .DIN2(n1434), .DIN3(n12734), .Q(n11184) );
  nnd2s1 U13124 ( .DIN1(n10661), .DIN2(n10910), .Q(n12751) );
  hi1s1 U13125 ( .DIN(n11186), .Q(n10910) );
  hi1s1 U13126 ( .DIN(n10912), .Q(n10661) );
  nnd2s1 U13127 ( .DIN1(n10904), .DIN2(n10662), .Q(n12750) );
  hi1s1 U13128 ( .DIN(n10886), .Q(n10904) );
  nnd2s1 U13129 ( .DIN1(n12755), .DIN2(n12756), .Q(n10886) );
  nnd3s1 U13130 ( .DIN1(n12757), .DIN2(n12758), .DIN3(n12759), .Q(n12748) );
  nnd2s1 U13131 ( .DIN1(n10877), .DIN2(n12760), .Q(n12759) );
  nnd3s1 U13132 ( .DIN1(n10916), .DIN2(n11216), .DIN3(n11186), .Q(n12760) );
  nnd3s1 U13133 ( .DIN1(n12761), .DIN2(n1447), .DIN3(sa01[0]), .Q(n11186) );
  nnd3s1 U13134 ( .DIN1(sa01[0]), .DIN2(n1434), .DIN3(n12762), .Q(n10916) );
  hi1s1 U13135 ( .DIN(n11646), .Q(n10877) );
  nnd2s1 U13136 ( .DIN1(n10878), .DIN2(n12763), .Q(n12758) );
  nnd2s1 U13137 ( .DIN1(n11215), .DIN2(n11675), .Q(n12763) );
  nnd3s1 U13138 ( .DIN1(n1366), .DIN2(n1434), .DIN3(n12762), .Q(n11215) );
  hi1s1 U13139 ( .DIN(n10668), .Q(n10878) );
  nnd2s1 U13140 ( .DIN1(n10901), .DIN2(n12764), .Q(n12757) );
  nnd2s1 U13141 ( .DIN1(n11180), .DIN2(n11185), .Q(n12764) );
  nnd2s1 U13142 ( .DIN1(n12755), .DIN2(n12741), .Q(n11180) );
  hi1s1 U13143 ( .DIN(n11637), .Q(n10901) );
  nnd3s1 U13144 ( .DIN1(sa01[0]), .DIN2(n1434), .DIN3(n12734), .Q(n11637) );
  nor2s1 U13145 ( .DIN1(n10895), .DIN2(n11220), .Q(n12747) );
  nnd2s1 U13146 ( .DIN1(n12740), .DIN2(n12765), .Q(n10895) );
  and2s1 U13147 ( .DIN1(n11199), .DIN2(n12766), .Q(n12746) );
  nnd4s1 U13148 ( .DIN1(n10684), .DIN2(n10680), .DIN3(n10912), .DIN4(n10683), 
        .Q(n12766) );
  nnd2s1 U13149 ( .DIN1(n12756), .DIN2(n12767), .Q(n10912) );
  nnd2s1 U13150 ( .DIN1(n12767), .DIN2(n12741), .Q(n10680) );
  nor2s1 U13151 ( .DIN1(n1522), .DIN2(n1404), .Q(n12741) );
  nnd2s1 U13152 ( .DIN1(n12765), .DIN2(n12754), .Q(n10684) );
  hi1s1 U13153 ( .DIN(n10892), .Q(n11199) );
  nnd3s1 U13154 ( .DIN1(sa01[1]), .DIN2(n1366), .DIN3(n12762), .Q(n10892) );
  nnd3s1 U13155 ( .DIN1(n12768), .DIN2(n12769), .DIN3(n12770), .Q(n12705) );
  nnd2s1 U13156 ( .DIN1(n10677), .DIN2(n11174), .Q(n12770) );
  hi1s1 U13157 ( .DIN(n10670), .Q(n11174) );
  hi1s1 U13158 ( .DIN(n11244), .Q(n10677) );
  nnd3s1 U13159 ( .DIN1(sa01[2]), .DIN2(n1366), .DIN3(n12771), .Q(n11244) );
  nnd2s1 U13160 ( .DIN1(n11710), .DIN2(n11172), .Q(n12769) );
  hi1s1 U13161 ( .DIN(n11220), .Q(n11172) );
  nnd3s1 U13162 ( .DIN1(sa01[1]), .DIN2(sa01[0]), .DIN3(n12762), .Q(n11220) );
  and2s1 U13163 ( .DIN1(sa01[3]), .DIN2(sa01[2]), .Q(n12762) );
  hi1s1 U13164 ( .DIN(n10679), .Q(n11710) );
  nnd2s1 U13165 ( .DIN1(n10866), .DIN2(n10664), .Q(n12768) );
  hi1s1 U13166 ( .DIN(n10874), .Q(n10664) );
  nnd2s1 U13167 ( .DIN1(n12765), .DIN2(n12767), .Q(n10874) );
  hi1s1 U13168 ( .DIN(n11638), .Q(n10866) );
  nnd4s1 U13169 ( .DIN1(n12772), .DIN2(n12773), .DIN3(n12774), .DIN4(n12775), 
        .Q(n12704) );
  nnd2s1 U13170 ( .DIN1(n11705), .DIN2(n12776), .Q(n12775) );
  nnd2s1 U13171 ( .DIN1(n11225), .DIN2(n11704), .Q(n12776) );
  nnd3s1 U13172 ( .DIN1(sa01[2]), .DIN2(sa01[0]), .DIN3(n12771), .Q(n11704) );
  hi1s1 U13173 ( .DIN(n11185), .Q(n11705) );
  nnd2s1 U13174 ( .DIN1(n12745), .DIN2(n12767), .Q(n11185) );
  and2s1 U13175 ( .DIN1(sa01[4]), .DIN2(sa01[6]), .Q(n12767) );
  nnd2s1 U13176 ( .DIN1(n11198), .DIN2(n12777), .Q(n12774) );
  nnd4s1 U13177 ( .DIN1(n11225), .DIN2(n11675), .DIN3(n11216), .DIN4(n11638), 
        .Q(n12777) );
  nnd3s1 U13178 ( .DIN1(sa01[0]), .DIN2(n12761), .DIN3(sa01[2]), .Q(n11638) );
  nnd3s1 U13179 ( .DIN1(n12734), .DIN2(sa01[0]), .DIN3(sa01[1]), .Q(n11216) );
  and2s1 U13180 ( .DIN1(sa01[3]), .DIN2(n1447), .Q(n12734) );
  nnd3s1 U13181 ( .DIN1(sa01[0]), .DIN2(n1447), .DIN3(n12771), .Q(n11675) );
  nnd3s1 U13182 ( .DIN1(n1366), .DIN2(n1447), .DIN3(n12761), .Q(n11225) );
  hi1s1 U13183 ( .DIN(n10683), .Q(n11198) );
  nnd2s1 U13184 ( .DIN1(n12745), .DIN2(n12755), .Q(n10683) );
  nnd2s1 U13185 ( .DIN1(n10913), .DIN2(n11679), .Q(n12773) );
  nnd2s1 U13186 ( .DIN1(n11646), .DIN2(n10670), .Q(n11679) );
  nnd2s1 U13187 ( .DIN1(n12756), .DIN2(n12754), .Q(n10670) );
  nnd2s1 U13188 ( .DIN1(n12745), .DIN2(n12754), .Q(n11646) );
  and2s1 U13189 ( .DIN1(sa01[6]), .DIN2(n1535), .Q(n12754) );
  nor2s1 U13190 ( .DIN1(sa01[7]), .DIN2(sa01[5]), .Q(n12745) );
  hi1s1 U13191 ( .DIN(n11219), .Q(n10913) );
  nnd3s1 U13192 ( .DIN1(n12761), .DIN2(n1366), .DIN3(sa01[2]), .Q(n11219) );
  nor2s1 U13193 ( .DIN1(sa01[3]), .DIN2(sa01[1]), .Q(n12761) );
  nnd2s1 U13194 ( .DIN1(n10662), .DIN2(n11208), .Q(n12772) );
  nnd2s1 U13195 ( .DIN1(n10668), .DIN2(n10679), .Q(n11208) );
  nnd2s1 U13196 ( .DIN1(n12755), .DIN2(n12765), .Q(n10679) );
  nor2s1 U13197 ( .DIN1(n1522), .DIN2(sa01[5]), .Q(n12765) );
  nor2s1 U13198 ( .DIN1(sa01[6]), .DIN2(sa01[4]), .Q(n12755) );
  nnd2s1 U13199 ( .DIN1(n12740), .DIN2(n12756), .Q(n10668) );
  nor2s1 U13200 ( .DIN1(n1404), .DIN2(sa01[7]), .Q(n12756) );
  nor2s1 U13201 ( .DIN1(n1535), .DIN2(sa01[6]), .Q(n12740) );
  hi1s1 U13202 ( .DIN(n11218), .Q(n10662) );
  nnd3s1 U13203 ( .DIN1(n1366), .DIN2(n1447), .DIN3(n12771), .Q(n11218) );
  nor2s1 U13204 ( .DIN1(n1434), .DIN2(sa01[3]), .Q(n12771) );
  xor2s1 U13205 ( .DIN1(n1497), .DIN2(n5045), .Q(n12310) );
  nor4s1 U13206 ( .DIN1(n12778), .DIN2(n12779), .DIN3(n12780), .DIN4(n12781), 
        .Q(n5045) );
  nnd4s1 U13207 ( .DIN1(n11394), .DIN2(n12782), .DIN3(n12783), .DIN4(n12784), 
        .Q(n12781) );
  nnd2s1 U13208 ( .DIN1(n11019), .DIN2(n11921), .Q(n12784) );
  nnd2s1 U13209 ( .DIN1(n11448), .DIN2(n10599), .Q(n11921) );
  nnd2s1 U13210 ( .DIN1(n11060), .DIN2(n10601), .Q(n12783) );
  nnd2s1 U13211 ( .DIN1(n11039), .DIN2(n11417), .Q(n10601) );
  nnd2s1 U13212 ( .DIN1(n11870), .DIN2(n11030), .Q(n12782) );
  nnd2s1 U13213 ( .DIN1(n11053), .DIN2(n10581), .Q(n11394) );
  nnd4s1 U13214 ( .DIN1(n12785), .DIN2(n12786), .DIN3(n12787), .DIN4(n12788), 
        .Q(n12780) );
  nnd2s1 U13215 ( .DIN1(n10572), .DIN2(n12789), .Q(n12788) );
  nnd2s1 U13216 ( .DIN1(n10785), .DIN2(n11027), .Q(n12789) );
  nnd2s1 U13217 ( .DIN1(n11018), .DIN2(n12790), .Q(n12787) );
  nnd2s1 U13218 ( .DIN1(n11452), .DIN2(n11444), .Q(n12790) );
  or2s1 U13219 ( .DIN1(n11059), .DIN2(n11041), .Q(n12786) );
  nor2s1 U13220 ( .DIN1(n10592), .DIN2(n11030), .Q(n11041) );
  nnd2s1 U13221 ( .DIN1(n11428), .DIN2(n11051), .Q(n12785) );
  nnd2s1 U13222 ( .DIN1(n11036), .DIN2(n10784), .Q(n11051) );
  nnd3s1 U13223 ( .DIN1(n12044), .DIN2(n12052), .DIN3(n10563), .Q(n12779) );
  nor4s1 U13224 ( .DIN1(n12791), .DIN2(n12792), .DIN3(n12793), .DIN4(n12794), 
        .Q(n10563) );
  nnd4s1 U13225 ( .DIN1(n12795), .DIN2(n12796), .DIN3(n12797), .DIN4(n12798), 
        .Q(n12794) );
  nnd2s1 U13226 ( .DIN1(n10596), .DIN2(n10580), .Q(n12798) );
  nor2s1 U13227 ( .DIN1(n12799), .DIN2(n11840), .Q(n12797) );
  nor2s1 U13228 ( .DIN1(n11039), .DIN2(n10598), .Q(n11840) );
  nor2s1 U13229 ( .DIN1(n11027), .DIN2(n11063), .Q(n12799) );
  nnd2s1 U13230 ( .DIN1(n11050), .DIN2(n10579), .Q(n12796) );
  nnd2s1 U13231 ( .DIN1(n11019), .DIN2(n11037), .Q(n12795) );
  hi1s1 U13232 ( .DIN(n10594), .Q(n11019) );
  nnd3s1 U13233 ( .DIN1(n12800), .DIN2(n12801), .DIN3(n12802), .Q(n12793) );
  nnd2s1 U13234 ( .DIN1(n11030), .DIN2(n11435), .Q(n12802) );
  nnd2s1 U13235 ( .DIN1(n11036), .DIN2(n11027), .Q(n11435) );
  nnd2s1 U13236 ( .DIN1(n10581), .DIN2(n12803), .Q(n12801) );
  nnd3s1 U13237 ( .DIN1(n11445), .DIN2(n11805), .DIN3(n11452), .Q(n12803) );
  nnd2s1 U13238 ( .DIN1(n11029), .DIN2(n12804), .Q(n12800) );
  nnd3s1 U13239 ( .DIN1(n11447), .DIN2(n11804), .DIN3(n11415), .Q(n12804) );
  nor2s1 U13240 ( .DIN1(n11415), .DIN2(n11044), .Q(n12792) );
  nor2s1 U13241 ( .DIN1(n11911), .DIN2(n11414), .Q(n12791) );
  nor2s1 U13242 ( .DIN1(n10782), .DIN2(n10600), .Q(n11911) );
  and4s1 U13243 ( .DIN1(n12805), .DIN2(n12806), .DIN3(n12807), .DIN4(n12808), 
        .Q(n12052) );
  and4s1 U13244 ( .DIN1(n12809), .DIN2(n11854), .DIN3(n12810), .DIN4(n12811), 
        .Q(n12808) );
  nnd2s1 U13245 ( .DIN1(n11053), .DIN2(n11870), .Q(n12811) );
  nnd2s1 U13246 ( .DIN1(n10580), .DIN2(n10771), .Q(n12810) );
  nnd2s1 U13247 ( .DIN1(n10592), .DIN2(n11875), .Q(n11854) );
  nnd2s1 U13248 ( .DIN1(n10572), .DIN2(n10596), .Q(n12809) );
  and3s1 U13249 ( .DIN1(n12812), .DIN2(n12813), .DIN3(n12814), .Q(n12807) );
  nnd2s1 U13250 ( .DIN1(n11050), .DIN2(n12815), .Q(n12814) );
  nnd2s1 U13251 ( .DIN1(n10789), .DIN2(n11036), .Q(n12815) );
  nnd2s1 U13252 ( .DIN1(n10571), .DIN2(n12816), .Q(n12813) );
  nnd2s1 U13253 ( .DIN1(n10594), .DIN2(n10789), .Q(n12816) );
  nnd2s1 U13254 ( .DIN1(n11020), .DIN2(n11903), .Q(n12812) );
  nnd2s1 U13255 ( .DIN1(n11039), .DIN2(n11059), .Q(n11903) );
  nnd2s1 U13256 ( .DIN1(n10786), .DIN2(n12817), .Q(n12806) );
  nnd3s1 U13257 ( .DIN1(n11059), .DIN2(n10788), .DIN3(n10595), .Q(n12817) );
  hi1s1 U13258 ( .DIN(n10598), .Q(n10786) );
  or2s1 U13259 ( .DIN1(n11036), .DIN2(n12294), .Q(n12805) );
  nor2s1 U13260 ( .DIN1(n10582), .DIN2(n10600), .Q(n12294) );
  nor4s1 U13261 ( .DIN1(n12818), .DIN2(n12819), .DIN3(n12820), .DIN4(n12821), 
        .Q(n12044) );
  nnd4s1 U13262 ( .DIN1(n12822), .DIN2(n12823), .DIN3(n12824), .DIN4(n12825), 
        .Q(n12821) );
  nor2s1 U13263 ( .DIN1(n12826), .DIN2(n12827), .Q(n12825) );
  nor2s1 U13264 ( .DIN1(n11445), .DIN2(n10784), .Q(n12827) );
  nor2s1 U13265 ( .DIN1(n11447), .DIN2(n10789), .Q(n12826) );
  nnd2s1 U13266 ( .DIN1(n11037), .DIN2(n11404), .Q(n12824) );
  or2s1 U13267 ( .DIN1(n11841), .DIN2(n11409), .Q(n12823) );
  nor2s1 U13268 ( .DIN1(n10596), .DIN2(n11404), .Q(n11409) );
  nnd2s1 U13269 ( .DIN1(n10570), .DIN2(n10578), .Q(n12822) );
  nnd3s1 U13270 ( .DIN1(n12828), .DIN2(n12829), .DIN3(n12830), .Q(n12820) );
  nnd2s1 U13271 ( .DIN1(n10571), .DIN2(n11468), .Q(n12830) );
  nnd2s1 U13272 ( .DIN1(n10784), .DIN2(n11417), .Q(n11468) );
  hi1s1 U13273 ( .DIN(n11063), .Q(n10571) );
  nnd2s1 U13274 ( .DIN1(n10771), .DIN2(n12831), .Q(n12829) );
  nnd2s1 U13275 ( .DIN1(n11804), .DIN2(n11042), .Q(n12831) );
  nnd2s1 U13276 ( .DIN1(n11029), .DIN2(n12832), .Q(n12828) );
  nnd2s1 U13277 ( .DIN1(n10591), .DIN2(n11841), .Q(n12832) );
  nor2s1 U13278 ( .DIN1(n12833), .DIN2(n10595), .Q(n12819) );
  nor2s1 U13279 ( .DIN1(n10572), .DIN2(n11020), .Q(n12833) );
  nor2s1 U13280 ( .DIN1(n12834), .DIN2(n10775), .Q(n12818) );
  nor2s1 U13281 ( .DIN1(n10578), .DIN2(n10782), .Q(n12834) );
  nnd4s1 U13282 ( .DIN1(n12251), .DIN2(n12835), .DIN3(n12836), .DIN4(n12837), 
        .Q(n12778) );
  nnd2s1 U13283 ( .DIN1(n10570), .DIN2(n11037), .Q(n12837) );
  nnd2s1 U13284 ( .DIN1(n11020), .DIN2(n10596), .Q(n12836) );
  nnd2s1 U13285 ( .DIN1(n11427), .DIN2(n11050), .Q(n12835) );
  nor3s1 U13286 ( .DIN1(n12838), .DIN2(n12839), .DIN3(n12840), .Q(n12251) );
  nnd4s1 U13287 ( .DIN1(n10566), .DIN2(n12053), .DIN3(n12048), .DIN4(n12841), 
        .Q(n12840) );
  and3s1 U13288 ( .DIN1(n12842), .DIN2(n12843), .DIN3(n12844), .Q(n12841) );
  nnd2s1 U13289 ( .DIN1(n11018), .DIN2(n11050), .Q(n12844) );
  nnd2s1 U13290 ( .DIN1(n10573), .DIN2(n11037), .Q(n12843) );
  hi1s1 U13291 ( .DIN(n11444), .Q(n11037) );
  hi1s1 U13292 ( .DIN(n10789), .Q(n10573) );
  nnd2s1 U13293 ( .DIN1(n11428), .DIN2(n10588), .Q(n12842) );
  hi1s1 U13294 ( .DIN(n11044), .Q(n10588) );
  and4s1 U13295 ( .DIN1(n12845), .DIN2(n12846), .DIN3(n12847), .DIN4(n12848), 
        .Q(n12048) );
  and4s1 U13296 ( .DIN1(n12849), .DIN2(n12850), .DIN3(n11819), .DIN4(n11402), 
        .Q(n12848) );
  nnd2s1 U13297 ( .DIN1(n10582), .DIN2(n10771), .Q(n11402) );
  nnd2s1 U13298 ( .DIN1(n11020), .DIN2(n10570), .Q(n11819) );
  nnd2s1 U13299 ( .DIN1(n10782), .DIN2(n10596), .Q(n12850) );
  nnd2s1 U13300 ( .DIN1(n11018), .DIN2(n11428), .Q(n12849) );
  and3s1 U13301 ( .DIN1(n12851), .DIN2(n12852), .DIN3(n12853), .Q(n12847) );
  nnd2s1 U13302 ( .DIN1(n10583), .DIN2(n12263), .Q(n12853) );
  nnd2s1 U13303 ( .DIN1(n11413), .DIN2(n11063), .Q(n12263) );
  nnd2s1 U13304 ( .DIN1(n10580), .DIN2(n12854), .Q(n12852) );
  nnd2s1 U13305 ( .DIN1(n11848), .DIN2(n11044), .Q(n12854) );
  nor2s1 U13306 ( .DIN1(n11427), .DIN2(n11404), .Q(n11848) );
  hi1s1 U13307 ( .DIN(n11039), .Q(n11404) );
  nnd2s1 U13308 ( .DIN1(n11875), .DIN2(n12855), .Q(n12851) );
  nnd2s1 U13309 ( .DIN1(n11448), .DIN2(n10598), .Q(n12855) );
  nnd2s1 U13310 ( .DIN1(n11427), .DIN2(n12856), .Q(n12846) );
  nnd2s1 U13311 ( .DIN1(n11470), .DIN2(n10591), .Q(n12856) );
  nnd2s1 U13312 ( .DIN1(n11030), .DIN2(n12857), .Q(n12845) );
  nnd3s1 U13313 ( .DIN1(n10785), .DIN2(n10595), .DIN3(n10789), .Q(n12857) );
  and4s1 U13314 ( .DIN1(n12858), .DIN2(n12859), .DIN3(n12860), .DIN4(n12861), 
        .Q(n12053) );
  nor4s1 U13315 ( .DIN1(n12862), .DIN2(n12863), .DIN3(n12864), .DIN4(n12865), 
        .Q(n12861) );
  nor2s1 U13316 ( .DIN1(n12866), .DIN2(n10784), .Q(n12865) );
  nor2s1 U13317 ( .DIN1(n11020), .DIN2(n11050), .Q(n12866) );
  nor2s1 U13318 ( .DIN1(n12867), .DIN2(n11417), .Q(n12864) );
  nor2s1 U13319 ( .DIN1(n10578), .DIN2(n10582), .Q(n12867) );
  hi1s1 U13320 ( .DIN(n10591), .Q(n10582) );
  nnd3s1 U13321 ( .DIN1(n12868), .DIN2(n1367), .DIN3(sa23[1]), .Q(n10591) );
  nor2s1 U13322 ( .DIN1(n12869), .DIN2(n11063), .Q(n12863) );
  nor2s1 U13323 ( .DIN1(n10770), .DIN2(n11427), .Q(n12869) );
  nnd3s1 U13324 ( .DIN1(n12870), .DIN2(n12871), .DIN3(n12872), .Q(n12862) );
  nnd2s1 U13325 ( .DIN1(n10578), .DIN2(n11870), .Q(n12872) );
  nnd2s1 U13326 ( .DIN1(n10579), .DIN2(n12873), .Q(n12871) );
  nnd2s1 U13327 ( .DIN1(n11042), .DIN2(n11415), .Q(n12873) );
  nnd2s1 U13328 ( .DIN1(n10592), .DIN2(n12078), .Q(n12870) );
  nnd2s1 U13329 ( .DIN1(n11036), .DIN2(n11039), .Q(n12078) );
  nnd2s1 U13330 ( .DIN1(n12874), .DIN2(n12875), .Q(n11039) );
  hi1s1 U13331 ( .DIN(n11452), .Q(n10592) );
  and3s1 U13332 ( .DIN1(n12876), .DIN2(n12877), .DIN3(n12878), .Q(n12860) );
  nnd2s1 U13333 ( .DIN1(n11060), .DIN2(n11029), .Q(n12878) );
  hi1s1 U13334 ( .DIN(n10785), .Q(n11029) );
  nnd2s1 U13335 ( .DIN1(n10770), .DIN2(n11053), .Q(n12877) );
  nnd2s1 U13336 ( .DIN1(n10583), .DIN2(n10600), .Q(n12876) );
  nnd2s1 U13337 ( .DIN1(n10782), .DIN2(n10570), .Q(n12859) );
  nnd2s1 U13338 ( .DIN1(n10596), .DIN2(n11030), .Q(n12858) );
  hi1s1 U13339 ( .DIN(n11445), .Q(n11030) );
  hi1s1 U13340 ( .DIN(n11865), .Q(n10596) );
  nnd2s1 U13341 ( .DIN1(n12874), .DIN2(n12879), .Q(n11865) );
  nor4s1 U13342 ( .DIN1(n12880), .DIN2(n12881), .DIN3(n12882), .DIN4(n12883), 
        .Q(n10566) );
  nnd4s1 U13343 ( .DIN1(n12884), .DIN2(n12885), .DIN3(n12886), .DIN4(n12887), 
        .Q(n12883) );
  nnd2s1 U13344 ( .DIN1(n11053), .DIN2(n10579), .Q(n12887) );
  hi1s1 U13345 ( .DIN(n11841), .Q(n11053) );
  nnd2s1 U13346 ( .DIN1(n10572), .DIN2(n10581), .Q(n12886) );
  hi1s1 U13347 ( .DIN(n11417), .Q(n10581) );
  nnd2s1 U13348 ( .DIN1(n12888), .DIN2(n12875), .Q(n11417) );
  hi1s1 U13349 ( .DIN(n11413), .Q(n10572) );
  nnd3s1 U13350 ( .DIN1(n1367), .DIN2(n1435), .DIN3(n12868), .Q(n11413) );
  nnd2s1 U13351 ( .DIN1(n10770), .DIN2(n10600), .Q(n12885) );
  hi1s1 U13352 ( .DIN(n11415), .Q(n10600) );
  hi1s1 U13353 ( .DIN(n11059), .Q(n10770) );
  nnd2s1 U13354 ( .DIN1(n10570), .DIN2(n10580), .Q(n12884) );
  hi1s1 U13355 ( .DIN(n11036), .Q(n10570) );
  nnd2s1 U13356 ( .DIN1(n12889), .DIN2(n12890), .Q(n11036) );
  nnd3s1 U13357 ( .DIN1(n12891), .DIN2(n12892), .DIN3(n12893), .Q(n12882) );
  nnd2s1 U13358 ( .DIN1(n11018), .DIN2(n12894), .Q(n12893) );
  nnd3s1 U13359 ( .DIN1(n11063), .DIN2(n11445), .DIN3(n11415), .Q(n12894) );
  nnd3s1 U13360 ( .DIN1(n12895), .DIN2(n1448), .DIN3(sa23[0]), .Q(n11415) );
  nnd3s1 U13361 ( .DIN1(sa23[0]), .DIN2(n1435), .DIN3(n12896), .Q(n11063) );
  hi1s1 U13362 ( .DIN(n11812), .Q(n11018) );
  nnd2s1 U13363 ( .DIN1(n10583), .DIN2(n12897), .Q(n12892) );
  nnd2s1 U13364 ( .DIN1(n11444), .DIN2(n11841), .Q(n12897) );
  nnd3s1 U13365 ( .DIN1(n1367), .DIN2(n1435), .DIN3(n12896), .Q(n11444) );
  hi1s1 U13366 ( .DIN(n10775), .Q(n10583) );
  nnd2s1 U13367 ( .DIN1(n11050), .DIN2(n12898), .Q(n12891) );
  nnd2s1 U13368 ( .DIN1(n10594), .DIN2(n11414), .Q(n12898) );
  nnd2s1 U13369 ( .DIN1(n12889), .DIN2(n12875), .Q(n10594) );
  hi1s1 U13370 ( .DIN(n11804), .Q(n11050) );
  nnd3s1 U13371 ( .DIN1(sa23[0]), .DIN2(n1435), .DIN3(n12868), .Q(n11804) );
  nor2s1 U13372 ( .DIN1(n11044), .DIN2(n10599), .Q(n12881) );
  nnd2s1 U13373 ( .DIN1(n12874), .DIN2(n12899), .Q(n11044) );
  and2s1 U13374 ( .DIN1(n11428), .DIN2(n12900), .Q(n12880) );
  nnd4s1 U13375 ( .DIN1(n10789), .DIN2(n10785), .DIN3(n11059), .DIN4(n10788), 
        .Q(n12900) );
  nnd2s1 U13376 ( .DIN1(n12890), .DIN2(n12901), .Q(n11059) );
  nnd2s1 U13377 ( .DIN1(n12901), .DIN2(n12875), .Q(n10785) );
  nor2s1 U13378 ( .DIN1(n1523), .DIN2(n1405), .Q(n12875) );
  nnd2s1 U13379 ( .DIN1(n12899), .DIN2(n12888), .Q(n10789) );
  hi1s1 U13380 ( .DIN(n11042), .Q(n11428) );
  nnd3s1 U13381 ( .DIN1(sa23[1]), .DIN2(n1367), .DIN3(n12896), .Q(n11042) );
  nnd3s1 U13382 ( .DIN1(n12902), .DIN2(n12903), .DIN3(n12904), .Q(n12839) );
  nnd2s1 U13383 ( .DIN1(n10782), .DIN2(n10579), .Q(n12904) );
  hi1s1 U13384 ( .DIN(n10595), .Q(n10579) );
  hi1s1 U13385 ( .DIN(n11470), .Q(n10782) );
  nnd3s1 U13386 ( .DIN1(sa23[2]), .DIN2(n1367), .DIN3(n12905), .Q(n11470) );
  nnd2s1 U13387 ( .DIN1(n11875), .DIN2(n10578), .Q(n12903) );
  hi1s1 U13388 ( .DIN(n10599), .Q(n10578) );
  nnd3s1 U13389 ( .DIN1(sa23[1]), .DIN2(sa23[0]), .DIN3(n12896), .Q(n10599) );
  and2s1 U13390 ( .DIN1(sa23[3]), .DIN2(sa23[2]), .Q(n12896) );
  hi1s1 U13391 ( .DIN(n10784), .Q(n11875) );
  nnd2s1 U13392 ( .DIN1(n11020), .DIN2(n10771), .Q(n12902) );
  hi1s1 U13393 ( .DIN(n11027), .Q(n10771) );
  nnd2s1 U13394 ( .DIN1(n12899), .DIN2(n12901), .Q(n11027) );
  hi1s1 U13395 ( .DIN(n11805), .Q(n11020) );
  nnd4s1 U13396 ( .DIN1(n12906), .DIN2(n12907), .DIN3(n12908), .DIN4(n12909), 
        .Q(n12838) );
  nnd2s1 U13397 ( .DIN1(n11870), .DIN2(n12910), .Q(n12909) );
  nnd2s1 U13398 ( .DIN1(n11452), .DIN2(n10598), .Q(n12910) );
  nnd3s1 U13399 ( .DIN1(sa23[2]), .DIN2(sa23[0]), .DIN3(n12905), .Q(n10598) );
  hi1s1 U13400 ( .DIN(n11414), .Q(n11870) );
  nnd2s1 U13401 ( .DIN1(n12879), .DIN2(n12901), .Q(n11414) );
  and2s1 U13402 ( .DIN1(sa23[4]), .DIN2(sa23[6]), .Q(n12901) );
  nnd2s1 U13403 ( .DIN1(n11427), .DIN2(n12911), .Q(n12908) );
  nnd4s1 U13404 ( .DIN1(n11452), .DIN2(n11841), .DIN3(n11445), .DIN4(n11805), 
        .Q(n12911) );
  nnd3s1 U13405 ( .DIN1(sa23[0]), .DIN2(n12895), .DIN3(sa23[2]), .Q(n11805) );
  nnd3s1 U13406 ( .DIN1(n12868), .DIN2(sa23[0]), .DIN3(sa23[1]), .Q(n11445) );
  and2s1 U13407 ( .DIN1(sa23[3]), .DIN2(n1448), .Q(n12868) );
  nnd3s1 U13408 ( .DIN1(sa23[0]), .DIN2(n1448), .DIN3(n12905), .Q(n11841) );
  nnd3s1 U13409 ( .DIN1(n1367), .DIN2(n1448), .DIN3(n12895), .Q(n11452) );
  hi1s1 U13410 ( .DIN(n10788), .Q(n11427) );
  nnd2s1 U13411 ( .DIN1(n12879), .DIN2(n12889), .Q(n10788) );
  nnd2s1 U13412 ( .DIN1(n11060), .DIN2(n11845), .Q(n12907) );
  nnd2s1 U13413 ( .DIN1(n11812), .DIN2(n10595), .Q(n11845) );
  nnd2s1 U13414 ( .DIN1(n12890), .DIN2(n12888), .Q(n10595) );
  nnd2s1 U13415 ( .DIN1(n12879), .DIN2(n12888), .Q(n11812) );
  and2s1 U13416 ( .DIN1(sa23[6]), .DIN2(n1536), .Q(n12888) );
  nor2s1 U13417 ( .DIN1(sa23[7]), .DIN2(sa23[5]), .Q(n12879) );
  hi1s1 U13418 ( .DIN(n11448), .Q(n11060) );
  nnd3s1 U13419 ( .DIN1(n12895), .DIN2(n1367), .DIN3(sa23[2]), .Q(n11448) );
  nor2s1 U13420 ( .DIN1(sa23[3]), .DIN2(sa23[1]), .Q(n12895) );
  nnd2s1 U13421 ( .DIN1(n10580), .DIN2(n11437), .Q(n12906) );
  nnd2s1 U13422 ( .DIN1(n10775), .DIN2(n10784), .Q(n11437) );
  nnd2s1 U13423 ( .DIN1(n12889), .DIN2(n12899), .Q(n10784) );
  nor2s1 U13424 ( .DIN1(n1523), .DIN2(sa23[5]), .Q(n12899) );
  nor2s1 U13425 ( .DIN1(sa23[6]), .DIN2(sa23[4]), .Q(n12889) );
  nnd2s1 U13426 ( .DIN1(n12874), .DIN2(n12890), .Q(n10775) );
  nor2s1 U13427 ( .DIN1(n1405), .DIN2(sa23[7]), .Q(n12890) );
  nor2s1 U13428 ( .DIN1(n1536), .DIN2(sa23[6]), .Q(n12874) );
  hi1s1 U13429 ( .DIN(n11447), .Q(n10580) );
  nnd3s1 U13430 ( .DIN1(n1367), .DIN2(n1448), .DIN3(n12905), .Q(n11447) );
  nor2s1 U13431 ( .DIN1(n1435), .DIN2(sa23[3]), .Q(n12905) );
  nnd2s1 U13432 ( .DIN1(n12912), .DIN2(n1601), .Q(n12307) );
  xor2s1 U13433 ( .DIN1(w1[0]), .DIN2(text_in_r[64]), .Q(n12912) );
  nnd2s1 U13434 ( .DIN1(n12913), .DIN2(n12914), .Q(N153) );
  nnd2s1 U13435 ( .DIN1(n12915), .DIN2(n1632), .Q(n12914) );
  xor2s1 U13436 ( .DIN1(n12916), .DIN2(n12917), .Q(n12915) );
  xor2s1 U13437 ( .DIN1(n12918), .DIN2(n12919), .Q(n12917) );
  xor2s1 U13438 ( .DIN1(n1451), .DIN2(n12920), .Q(n12916) );
  hi1s1 U13439 ( .DIN(n5068), .Q(n12920) );
  nnd2s1 U13440 ( .DIN1(n12921), .DIN2(n1600), .Q(n12913) );
  xor2s1 U13441 ( .DIN1(w2[31]), .DIN2(text_in_r[63]), .Q(n12921) );
  nnd2s1 U13442 ( .DIN1(n12922), .DIN2(n12923), .Q(N152) );
  nnd2s1 U13443 ( .DIN1(n12924), .DIN2(n1633), .Q(n12923) );
  xor2s1 U13444 ( .DIN1(n12925), .DIN2(n12926), .Q(n12924) );
  xor2s1 U13445 ( .DIN1(n12927), .DIN2(n12928), .Q(n12926) );
  xor2s1 U13446 ( .DIN1(n5067), .DIN2(w2[30]), .Q(n12925) );
  nnd2s1 U13447 ( .DIN1(n12929), .DIN2(n1600), .Q(n12922) );
  xor2s1 U13448 ( .DIN1(w2[30]), .DIN2(text_in_r[62]), .Q(n12929) );
  nnd2s1 U13449 ( .DIN1(n12930), .DIN2(n12931), .Q(N151) );
  nnd2s1 U13450 ( .DIN1(n12932), .DIN2(n1632), .Q(n12931) );
  xor2s1 U13451 ( .DIN1(n12933), .DIN2(n12934), .Q(n12932) );
  xor2s1 U13452 ( .DIN1(n12935), .DIN2(n12936), .Q(n12934) );
  xor2s1 U13453 ( .DIN1(n1452), .DIN2(n5066), .Q(n12933) );
  nnd2s1 U13454 ( .DIN1(n12937), .DIN2(n1601), .Q(n12930) );
  xor2s1 U13455 ( .DIN1(w2[29]), .DIN2(text_in_r[61]), .Q(n12937) );
  nnd3s1 U13456 ( .DIN1(n12938), .DIN2(n12939), .DIN3(n12940), .Q(N150) );
  nnd2s1 U13457 ( .DIN1(n1598), .DIN2(n12941), .Q(n12940) );
  xor2s1 U13458 ( .DIN1(w2[28]), .DIN2(text_in_r[60]), .Q(n12941) );
  nnd2s1 U13459 ( .DIN1(n12942), .DIN2(n12943), .Q(n12939) );
  nnd2s1 U13460 ( .DIN1(n12944), .DIN2(n12945), .Q(n12942) );
  nnd2s1 U13461 ( .DIN1(n12946), .DIN2(n12947), .Q(n12945) );
  nnd2s1 U13462 ( .DIN1(n12948), .DIN2(n12949), .Q(n12944) );
  nnd2s1 U13463 ( .DIN1(n12950), .DIN2(n12951), .Q(n12938) );
  nnd2s1 U13464 ( .DIN1(n12952), .DIN2(n12953), .Q(n12951) );
  nnd2s1 U13465 ( .DIN1(n12948), .DIN2(n12947), .Q(n12953) );
  nnd2s1 U13466 ( .DIN1(n12949), .DIN2(n12946), .Q(n12952) );
  hi1s1 U13467 ( .DIN(n12947), .Q(n12949) );
  xor2s1 U13468 ( .DIN1(n12954), .DIN2(n12955), .Q(n12947) );
  xor2s1 U13469 ( .DIN1(n1477), .DIN2(n5065), .Q(n12954) );
  nnd3s1 U13470 ( .DIN1(n12956), .DIN2(n12957), .DIN3(n12958), .Q(N149) );
  nnd2s1 U13471 ( .DIN1(n1598), .DIN2(n12959), .Q(n12958) );
  xor2s1 U13472 ( .DIN1(w2[27]), .DIN2(text_in_r[59]), .Q(n12959) );
  nnd2s1 U13473 ( .DIN1(n12960), .DIN2(n12961), .Q(n12957) );
  nnd2s1 U13474 ( .DIN1(n12962), .DIN2(n12963), .Q(n12960) );
  nnd2s1 U13475 ( .DIN1(n12964), .DIN2(n12965), .Q(n12963) );
  nnd2s1 U13476 ( .DIN1(n12966), .DIN2(n12967), .Q(n12962) );
  nnd2s1 U13477 ( .DIN1(n12968), .DIN2(n12969), .Q(n12956) );
  nnd2s1 U13478 ( .DIN1(n12970), .DIN2(n12971), .Q(n12969) );
  nnd2s1 U13479 ( .DIN1(n12966), .DIN2(n12965), .Q(n12971) );
  nnd2s1 U13480 ( .DIN1(n12967), .DIN2(n12964), .Q(n12970) );
  hi1s1 U13481 ( .DIN(n12965), .Q(n12967) );
  xor2s1 U13482 ( .DIN1(n12972), .DIN2(n12973), .Q(n12965) );
  xor2s1 U13483 ( .DIN1(n5064), .DIN2(w2[27]), .Q(n12972) );
  nnd2s1 U13484 ( .DIN1(n12974), .DIN2(n12975), .Q(N148) );
  nnd2s1 U13485 ( .DIN1(n12976), .DIN2(n1634), .Q(n12975) );
  xor2s1 U13486 ( .DIN1(n12977), .DIN2(n12978), .Q(n12976) );
  xor2s1 U13487 ( .DIN1(n4742), .DIN2(n12979), .Q(n12978) );
  xor2s1 U13488 ( .DIN1(n1453), .DIN2(n12980), .Q(n12977) );
  hi1s1 U13489 ( .DIN(n5063), .Q(n12980) );
  nnd2s1 U13490 ( .DIN1(n12981), .DIN2(n1600), .Q(n12974) );
  xor2s1 U13491 ( .DIN1(w2[26]), .DIN2(text_in_r[58]), .Q(n12981) );
  nnd3s1 U13492 ( .DIN1(n12982), .DIN2(n12983), .DIN3(n12984), .Q(N147) );
  nnd2s1 U13493 ( .DIN1(n1598), .DIN2(n12985), .Q(n12984) );
  xor2s1 U13494 ( .DIN1(w2[25]), .DIN2(text_in_r[57]), .Q(n12985) );
  nnd2s1 U13495 ( .DIN1(n12986), .DIN2(n12987), .Q(n12983) );
  nnd2s1 U13496 ( .DIN1(n12988), .DIN2(n12989), .Q(n12986) );
  nnd2s1 U13497 ( .DIN1(n12946), .DIN2(n12990), .Q(n12989) );
  nnd2s1 U13498 ( .DIN1(n12991), .DIN2(n12948), .Q(n12988) );
  nnd2s1 U13499 ( .DIN1(n12992), .DIN2(n12993), .Q(n12982) );
  nnd2s1 U13500 ( .DIN1(n12994), .DIN2(n12995), .Q(n12993) );
  nnd2s1 U13501 ( .DIN1(n12948), .DIN2(n12990), .Q(n12995) );
  nnd2s1 U13502 ( .DIN1(n12991), .DIN2(n12946), .Q(n12994) );
  hi1s1 U13503 ( .DIN(n12990), .Q(n12991) );
  xor2s1 U13504 ( .DIN1(n12996), .DIN2(n4753), .Q(n12990) );
  xnr2s1 U13505 ( .DIN1(w2[25]), .DIN2(n5062), .Q(n12996) );
  nnd2s1 U13506 ( .DIN1(n12997), .DIN2(n12998), .Q(N146) );
  nnd2s1 U13507 ( .DIN1(n12999), .DIN2(n1633), .Q(n12998) );
  xor2s1 U13508 ( .DIN1(n13000), .DIN2(n13001), .Q(n12999) );
  xor2s1 U13509 ( .DIN1(n12973), .DIN2(n13002), .Q(n13001) );
  xor2s1 U13510 ( .DIN1(n1454), .DIN2(n5061), .Q(n13000) );
  nnd2s1 U13511 ( .DIN1(n13003), .DIN2(n1600), .Q(n12997) );
  xor2s1 U13512 ( .DIN1(w2[24]), .DIN2(text_in_r[56]), .Q(n13003) );
  nnd3s1 U13513 ( .DIN1(n13004), .DIN2(n13005), .DIN3(n13006), .Q(N137) );
  nnd2s1 U13514 ( .DIN1(n1597), .DIN2(n13007), .Q(n13006) );
  xor2s1 U13515 ( .DIN1(w2[23]), .DIN2(text_in_r[55]), .Q(n13007) );
  nnd2s1 U13516 ( .DIN1(n13008), .DIN2(n13009), .Q(n13005) );
  nnd2s1 U13517 ( .DIN1(n13010), .DIN2(n13011), .Q(n13008) );
  nnd2s1 U13518 ( .DIN1(n13012), .DIN2(n13013), .Q(n13011) );
  nnd2s1 U13519 ( .DIN1(n13014), .DIN2(n13015), .Q(n13010) );
  nnd2s1 U13520 ( .DIN1(n5421), .DIN2(n13016), .Q(n13004) );
  nnd2s1 U13521 ( .DIN1(n13017), .DIN2(n13018), .Q(n13016) );
  nnd2s1 U13522 ( .DIN1(n13014), .DIN2(n13013), .Q(n13018) );
  nnd2s1 U13523 ( .DIN1(n13015), .DIN2(n13012), .Q(n13017) );
  hi1s1 U13524 ( .DIN(n13013), .Q(n13015) );
  xor2s1 U13525 ( .DIN1(n5067), .DIN2(n13019), .Q(n13013) );
  xnr2s1 U13526 ( .DIN1(w2[23]), .DIN2(n5043), .Q(n13019) );
  nnd2s1 U13527 ( .DIN1(n13020), .DIN2(n13021), .Q(N136) );
  nnd2s1 U13528 ( .DIN1(n13022), .DIN2(n1635), .Q(n13021) );
  xor2s1 U13529 ( .DIN1(n13023), .DIN2(n13024), .Q(n13022) );
  xor2s1 U13530 ( .DIN1(n13025), .DIN2(n12927), .Q(n13024) );
  xnr2s1 U13531 ( .DIN1(n5066), .DIN2(n13026), .Q(n13023) );
  xor2s1 U13532 ( .DIN1(n1482), .DIN2(n13027), .Q(n13026) );
  nnd2s1 U13533 ( .DIN1(n13028), .DIN2(n1600), .Q(n13020) );
  xor2s1 U13534 ( .DIN1(w2[22]), .DIN2(text_in_r[54]), .Q(n13028) );
  nnd3s1 U13535 ( .DIN1(n13029), .DIN2(n13030), .DIN3(n13031), .Q(N135) );
  nnd2s1 U13536 ( .DIN1(n1597), .DIN2(n13032), .Q(n13031) );
  xor2s1 U13537 ( .DIN1(w2[21]), .DIN2(text_in_r[53]), .Q(n13032) );
  nnd2s1 U13538 ( .DIN1(n13033), .DIN2(n13034), .Q(n13030) );
  hi1s1 U13539 ( .DIN(n12935), .Q(n13034) );
  nnd2s1 U13540 ( .DIN1(n13035), .DIN2(n13036), .Q(n13033) );
  nnd2s1 U13541 ( .DIN1(n13037), .DIN2(n13038), .Q(n13036) );
  nnd2s1 U13542 ( .DIN1(n13039), .DIN2(n13040), .Q(n13035) );
  nnd2s1 U13543 ( .DIN1(n12935), .DIN2(n13041), .Q(n13029) );
  nnd2s1 U13544 ( .DIN1(n13042), .DIN2(n13043), .Q(n13041) );
  nnd2s1 U13545 ( .DIN1(n13039), .DIN2(n13038), .Q(n13043) );
  nnd2s1 U13546 ( .DIN1(n13040), .DIN2(n13037), .Q(n13042) );
  hi1s1 U13547 ( .DIN(n13038), .Q(n13040) );
  xor2s1 U13548 ( .DIN1(n13044), .DIN2(n13045), .Q(n13038) );
  xor2s1 U13549 ( .DIN1(w2[21]), .DIN2(n5041), .Q(n13045) );
  nnd2s1 U13550 ( .DIN1(n13046), .DIN2(n13047), .Q(N134) );
  nnd2s1 U13551 ( .DIN1(n13048), .DIN2(n1634), .Q(n13047) );
  xor2s1 U13552 ( .DIN1(n13049), .DIN2(n13050), .Q(n13048) );
  xor2s1 U13553 ( .DIN1(n13051), .DIN2(n13052), .Q(n13050) );
  xor2s1 U13554 ( .DIN1(n5418), .DIN2(n13053), .Q(n13052) );
  xor2s1 U13555 ( .DIN1(n5064), .DIN2(n13054), .Q(n13049) );
  xor2s1 U13556 ( .DIN1(n1455), .DIN2(n5040), .Q(n13054) );
  nnd2s1 U13557 ( .DIN1(n13055), .DIN2(n1600), .Q(n13046) );
  xor2s1 U13558 ( .DIN1(w2[20]), .DIN2(text_in_r[52]), .Q(n13055) );
  nnd2s1 U13559 ( .DIN1(n13056), .DIN2(n13057), .Q(N133) );
  nnd2s1 U13560 ( .DIN1(n13058), .DIN2(n1635), .Q(n13057) );
  xor2s1 U13561 ( .DIN1(n13059), .DIN2(n13060), .Q(n13058) );
  xor2s1 U13562 ( .DIN1(n13061), .DIN2(n13062), .Q(n13060) );
  xor2s1 U13563 ( .DIN1(n5417), .DIN2(n12968), .Q(n13062) );
  hi1s1 U13564 ( .DIN(n12961), .Q(n12968) );
  xor2s1 U13565 ( .DIN1(n5063), .DIN2(n13063), .Q(n13059) );
  xor2s1 U13566 ( .DIN1(n1483), .DIN2(n5039), .Q(n13063) );
  nnd2s1 U13567 ( .DIN1(n13064), .DIN2(n1600), .Q(n13056) );
  xor2s1 U13568 ( .DIN1(w2[19]), .DIN2(text_in_r[51]), .Q(n13064) );
  nnd3s1 U13569 ( .DIN1(n13065), .DIN2(n13066), .DIN3(n13067), .Q(N132) );
  nnd2s1 U13570 ( .DIN1(n1598), .DIN2(n13068), .Q(n13067) );
  xor2s1 U13571 ( .DIN1(w2[18]), .DIN2(text_in_r[50]), .Q(n13068) );
  nnd2s1 U13572 ( .DIN1(n13069), .DIN2(n13070), .Q(n13066) );
  nnd2s1 U13573 ( .DIN1(n13071), .DIN2(n13072), .Q(n13069) );
  nnd2s1 U13574 ( .DIN1(n13073), .DIN2(n13074), .Q(n13072) );
  nnd2s1 U13575 ( .DIN1(n13075), .DIN2(n13076), .Q(n13071) );
  nnd2s1 U13576 ( .DIN1(n5416), .DIN2(n13077), .Q(n13065) );
  nnd2s1 U13577 ( .DIN1(n13078), .DIN2(n13079), .Q(n13077) );
  nnd2s1 U13578 ( .DIN1(n13075), .DIN2(n13074), .Q(n13079) );
  nnd2s1 U13579 ( .DIN1(n13076), .DIN2(n13073), .Q(n13078) );
  hi1s1 U13580 ( .DIN(n13074), .Q(n13076) );
  xnr2s1 U13581 ( .DIN1(n5062), .DIN2(n13080), .Q(n13074) );
  xor2s1 U13582 ( .DIN1(w2[18]), .DIN2(n4744), .Q(n13080) );
  hi1s1 U13583 ( .DIN(n13070), .Q(n5416) );
  nnd2s1 U13584 ( .DIN1(n13081), .DIN2(n13082), .Q(N131) );
  nnd2s1 U13585 ( .DIN1(n13083), .DIN2(n1634), .Q(n13082) );
  xor2s1 U13586 ( .DIN1(n13084), .DIN2(n13085), .Q(n13083) );
  xor2s1 U13587 ( .DIN1(n13051), .DIN2(n13086), .Q(n13085) );
  xor2s1 U13588 ( .DIN1(n13087), .DIN2(n12987), .Q(n13086) );
  xor2s1 U13589 ( .DIN1(n13088), .DIN2(n4754), .Q(n13084) );
  xor2s1 U13590 ( .DIN1(n1456), .DIN2(n13089), .Q(n13088) );
  nnd2s1 U13591 ( .DIN1(n13090), .DIN2(n1601), .Q(n13081) );
  xor2s1 U13592 ( .DIN1(w2[17]), .DIN2(text_in_r[49]), .Q(n13090) );
  nnd2s1 U13593 ( .DIN1(n13091), .DIN2(n13092), .Q(N130) );
  nnd2s1 U13594 ( .DIN1(n13093), .DIN2(n1636), .Q(n13092) );
  xor2s1 U13595 ( .DIN1(n13094), .DIN2(n13095), .Q(n13093) );
  xor2s1 U13596 ( .DIN1(n13002), .DIN2(n13051), .Q(n13095) );
  hi1s1 U13597 ( .DIN(n13061), .Q(n13051) );
  xor2s1 U13598 ( .DIN1(n5068), .DIN2(n5044), .Q(n13061) );
  xor2s1 U13599 ( .DIN1(n1457), .DIN2(n4741), .Q(n13094) );
  nnd2s1 U13600 ( .DIN1(n13096), .DIN2(n1600), .Q(n13091) );
  xor2s1 U13601 ( .DIN1(w2[16]), .DIN2(text_in_r[48]), .Q(n13096) );
  nnd2s1 U13602 ( .DIN1(n13097), .DIN2(n13098), .Q(N121) );
  nnd2s1 U13603 ( .DIN1(n13099), .DIN2(n1635), .Q(n13098) );
  xor2s1 U13604 ( .DIN1(n13100), .DIN2(n13101), .Q(n13099) );
  xor2s1 U13605 ( .DIN1(n12927), .DIN2(n12973), .Q(n13101) );
  xnr2s1 U13606 ( .DIN1(n5043), .DIN2(n5020), .Q(n12927) );
  xor2s1 U13607 ( .DIN1(n1458), .DIN2(n5021), .Q(n13100) );
  nnd2s1 U13608 ( .DIN1(n13102), .DIN2(n1600), .Q(n13097) );
  xor2s1 U13609 ( .DIN1(w2[15]), .DIN2(text_in_r[47]), .Q(n13102) );
  nnd2s1 U13610 ( .DIN1(n13103), .DIN2(n13104), .Q(N120) );
  nnd2s1 U13611 ( .DIN1(n13105), .DIN2(n1637), .Q(n13104) );
  xor2s1 U13612 ( .DIN1(n13106), .DIN2(n13107), .Q(n13105) );
  xor2s1 U13613 ( .DIN1(n12919), .DIN2(n12935), .Q(n13107) );
  xnr2s1 U13614 ( .DIN1(n13108), .DIN2(n5042), .Q(n12935) );
  hi1s1 U13615 ( .DIN(n13027), .Q(n5042) );
  xnr2s1 U13616 ( .DIN1(n5020), .DIN2(w2[14]), .Q(n13106) );
  nnd2s1 U13617 ( .DIN1(n13109), .DIN2(n1601), .Q(n13103) );
  xor2s1 U13618 ( .DIN1(w2[14]), .DIN2(text_in_r[46]), .Q(n13109) );
  nnd2s1 U13619 ( .DIN1(n13110), .DIN2(n13111), .Q(N119) );
  nnd2s1 U13620 ( .DIN1(n13112), .DIN2(n1637), .Q(n13111) );
  xor2s1 U13621 ( .DIN1(n13113), .DIN2(n13114), .Q(n13112) );
  xor2s1 U13622 ( .DIN1(n12928), .DIN2(n12955), .Q(n13114) );
  hi1s1 U13623 ( .DIN(n13053), .Q(n12955) );
  xor2s1 U13624 ( .DIN1(n5018), .DIN2(n5041), .Q(n13053) );
  hi1s1 U13625 ( .DIN(n13115), .Q(n5041) );
  xor2s1 U13626 ( .DIN1(n1459), .DIN2(n5019), .Q(n13113) );
  nnd2s1 U13627 ( .DIN1(n13116), .DIN2(n1599), .Q(n13110) );
  xor2s1 U13628 ( .DIN1(w2[13]), .DIN2(text_in_r[45]), .Q(n13116) );
  nnd2s1 U13629 ( .DIN1(n13117), .DIN2(n13118), .Q(N118) );
  nnd2s1 U13630 ( .DIN1(n13119), .DIN2(n1636), .Q(n13118) );
  xor2s1 U13631 ( .DIN1(n13120), .DIN2(n13121), .Q(n13119) );
  xor2s1 U13632 ( .DIN1(n12918), .DIN2(n13122), .Q(n13121) );
  xor2s1 U13633 ( .DIN1(n1460), .DIN2(n5018), .Q(n13122) );
  xor2s1 U13634 ( .DIN1(n12936), .DIN2(n12961), .Q(n13120) );
  xor2s1 U13635 ( .DIN1(n5040), .DIN2(n13123), .Q(n12961) );
  hi1s1 U13636 ( .DIN(n5017), .Q(n13123) );
  nnd2s1 U13637 ( .DIN1(n13124), .DIN2(n1599), .Q(n13117) );
  xor2s1 U13638 ( .DIN1(w2[12]), .DIN2(text_in_r[44]), .Q(n13124) );
  nnd3s1 U13639 ( .DIN1(n13125), .DIN2(n13126), .DIN3(n13127), .Q(N117) );
  nnd2s1 U13640 ( .DIN1(n1597), .DIN2(n13128), .Q(n13127) );
  xor2s1 U13641 ( .DIN1(w2[11]), .DIN2(text_in_r[43]), .Q(n13128) );
  nnd2s1 U13642 ( .DIN1(n13129), .DIN2(n12943), .Q(n13126) );
  nnd2s1 U13643 ( .DIN1(n13130), .DIN2(n13131), .Q(n13129) );
  nnd2s1 U13644 ( .DIN1(n13073), .DIN2(n13132), .Q(n13131) );
  nnd2s1 U13645 ( .DIN1(n13133), .DIN2(n13075), .Q(n13130) );
  nnd2s1 U13646 ( .DIN1(n13134), .DIN2(n12950), .Q(n13125) );
  nnd2s1 U13647 ( .DIN1(n13135), .DIN2(n13136), .Q(n13134) );
  nnd2s1 U13648 ( .DIN1(n13075), .DIN2(n13132), .Q(n13136) );
  and2s1 U13649 ( .DIN1(n12979), .DIN2(n1641), .Q(n13075) );
  nnd2s1 U13650 ( .DIN1(n13133), .DIN2(n13073), .Q(n13135) );
  nor2s1 U13651 ( .DIN1(n12979), .DIN2(n1595), .Q(n13073) );
  xor2s1 U13652 ( .DIN1(n5016), .DIN2(n5039), .Q(n12979) );
  hi1s1 U13653 ( .DIN(n13132), .Q(n13133) );
  xor2s1 U13654 ( .DIN1(n13137), .DIN2(n12918), .Q(n13132) );
  xor2s1 U13655 ( .DIN1(n5017), .DIN2(w2[11]), .Q(n13137) );
  nnd2s1 U13656 ( .DIN1(n13138), .DIN2(n13139), .Q(N116) );
  nnd2s1 U13657 ( .DIN1(n13140), .DIN2(n1636), .Q(n13139) );
  xor2s1 U13658 ( .DIN1(n13141), .DIN2(n13142), .Q(n13140) );
  xor2s1 U13659 ( .DIN1(n13143), .DIN2(n12992), .Q(n13142) );
  hi1s1 U13660 ( .DIN(n12987), .Q(n12992) );
  xor2s1 U13661 ( .DIN1(n5015), .DIN2(n4744), .Q(n12987) );
  hi1s1 U13662 ( .DIN(n5038), .Q(n4744) );
  or3s1 U13663 ( .DIN1(n13144), .DIN2(n13145), .DIN3(n13146), .Q(n5038) );
  nnd4s1 U13664 ( .DIN1(n13147), .DIN2(n13148), .DIN3(n13149), .DIN4(n13150), 
        .Q(n13146) );
  and4s1 U13665 ( .DIN1(n13151), .DIN2(n13152), .DIN3(n13153), .DIN4(n13154), 
        .Q(n13150) );
  nnd2s1 U13666 ( .DIN1(n13155), .DIN2(n13156), .Q(n13154) );
  nnd2s1 U13667 ( .DIN1(n13157), .DIN2(n13158), .Q(n13156) );
  nnd2s1 U13668 ( .DIN1(n13159), .DIN2(n13160), .Q(n13153) );
  nnd2s1 U13669 ( .DIN1(n13161), .DIN2(n13162), .Q(n13160) );
  nnd2s1 U13670 ( .DIN1(n13163), .DIN2(n13164), .Q(n13152) );
  nnd3s1 U13671 ( .DIN1(n13165), .DIN2(n13166), .DIN3(n13167), .Q(n13164) );
  nnd2s1 U13672 ( .DIN1(n13168), .DIN2(n13169), .Q(n13151) );
  nnd2s1 U13673 ( .DIN1(n13170), .DIN2(n13171), .Q(n13149) );
  nnd2s1 U13674 ( .DIN1(n13172), .DIN2(n13173), .Q(n13148) );
  nnd3s1 U13675 ( .DIN1(n13174), .DIN2(n13175), .DIN3(n13176), .Q(n13145) );
  nnd4s1 U13676 ( .DIN1(n13177), .DIN2(n13178), .DIN3(n13179), .DIN4(n13180), 
        .Q(n13144) );
  nnd2s1 U13677 ( .DIN1(n13181), .DIN2(n13182), .Q(n13180) );
  nnd2s1 U13678 ( .DIN1(n13183), .DIN2(n13184), .Q(n13179) );
  nnd2s1 U13679 ( .DIN1(n13185), .DIN2(n13186), .Q(n13178) );
  xor2s1 U13680 ( .DIN1(w2[10]), .DIN2(n5016), .Q(n13141) );
  nnd2s1 U13681 ( .DIN1(n13187), .DIN2(n1599), .Q(n13138) );
  xor2s1 U13682 ( .DIN1(w2[10]), .DIN2(text_in_r[42]), .Q(n13187) );
  nnd3s1 U13683 ( .DIN1(n13188), .DIN2(n13189), .DIN3(n13190), .Q(N115) );
  nnd2s1 U13684 ( .DIN1(n1597), .DIN2(n13191), .Q(n13190) );
  xor2s1 U13685 ( .DIN1(w2[9]), .DIN2(text_in_r[41]), .Q(n13191) );
  nnd2s1 U13686 ( .DIN1(n13192), .DIN2(n13193), .Q(n13189) );
  nnd2s1 U13687 ( .DIN1(n13194), .DIN2(n13195), .Q(n13192) );
  nnd2s1 U13688 ( .DIN1(n13012), .DIN2(n13196), .Q(n13195) );
  nnd2s1 U13689 ( .DIN1(n13002), .DIN2(n13014), .Q(n13194) );
  nnd2s1 U13690 ( .DIN1(n13197), .DIN2(n13198), .Q(n13188) );
  nnd2s1 U13691 ( .DIN1(n13199), .DIN2(n13200), .Q(n13198) );
  nnd2s1 U13692 ( .DIN1(n13014), .DIN2(n13196), .Q(n13200) );
  nor2s1 U13693 ( .DIN1(n13201), .DIN2(n1595), .Q(n13014) );
  nnd2s1 U13694 ( .DIN1(n13002), .DIN2(n13012), .Q(n13199) );
  nor2s1 U13695 ( .DIN1(n12918), .DIN2(n1594), .Q(n13012) );
  hi1s1 U13696 ( .DIN(n13196), .Q(n13002) );
  xnr2s1 U13697 ( .DIN1(n4745), .DIN2(n4754), .Q(n13196) );
  nor3s1 U13698 ( .DIN1(n13202), .DIN2(n13203), .DIN3(n13204), .Q(n4754) );
  nnd4s1 U13699 ( .DIN1(n13205), .DIN2(n13206), .DIN3(n13207), .DIN4(n13208), 
        .Q(n13204) );
  and4s1 U13700 ( .DIN1(n13209), .DIN2(n13210), .DIN3(n13211), .DIN4(n13212), 
        .Q(n13208) );
  nnd2s1 U13701 ( .DIN1(n13168), .DIN2(n13213), .Q(n13212) );
  nnd2s1 U13702 ( .DIN1(n13161), .DIN2(n13214), .Q(n13213) );
  nnd2s1 U13703 ( .DIN1(n13186), .DIN2(n13215), .Q(n13211) );
  nnd2s1 U13704 ( .DIN1(n13216), .DIN2(n13162), .Q(n13215) );
  nnd2s1 U13705 ( .DIN1(n13172), .DIN2(n13217), .Q(n13210) );
  or2s1 U13706 ( .DIN1(n13218), .DIN2(n13219), .Q(n13209) );
  nnd2s1 U13707 ( .DIN1(n13220), .DIN2(n13221), .Q(n13207) );
  nnd2s1 U13708 ( .DIN1(n13163), .DIN2(n13222), .Q(n13206) );
  nnd2s1 U13709 ( .DIN1(n13223), .DIN2(n13224), .Q(n13205) );
  nnd3s1 U13710 ( .DIN1(n13225), .DIN2(n13226), .DIN3(n13227), .Q(n13203) );
  nnd4s1 U13711 ( .DIN1(n13177), .DIN2(n13228), .DIN3(n13229), .DIN4(n13230), 
        .Q(n13202) );
  nnd2s1 U13712 ( .DIN1(n13173), .DIN2(n13231), .Q(n13230) );
  nnd2s1 U13713 ( .DIN1(n13185), .DIN2(n13232), .Q(n13228) );
  nor3s1 U13714 ( .DIN1(n13233), .DIN2(n13234), .DIN3(n13235), .Q(n13177) );
  nnd4s1 U13715 ( .DIN1(n13236), .DIN2(n13237), .DIN3(n13238), .DIN4(n13239), 
        .Q(n13235) );
  and3s1 U13716 ( .DIN1(n13240), .DIN2(n13241), .DIN3(n13242), .Q(n13239) );
  nnd2s1 U13717 ( .DIN1(n13183), .DIN2(n13159), .Q(n13242) );
  nnd2s1 U13718 ( .DIN1(n13170), .DIN2(n13221), .Q(n13241) );
  nnd2s1 U13719 ( .DIN1(n13186), .DIN2(n13243), .Q(n13240) );
  nnd3s1 U13720 ( .DIN1(n13244), .DIN2(n13245), .DIN3(n13246), .Q(n13234) );
  nnd2s1 U13721 ( .DIN1(n13172), .DIN2(n13155), .Q(n13246) );
  nnd2s1 U13722 ( .DIN1(n13231), .DIN2(n13247), .Q(n13245) );
  nnd2s1 U13723 ( .DIN1(n13248), .DIN2(n13249), .Q(n13244) );
  nnd4s1 U13724 ( .DIN1(n13250), .DIN2(n13251), .DIN3(n13252), .DIN4(n13253), 
        .Q(n13233) );
  nnd2s1 U13725 ( .DIN1(n13185), .DIN2(n13254), .Q(n13253) );
  nnd2s1 U13726 ( .DIN1(n13255), .DIN2(n13256), .Q(n13254) );
  nnd2s1 U13727 ( .DIN1(n13220), .DIN2(n13257), .Q(n13252) );
  nnd4s1 U13728 ( .DIN1(n13256), .DIN2(n13166), .DIN3(n13158), .DIN4(n13258), 
        .Q(n13257) );
  nnd2s1 U13729 ( .DIN1(n13259), .DIN2(n13260), .Q(n13251) );
  nnd2s1 U13730 ( .DIN1(n13261), .DIN2(n13262), .Q(n13250) );
  hi1s1 U13731 ( .DIN(n13193), .Q(n13197) );
  xor2s1 U13732 ( .DIN1(n13263), .DIN2(n4742), .Q(n13193) );
  xor2s1 U13733 ( .DIN1(n13089), .DIN2(n5062), .Q(n4742) );
  nor3s1 U13734 ( .DIN1(n13264), .DIN2(n13265), .DIN3(n13266), .Q(n5062) );
  nnd4s1 U13735 ( .DIN1(n13267), .DIN2(n13268), .DIN3(n13269), .DIN4(n13270), 
        .Q(n13266) );
  and4s1 U13736 ( .DIN1(n13271), .DIN2(n13272), .DIN3(n13273), .DIN4(n13274), 
        .Q(n13270) );
  nnd2s1 U13737 ( .DIN1(n13275), .DIN2(n13276), .Q(n13274) );
  nnd2s1 U13738 ( .DIN1(n13277), .DIN2(n13278), .Q(n13276) );
  nnd2s1 U13739 ( .DIN1(n13279), .DIN2(n13280), .Q(n13273) );
  nnd2s1 U13740 ( .DIN1(n13281), .DIN2(n13282), .Q(n13280) );
  nnd2s1 U13741 ( .DIN1(n13283), .DIN2(n13284), .Q(n13272) );
  nnd3s1 U13742 ( .DIN1(n13285), .DIN2(n13286), .DIN3(n13287), .Q(n13284) );
  nnd2s1 U13743 ( .DIN1(n13288), .DIN2(n13289), .Q(n13271) );
  nnd2s1 U13744 ( .DIN1(n13290), .DIN2(n13291), .Q(n13269) );
  nnd2s1 U13745 ( .DIN1(n13292), .DIN2(n13293), .Q(n13268) );
  nnd3s1 U13746 ( .DIN1(n13294), .DIN2(n13295), .DIN3(n13296), .Q(n13265) );
  nnd4s1 U13747 ( .DIN1(n13297), .DIN2(n13298), .DIN3(n13299), .DIN4(n13300), 
        .Q(n13264) );
  nnd2s1 U13748 ( .DIN1(n13301), .DIN2(n13302), .Q(n13300) );
  nnd2s1 U13749 ( .DIN1(n13303), .DIN2(n13304), .Q(n13299) );
  nnd2s1 U13750 ( .DIN1(n13305), .DIN2(n13306), .Q(n13298) );
  xor2s1 U13751 ( .DIN1(n5015), .DIN2(w2[9]), .Q(n13263) );
  nnd2s1 U13752 ( .DIN1(n13307), .DIN2(n13308), .Q(N114) );
  nnd2s1 U13753 ( .DIN1(n13309), .DIN2(n1638), .Q(n13308) );
  xor2s1 U13754 ( .DIN1(n13310), .DIN2(n13311), .Q(n13309) );
  xor2s1 U13755 ( .DIN1(n4753), .DIN2(n12918), .Q(n13311) );
  hi1s1 U13756 ( .DIN(n13201), .Q(n12918) );
  xnr2s1 U13757 ( .DIN1(n5021), .DIN2(n5044), .Q(n13201) );
  xor2s1 U13758 ( .DIN1(n4741), .DIN2(n5061), .Q(n4753) );
  hi1s1 U13759 ( .DIN(n13087), .Q(n5061) );
  or3s1 U13760 ( .DIN1(n13312), .DIN2(n13313), .DIN3(n13314), .Q(n13087) );
  nnd4s1 U13761 ( .DIN1(n13315), .DIN2(n13316), .DIN3(n13317), .DIN4(n13318), 
        .Q(n13314) );
  and4s1 U13762 ( .DIN1(n13319), .DIN2(n13320), .DIN3(n13321), .DIN4(n13322), 
        .Q(n13318) );
  nnd2s1 U13763 ( .DIN1(n13288), .DIN2(n13323), .Q(n13322) );
  nnd2s1 U13764 ( .DIN1(n13281), .DIN2(n13324), .Q(n13323) );
  nnd2s1 U13765 ( .DIN1(n13306), .DIN2(n13325), .Q(n13321) );
  nnd2s1 U13766 ( .DIN1(n13326), .DIN2(n13282), .Q(n13325) );
  nnd2s1 U13767 ( .DIN1(n13292), .DIN2(n13327), .Q(n13320) );
  or2s1 U13768 ( .DIN1(n13328), .DIN2(n13329), .Q(n13319) );
  nnd2s1 U13769 ( .DIN1(n13330), .DIN2(n13331), .Q(n13317) );
  nnd2s1 U13770 ( .DIN1(n13283), .DIN2(n13332), .Q(n13316) );
  nnd2s1 U13771 ( .DIN1(n13333), .DIN2(n13334), .Q(n13315) );
  nnd3s1 U13772 ( .DIN1(n13335), .DIN2(n13336), .DIN3(n13337), .Q(n13313) );
  nnd4s1 U13773 ( .DIN1(n13297), .DIN2(n13338), .DIN3(n13339), .DIN4(n13340), 
        .Q(n13312) );
  nnd2s1 U13774 ( .DIN1(n13293), .DIN2(n13341), .Q(n13340) );
  nnd2s1 U13775 ( .DIN1(n13305), .DIN2(n13342), .Q(n13338) );
  nor3s1 U13776 ( .DIN1(n13343), .DIN2(n13344), .DIN3(n13345), .Q(n13297) );
  nnd4s1 U13777 ( .DIN1(n13346), .DIN2(n13347), .DIN3(n13348), .DIN4(n13349), 
        .Q(n13345) );
  and3s1 U13778 ( .DIN1(n13350), .DIN2(n13351), .DIN3(n13352), .Q(n13349) );
  nnd2s1 U13779 ( .DIN1(n13303), .DIN2(n13279), .Q(n13352) );
  nnd2s1 U13780 ( .DIN1(n13290), .DIN2(n13331), .Q(n13351) );
  nnd2s1 U13781 ( .DIN1(n13306), .DIN2(n13353), .Q(n13350) );
  nnd3s1 U13782 ( .DIN1(n13354), .DIN2(n13355), .DIN3(n13356), .Q(n13344) );
  nnd2s1 U13783 ( .DIN1(n13292), .DIN2(n13275), .Q(n13356) );
  nnd2s1 U13784 ( .DIN1(n13341), .DIN2(n13357), .Q(n13355) );
  nnd2s1 U13785 ( .DIN1(n13358), .DIN2(n13359), .Q(n13354) );
  nnd4s1 U13786 ( .DIN1(n13360), .DIN2(n13361), .DIN3(n13362), .DIN4(n13363), 
        .Q(n13343) );
  nnd2s1 U13787 ( .DIN1(n13305), .DIN2(n13364), .Q(n13363) );
  nnd2s1 U13788 ( .DIN1(n13365), .DIN2(n13366), .Q(n13364) );
  nnd2s1 U13789 ( .DIN1(n13330), .DIN2(n13367), .Q(n13362) );
  nnd4s1 U13790 ( .DIN1(n13366), .DIN2(n13286), .DIN3(n13278), .DIN4(n13368), 
        .Q(n13367) );
  nnd2s1 U13791 ( .DIN1(n13369), .DIN2(n13370), .Q(n13361) );
  nnd2s1 U13792 ( .DIN1(n13371), .DIN2(n13372), .Q(n13360) );
  nor4s1 U13793 ( .DIN1(n13373), .DIN2(n13374), .DIN3(n13375), .DIN4(n13376), 
        .Q(n4741) );
  nnd4s1 U13794 ( .DIN1(n13377), .DIN2(n13378), .DIN3(n13379), .DIN4(n13380), 
        .Q(n13376) );
  nnd2s1 U13795 ( .DIN1(n13381), .DIN2(n13382), .Q(n13380) );
  nnd2s1 U13796 ( .DIN1(n13383), .DIN2(n13384), .Q(n13379) );
  nnd2s1 U13797 ( .DIN1(n13385), .DIN2(n13386), .Q(n13378) );
  nnd2s1 U13798 ( .DIN1(n13387), .DIN2(n13388), .Q(n13377) );
  nnd4s1 U13799 ( .DIN1(n13389), .DIN2(n13390), .DIN3(n13391), .DIN4(n13392), 
        .Q(n13375) );
  nnd2s1 U13800 ( .DIN1(n13393), .DIN2(n13394), .Q(n13392) );
  nnd2s1 U13801 ( .DIN1(n13395), .DIN2(n13396), .Q(n13394) );
  nnd2s1 U13802 ( .DIN1(n13397), .DIN2(n13398), .Q(n13391) );
  nnd2s1 U13803 ( .DIN1(n13399), .DIN2(n13400), .Q(n13398) );
  or2s1 U13804 ( .DIN1(n13401), .DIN2(n13402), .Q(n13390) );
  nnd2s1 U13805 ( .DIN1(n13403), .DIN2(n13404), .Q(n13389) );
  nnd3s1 U13806 ( .DIN1(n13405), .DIN2(n13406), .DIN3(n13407), .Q(n13374) );
  nnd4s1 U13807 ( .DIN1(n13408), .DIN2(n13409), .DIN3(n13410), .DIN4(n13411), 
        .Q(n13373) );
  nnd2s1 U13808 ( .DIN1(n13412), .DIN2(n13413), .Q(n13410) );
  nnd2s1 U13809 ( .DIN1(n13414), .DIN2(n13415), .Q(n13409) );
  xor2s1 U13810 ( .DIN1(n1461), .DIN2(n4745), .Q(n13310) );
  nor4s1 U13811 ( .DIN1(n13416), .DIN2(n13417), .DIN3(n13418), .DIN4(n13419), 
        .Q(n4745) );
  nnd4s1 U13812 ( .DIN1(n13420), .DIN2(n13421), .DIN3(n13422), .DIN4(n13423), 
        .Q(n13419) );
  nnd2s1 U13813 ( .DIN1(n13424), .DIN2(n13425), .Q(n13423) );
  nnd2s1 U13814 ( .DIN1(n13426), .DIN2(n13427), .Q(n13422) );
  nnd2s1 U13815 ( .DIN1(n13428), .DIN2(n13429), .Q(n13421) );
  nnd2s1 U13816 ( .DIN1(n13430), .DIN2(n13431), .Q(n13420) );
  nnd4s1 U13817 ( .DIN1(n13432), .DIN2(n13433), .DIN3(n13434), .DIN4(n13435), 
        .Q(n13418) );
  nnd2s1 U13818 ( .DIN1(n13436), .DIN2(n13437), .Q(n13435) );
  nnd2s1 U13819 ( .DIN1(n13438), .DIN2(n13439), .Q(n13437) );
  nnd2s1 U13820 ( .DIN1(n13440), .DIN2(n13441), .Q(n13434) );
  nnd2s1 U13821 ( .DIN1(n13442), .DIN2(n13443), .Q(n13441) );
  or2s1 U13822 ( .DIN1(n13444), .DIN2(n13445), .Q(n13433) );
  nnd2s1 U13823 ( .DIN1(n13446), .DIN2(n13447), .Q(n13432) );
  nnd3s1 U13824 ( .DIN1(n13448), .DIN2(n13449), .DIN3(n13450), .Q(n13417) );
  nnd4s1 U13825 ( .DIN1(n13451), .DIN2(n13452), .DIN3(n13453), .DIN4(n13454), 
        .Q(n13416) );
  nnd2s1 U13826 ( .DIN1(n13455), .DIN2(n13456), .Q(n13453) );
  nnd2s1 U13827 ( .DIN1(n13457), .DIN2(n13458), .Q(n13452) );
  nnd2s1 U13828 ( .DIN1(n13459), .DIN2(n1600), .Q(n13307) );
  xor2s1 U13829 ( .DIN1(w2[8]), .DIN2(text_in_r[40]), .Q(n13459) );
  nnd3s1 U13830 ( .DIN1(n13460), .DIN2(n13461), .DIN3(n13462), .Q(N105) );
  nnd2s1 U13831 ( .DIN1(n1596), .DIN2(n13463), .Q(n13462) );
  xor2s1 U13832 ( .DIN1(w2[7]), .DIN2(text_in_r[39]), .Q(n13463) );
  nnd2s1 U13833 ( .DIN1(n13464), .DIN2(n5420), .Q(n13461) );
  nnd2s1 U13834 ( .DIN1(n13465), .DIN2(n13466), .Q(n13464) );
  nnd2s1 U13835 ( .DIN1(n12946), .DIN2(n13467), .Q(n13466) );
  nnd2s1 U13836 ( .DIN1(n13468), .DIN2(n12948), .Q(n13465) );
  nnd2s1 U13837 ( .DIN1(n13025), .DIN2(n13469), .Q(n13460) );
  nnd2s1 U13838 ( .DIN1(n13470), .DIN2(n13471), .Q(n13469) );
  nnd2s1 U13839 ( .DIN1(n12948), .DIN2(n13467), .Q(n13471) );
  and2s1 U13840 ( .DIN1(n12973), .DIN2(n1543), .Q(n12948) );
  nnd2s1 U13841 ( .DIN1(n13468), .DIN2(n12946), .Q(n13470) );
  nor2s1 U13842 ( .DIN1(n12973), .DIN2(n1594), .Q(n12946) );
  xor2s1 U13843 ( .DIN1(n13009), .DIN2(n5068), .Q(n12973) );
  or3s1 U13844 ( .DIN1(n13472), .DIN2(n13473), .DIN3(n13474), .Q(n5068) );
  nnd4s1 U13845 ( .DIN1(n13337), .DIN2(n13294), .DIN3(n13475), .DIN4(n13476), 
        .Q(n13474) );
  and4s1 U13846 ( .DIN1(n13346), .DIN2(n13477), .DIN3(n13478), .DIN4(n13479), 
        .Q(n13476) );
  nnd2s1 U13847 ( .DIN1(n13301), .DIN2(n13480), .Q(n13479) );
  nnd2s1 U13848 ( .DIN1(n13288), .DIN2(n13353), .Q(n13478) );
  and4s1 U13849 ( .DIN1(n13481), .DIN2(n13482), .DIN3(n13483), .DIN4(n13484), 
        .Q(n13346) );
  and4s1 U13850 ( .DIN1(n13485), .DIN2(n13486), .DIN3(n13487), .DIN4(n13488), 
        .Q(n13484) );
  nnd2s1 U13851 ( .DIN1(n13333), .DIN2(n13288), .Q(n13488) );
  nnd2s1 U13852 ( .DIN1(n13489), .DIN2(n13490), .Q(n13487) );
  nnd2s1 U13853 ( .DIN1(n13303), .DIN2(n13291), .Q(n13486) );
  nnd2s1 U13854 ( .DIN1(n13371), .DIN2(n13480), .Q(n13485) );
  and3s1 U13855 ( .DIN1(n13491), .DIN2(n13492), .DIN3(n13493), .Q(n13483) );
  nnd2s1 U13856 ( .DIN1(n13290), .DIN2(n13494), .Q(n13493) );
  nnd3s1 U13857 ( .DIN1(n13495), .DIN2(n13496), .DIN3(n13286), .Q(n13494) );
  nnd2s1 U13858 ( .DIN1(n13331), .DIN2(n13497), .Q(n13492) );
  nnd2s1 U13859 ( .DIN1(n13498), .DIN2(n13499), .Q(n13497) );
  nnd2s1 U13860 ( .DIN1(n13500), .DIN2(n13501), .Q(n13491) );
  nnd2s1 U13861 ( .DIN1(n13502), .DIN2(n13368), .Q(n13501) );
  nnd2s1 U13862 ( .DIN1(n13292), .DIN2(n13503), .Q(n13482) );
  nnd4s1 U13863 ( .DIN1(n13328), .DIN2(n13504), .DIN3(n13281), .DIN4(n13505), 
        .Q(n13503) );
  nnd2s1 U13864 ( .DIN1(n13275), .DIN2(n13359), .Q(n13481) );
  nor2s1 U13865 ( .DIN1(n13506), .DIN2(n13507), .Q(n13294) );
  nnd4s1 U13866 ( .DIN1(n13508), .DIN2(n13509), .DIN3(n13510), .DIN4(n13511), 
        .Q(n13507) );
  nnd2s1 U13867 ( .DIN1(n13500), .DIN2(n13512), .Q(n13511) );
  nnd2s1 U13868 ( .DIN1(n13303), .DIN2(n13371), .Q(n13510) );
  nnd2s1 U13869 ( .DIN1(n13283), .DIN2(n13288), .Q(n13509) );
  nnd2s1 U13870 ( .DIN1(n13369), .DIN2(n13330), .Q(n13508) );
  nnd4s1 U13871 ( .DIN1(n13513), .DIN2(n13514), .DIN3(n13515), .DIN4(n13516), 
        .Q(n13506) );
  nnd2s1 U13872 ( .DIN1(n13490), .DIN2(n13517), .Q(n13516) );
  or2s1 U13873 ( .DIN1(n13332), .DIN2(n13304), .Q(n13517) );
  nnd2s1 U13874 ( .DIN1(n13342), .DIN2(n13518), .Q(n13515) );
  nnd2s1 U13875 ( .DIN1(n13519), .DIN2(n13520), .Q(n13518) );
  nnd2s1 U13876 ( .DIN1(n13353), .DIN2(n13521), .Q(n13514) );
  nnd2s1 U13877 ( .DIN1(n13293), .DIN2(n13522), .Q(n13513) );
  nnd3s1 U13878 ( .DIN1(n13366), .DIN2(n13277), .DIN3(n13523), .Q(n13522) );
  nor4s1 U13879 ( .DIN1(n13524), .DIN2(n13525), .DIN3(n13526), .DIN4(n13527), 
        .Q(n13337) );
  nnd4s1 U13880 ( .DIN1(n13528), .DIN2(n13529), .DIN3(n13530), .DIN4(n13531), 
        .Q(n13527) );
  nor2s1 U13881 ( .DIN1(n13532), .DIN2(n13533), .Q(n13531) );
  nor2s1 U13882 ( .DIN1(n13499), .DIN2(n13502), .Q(n13533) );
  nor2s1 U13883 ( .DIN1(n13519), .DIN2(n13365), .Q(n13532) );
  nnd2s1 U13884 ( .DIN1(n13489), .DIN2(n13275), .Q(n13530) );
  nnd2s1 U13885 ( .DIN1(n13303), .DIN2(n13331), .Q(n13529) );
  nnd2s1 U13886 ( .DIN1(n13371), .DIN2(n13293), .Q(n13528) );
  nnd3s1 U13887 ( .DIN1(n13534), .DIN2(n13535), .DIN3(n13536), .Q(n13526) );
  nnd2s1 U13888 ( .DIN1(n13342), .DIN2(n13537), .Q(n13536) );
  nnd2s1 U13889 ( .DIN1(n13333), .DIN2(n13538), .Q(n13535) );
  nnd3s1 U13890 ( .DIN1(n13286), .DIN2(n13278), .DIN3(n13366), .Q(n13538) );
  nnd2s1 U13891 ( .DIN1(n13539), .DIN2(n13540), .Q(n13534) );
  nnd3s1 U13892 ( .DIN1(n13495), .DIN2(n13541), .DIN3(n13285), .Q(n13540) );
  nor2s1 U13893 ( .DIN1(n13324), .DIN2(n13496), .Q(n13525) );
  nor2s1 U13894 ( .DIN1(n13542), .DIN2(n13498), .Q(n13524) );
  nnd4s1 U13895 ( .DIN1(n13543), .DIN2(n13544), .DIN3(n13545), .DIN4(n13546), 
        .Q(n13473) );
  nnd2s1 U13896 ( .DIN1(n13275), .DIN2(n13547), .Q(n13546) );
  nnd2s1 U13897 ( .DIN1(n13293), .DIN2(n13359), .Q(n13545) );
  nnd2s1 U13898 ( .DIN1(n13333), .DIN2(n13371), .Q(n13544) );
  nnd2s1 U13899 ( .DIN1(n13548), .DIN2(n13283), .Q(n13543) );
  nnd4s1 U13900 ( .DIN1(n13549), .DIN2(n13550), .DIN3(n13551), .DIN4(n13552), 
        .Q(n13472) );
  nnd2s1 U13901 ( .DIN1(n13553), .DIN2(n13554), .Q(n13552) );
  nnd2s1 U13902 ( .DIN1(n13282), .DIN2(n13555), .Q(n13554) );
  nnd2s1 U13903 ( .DIN1(n13304), .DIN2(n13556), .Q(n13551) );
  nnd2s1 U13904 ( .DIN1(n13557), .DIN2(n13520), .Q(n13556) );
  nnd2s1 U13905 ( .DIN1(n13303), .DIN2(n13521), .Q(n13550) );
  nnd2s1 U13906 ( .DIN1(n13366), .DIN2(n13558), .Q(n13521) );
  or2s1 U13907 ( .DIN1(n13495), .DIN2(n13559), .Q(n13549) );
  hi1s1 U13908 ( .DIN(n13467), .Q(n13468) );
  xor2s1 U13909 ( .DIN1(n13560), .DIN2(n5044), .Q(n13467) );
  nor3s1 U13910 ( .DIN1(n13561), .DIN2(n13562), .DIN3(n13563), .Q(n5044) );
  nnd4s1 U13911 ( .DIN1(n13227), .DIN2(n13174), .DIN3(n13564), .DIN4(n13565), 
        .Q(n13563) );
  and4s1 U13912 ( .DIN1(n13236), .DIN2(n13566), .DIN3(n13567), .DIN4(n13568), 
        .Q(n13565) );
  nnd2s1 U13913 ( .DIN1(n13181), .DIN2(n13569), .Q(n13568) );
  nnd2s1 U13914 ( .DIN1(n13168), .DIN2(n13243), .Q(n13567) );
  and4s1 U13915 ( .DIN1(n13570), .DIN2(n13571), .DIN3(n13572), .DIN4(n13573), 
        .Q(n13236) );
  and4s1 U13916 ( .DIN1(n13574), .DIN2(n13575), .DIN3(n13576), .DIN4(n13577), 
        .Q(n13573) );
  nnd2s1 U13917 ( .DIN1(n13223), .DIN2(n13168), .Q(n13577) );
  nnd2s1 U13918 ( .DIN1(n13578), .DIN2(n13579), .Q(n13576) );
  nnd2s1 U13919 ( .DIN1(n13183), .DIN2(n13171), .Q(n13575) );
  nnd2s1 U13920 ( .DIN1(n13261), .DIN2(n13569), .Q(n13574) );
  and3s1 U13921 ( .DIN1(n13580), .DIN2(n13581), .DIN3(n13582), .Q(n13572) );
  nnd2s1 U13922 ( .DIN1(n13170), .DIN2(n13583), .Q(n13582) );
  nnd3s1 U13923 ( .DIN1(n13584), .DIN2(n13585), .DIN3(n13166), .Q(n13583) );
  nnd2s1 U13924 ( .DIN1(n13221), .DIN2(n13586), .Q(n13581) );
  nnd2s1 U13925 ( .DIN1(n13587), .DIN2(n13588), .Q(n13586) );
  nnd2s1 U13926 ( .DIN1(n13589), .DIN2(n13590), .Q(n13580) );
  nnd2s1 U13927 ( .DIN1(n13591), .DIN2(n13258), .Q(n13590) );
  nnd2s1 U13928 ( .DIN1(n13172), .DIN2(n13592), .Q(n13571) );
  nnd4s1 U13929 ( .DIN1(n13218), .DIN2(n13593), .DIN3(n13161), .DIN4(n13594), 
        .Q(n13592) );
  nnd2s1 U13930 ( .DIN1(n13155), .DIN2(n13249), .Q(n13570) );
  nor2s1 U13931 ( .DIN1(n13595), .DIN2(n13596), .Q(n13174) );
  nnd4s1 U13932 ( .DIN1(n13597), .DIN2(n13598), .DIN3(n13599), .DIN4(n13600), 
        .Q(n13596) );
  nnd2s1 U13933 ( .DIN1(n13589), .DIN2(n13601), .Q(n13600) );
  nnd2s1 U13934 ( .DIN1(n13183), .DIN2(n13261), .Q(n13599) );
  nnd2s1 U13935 ( .DIN1(n13163), .DIN2(n13168), .Q(n13598) );
  nnd2s1 U13936 ( .DIN1(n13259), .DIN2(n13220), .Q(n13597) );
  nnd4s1 U13937 ( .DIN1(n13602), .DIN2(n13603), .DIN3(n13604), .DIN4(n13605), 
        .Q(n13595) );
  nnd2s1 U13938 ( .DIN1(n13579), .DIN2(n13606), .Q(n13605) );
  or2s1 U13939 ( .DIN1(n13222), .DIN2(n13184), .Q(n13606) );
  nnd2s1 U13940 ( .DIN1(n13232), .DIN2(n13607), .Q(n13604) );
  nnd2s1 U13941 ( .DIN1(n13608), .DIN2(n13609), .Q(n13607) );
  nnd2s1 U13942 ( .DIN1(n13243), .DIN2(n13610), .Q(n13603) );
  nnd2s1 U13943 ( .DIN1(n13173), .DIN2(n13611), .Q(n13602) );
  nnd3s1 U13944 ( .DIN1(n13256), .DIN2(n13157), .DIN3(n13612), .Q(n13611) );
  nor4s1 U13945 ( .DIN1(n13613), .DIN2(n13614), .DIN3(n13615), .DIN4(n13616), 
        .Q(n13227) );
  nnd4s1 U13946 ( .DIN1(n13617), .DIN2(n13618), .DIN3(n13619), .DIN4(n13620), 
        .Q(n13616) );
  nor2s1 U13947 ( .DIN1(n13621), .DIN2(n13622), .Q(n13620) );
  nor2s1 U13948 ( .DIN1(n13588), .DIN2(n13591), .Q(n13622) );
  nor2s1 U13949 ( .DIN1(n13608), .DIN2(n13255), .Q(n13621) );
  nnd2s1 U13950 ( .DIN1(n13578), .DIN2(n13155), .Q(n13619) );
  nnd2s1 U13951 ( .DIN1(n13183), .DIN2(n13221), .Q(n13618) );
  nnd2s1 U13952 ( .DIN1(n13261), .DIN2(n13173), .Q(n13617) );
  nnd3s1 U13953 ( .DIN1(n13623), .DIN2(n13624), .DIN3(n13625), .Q(n13615) );
  nnd2s1 U13954 ( .DIN1(n13232), .DIN2(n13626), .Q(n13625) );
  nnd2s1 U13955 ( .DIN1(n13223), .DIN2(n13627), .Q(n13624) );
  nnd3s1 U13956 ( .DIN1(n13166), .DIN2(n13158), .DIN3(n13256), .Q(n13627) );
  nnd2s1 U13957 ( .DIN1(n13628), .DIN2(n13629), .Q(n13623) );
  nnd3s1 U13958 ( .DIN1(n13584), .DIN2(n13630), .DIN3(n13165), .Q(n13629) );
  nor2s1 U13959 ( .DIN1(n13214), .DIN2(n13585), .Q(n13614) );
  nor2s1 U13960 ( .DIN1(n13631), .DIN2(n13587), .Q(n13613) );
  nnd4s1 U13961 ( .DIN1(n13632), .DIN2(n13633), .DIN3(n13634), .DIN4(n13635), 
        .Q(n13562) );
  nnd2s1 U13962 ( .DIN1(n13155), .DIN2(n13636), .Q(n13635) );
  nnd2s1 U13963 ( .DIN1(n13173), .DIN2(n13249), .Q(n13634) );
  nnd2s1 U13964 ( .DIN1(n13223), .DIN2(n13261), .Q(n13633) );
  nnd2s1 U13965 ( .DIN1(n13637), .DIN2(n13163), .Q(n13632) );
  nnd4s1 U13966 ( .DIN1(n13638), .DIN2(n13639), .DIN3(n13640), .DIN4(n13641), 
        .Q(n13561) );
  nnd2s1 U13967 ( .DIN1(n13642), .DIN2(n13643), .Q(n13641) );
  nnd2s1 U13968 ( .DIN1(n13162), .DIN2(n13644), .Q(n13643) );
  nnd2s1 U13969 ( .DIN1(n13184), .DIN2(n13645), .Q(n13640) );
  nnd2s1 U13970 ( .DIN1(n13646), .DIN2(n13609), .Q(n13645) );
  nnd2s1 U13971 ( .DIN1(n13183), .DIN2(n13610), .Q(n13639) );
  nnd2s1 U13972 ( .DIN1(n13256), .DIN2(n13647), .Q(n13610) );
  or2s1 U13973 ( .DIN1(n13584), .DIN2(n13648), .Q(n13638) );
  xnr2s1 U13974 ( .DIN1(n5020), .DIN2(w2[7]), .Q(n13560) );
  nor3s1 U13975 ( .DIN1(n13649), .DIN2(n13650), .DIN3(n13651), .Q(n5020) );
  nnd4s1 U13976 ( .DIN1(n13652), .DIN2(n13653), .DIN3(n13654), .DIN4(n13655), 
        .Q(n13651) );
  and3s1 U13977 ( .DIN1(n13656), .DIN2(n13657), .DIN3(n13658), .Q(n13655) );
  nnd2s1 U13978 ( .DIN1(n13659), .DIN2(n13660), .Q(n13653) );
  nnd3s1 U13979 ( .DIN1(n13661), .DIN2(n13662), .DIN3(n13663), .Q(n13650) );
  or2s1 U13980 ( .DIN1(n13664), .DIN2(n13665), .Q(n13663) );
  nnd2s1 U13981 ( .DIN1(n13429), .DIN2(n13666), .Q(n13662) );
  or2s1 U13982 ( .DIN1(n13667), .DIN2(n13668), .Q(n13661) );
  nnd3s1 U13983 ( .DIN1(n13669), .DIN2(n13670), .DIN3(n13671), .Q(n13649) );
  nnd2s1 U13984 ( .DIN1(n13436), .DIN2(n13672), .Q(n13671) );
  nnd2s1 U13985 ( .DIN1(n13673), .DIN2(n13674), .Q(n13672) );
  nnd2s1 U13986 ( .DIN1(n13675), .DIN2(n13676), .Q(n13670) );
  nnd2s1 U13987 ( .DIN1(n13438), .DIN2(n13677), .Q(n13675) );
  nnd2s1 U13988 ( .DIN1(n13678), .DIN2(n13679), .Q(n13669) );
  nnd2s1 U13989 ( .DIN1(n13680), .DIN2(n13681), .Q(n13679) );
  nnd3s1 U13990 ( .DIN1(n13682), .DIN2(n13683), .DIN3(n13684), .Q(N104) );
  nnd2s1 U13991 ( .DIN1(n1596), .DIN2(n13685), .Q(n13684) );
  xor2s1 U13992 ( .DIN1(w2[6]), .DIN2(text_in_r[38]), .Q(n13685) );
  nnd2s1 U13993 ( .DIN1(n13686), .DIN2(n13687), .Q(n13683) );
  nnd2s1 U13994 ( .DIN1(n13688), .DIN2(n13689), .Q(n13686) );
  nnd2s1 U13995 ( .DIN1(n13037), .DIN2(n13690), .Q(n13689) );
  nnd2s1 U13996 ( .DIN1(n12919), .DIN2(n13039), .Q(n13688) );
  nnd2s1 U13997 ( .DIN1(n13691), .DIN2(n13692), .Q(n13682) );
  nnd2s1 U13998 ( .DIN1(n13693), .DIN2(n13694), .Q(n13692) );
  nnd2s1 U13999 ( .DIN1(n13039), .DIN2(n13690), .Q(n13694) );
  nor2s1 U14000 ( .DIN1(n13695), .DIN2(n1594), .Q(n13039) );
  nnd2s1 U14001 ( .DIN1(n12919), .DIN2(n13037), .Q(n13693) );
  nor2s1 U14002 ( .DIN1(n5419), .DIN2(n1594), .Q(n13037) );
  hi1s1 U14003 ( .DIN(n13695), .Q(n5419) );
  hi1s1 U14004 ( .DIN(n13690), .Q(n12919) );
  xor2s1 U14005 ( .DIN1(n5067), .DIN2(n13025), .Q(n13690) );
  hi1s1 U14006 ( .DIN(n5420), .Q(n13025) );
  or3s1 U14007 ( .DIN1(n13696), .DIN2(n13697), .DIN3(n13698), .Q(n5420) );
  nnd4s1 U14008 ( .DIN1(n13699), .DIN2(n13700), .DIN3(n13701), .DIN4(n13702), 
        .Q(n13698) );
  and3s1 U14009 ( .DIN1(n13703), .DIN2(n13704), .DIN3(n13705), .Q(n13702) );
  nnd2s1 U14010 ( .DIN1(n13706), .DIN2(n13707), .Q(n13700) );
  nnd3s1 U14011 ( .DIN1(n13708), .DIN2(n13709), .DIN3(n13710), .Q(n13697) );
  or2s1 U14012 ( .DIN1(n13711), .DIN2(n13712), .Q(n13710) );
  nnd2s1 U14013 ( .DIN1(n13386), .DIN2(n13713), .Q(n13709) );
  or2s1 U14014 ( .DIN1(n13714), .DIN2(n13715), .Q(n13708) );
  nnd3s1 U14015 ( .DIN1(n13716), .DIN2(n13717), .DIN3(n13718), .Q(n13696) );
  nnd2s1 U14016 ( .DIN1(n13393), .DIN2(n13719), .Q(n13718) );
  nnd2s1 U14017 ( .DIN1(n13720), .DIN2(n13721), .Q(n13719) );
  nnd2s1 U14018 ( .DIN1(n13722), .DIN2(n13723), .Q(n13717) );
  nnd2s1 U14019 ( .DIN1(n13395), .DIN2(n13724), .Q(n13722) );
  nnd2s1 U14020 ( .DIN1(n13725), .DIN2(n13726), .Q(n13716) );
  nnd2s1 U14021 ( .DIN1(n13727), .DIN2(n13728), .Q(n13726) );
  or3s1 U14022 ( .DIN1(n13729), .DIN2(n13730), .DIN3(n13731), .Q(n5067) );
  nnd4s1 U14023 ( .DIN1(n13732), .DIN2(n13733), .DIN3(n13734), .DIN4(n13735), 
        .Q(n13731) );
  and3s1 U14024 ( .DIN1(n13736), .DIN2(n13737), .DIN3(n13738), .Q(n13735) );
  nnd2s1 U14025 ( .DIN1(n13301), .DIN2(n13357), .Q(n13733) );
  nnd2s1 U14026 ( .DIN1(n13371), .DIN2(n13490), .Q(n13732) );
  nnd3s1 U14027 ( .DIN1(n13739), .DIN2(n13740), .DIN3(n13741), .Q(n13730) );
  or2s1 U14028 ( .DIN1(n13520), .DIN2(n13287), .Q(n13741) );
  or2s1 U14029 ( .DIN1(n13742), .DIN2(n13743), .Q(n13740) );
  nnd2s1 U14030 ( .DIN1(n13293), .DIN2(n13744), .Q(n13739) );
  nnd3s1 U14031 ( .DIN1(n13745), .DIN2(n13746), .DIN3(n13747), .Q(n13729) );
  nnd2s1 U14032 ( .DIN1(n13279), .DIN2(n13748), .Q(n13747) );
  nnd2s1 U14033 ( .DIN1(n13281), .DIN2(n13749), .Q(n13748) );
  nnd2s1 U14034 ( .DIN1(n13288), .DIN2(n13750), .Q(n13746) );
  nnd2s1 U14035 ( .DIN1(n13751), .DIN2(n13752), .Q(n13750) );
  nnd2s1 U14036 ( .DIN1(n13553), .DIN2(n13753), .Q(n13745) );
  nnd2s1 U14037 ( .DIN1(n13505), .DIN2(n13504), .Q(n13753) );
  hi1s1 U14038 ( .DIN(n13687), .Q(n13691) );
  xor2s1 U14039 ( .DIN1(n5043), .DIN2(n13754), .Q(n13687) );
  xor2s1 U14040 ( .DIN1(w2[6]), .DIN2(n5019), .Q(n13754) );
  hi1s1 U14041 ( .DIN(n13108), .Q(n5019) );
  or3s1 U14042 ( .DIN1(n13755), .DIN2(n13756), .DIN3(n13757), .Q(n13108) );
  nnd4s1 U14043 ( .DIN1(n13758), .DIN2(n13759), .DIN3(n13658), .DIN4(n13760), 
        .Q(n13757) );
  and4s1 U14044 ( .DIN1(n13761), .DIN2(n13762), .DIN3(n13763), .DIN4(n13764), 
        .Q(n13760) );
  nnd2s1 U14045 ( .DIN1(n13455), .DIN2(n13765), .Q(n13764) );
  nnd2s1 U14046 ( .DIN1(n13440), .DIN2(n13678), .Q(n13763) );
  nnd2s1 U14047 ( .DIN1(n13766), .DIN2(n13424), .Q(n13762) );
  nor2s1 U14048 ( .DIN1(n13767), .DIN2(n13768), .Q(n13658) );
  nnd4s1 U14049 ( .DIN1(n13769), .DIN2(n13770), .DIN3(n13771), .DIN4(n13772), 
        .Q(n13768) );
  nnd2s1 U14050 ( .DIN1(n13773), .DIN2(n13774), .Q(n13772) );
  nnd3s1 U14051 ( .DIN1(n13673), .DIN2(n13681), .DIN3(n13775), .Q(n13774) );
  nnd2s1 U14052 ( .DIN1(n13776), .DIN2(n13458), .Q(n13771) );
  nnd2s1 U14053 ( .DIN1(n13428), .DIN2(n13777), .Q(n13770) );
  nnd2s1 U14054 ( .DIN1(n13440), .DIN2(n13778), .Q(n13769) );
  nnd4s1 U14055 ( .DIN1(n13779), .DIN2(n13780), .DIN3(n13781), .DIN4(n13782), 
        .Q(n13767) );
  nnd2s1 U14056 ( .DIN1(n13783), .DIN2(n13784), .Q(n13782) );
  nnd2s1 U14057 ( .DIN1(n13785), .DIN2(n13786), .Q(n13784) );
  nnd2s1 U14058 ( .DIN1(n13787), .DIN2(n13788), .Q(n13781) );
  nnd2s1 U14059 ( .DIN1(n13789), .DIN2(n13681), .Q(n13788) );
  nnd2s1 U14060 ( .DIN1(n13424), .DIN2(n13790), .Q(n13780) );
  nnd2s1 U14061 ( .DIN1(n13445), .DIN2(n13791), .Q(n13790) );
  nnd2s1 U14062 ( .DIN1(n13456), .DIN2(n13792), .Q(n13779) );
  nnd2s1 U14063 ( .DIN1(n13793), .DIN2(n13677), .Q(n13792) );
  nnd4s1 U14064 ( .DIN1(n13794), .DIN2(n13795), .DIN3(n13796), .DIN4(n13797), 
        .Q(n13756) );
  nnd2s1 U14065 ( .DIN1(n13431), .DIN2(n13447), .Q(n13797) );
  nnd2s1 U14066 ( .DIN1(n13776), .DIN2(n13798), .Q(n13796) );
  nnd2s1 U14067 ( .DIN1(n13659), .DIN2(n13458), .Q(n13795) );
  nnd2s1 U14068 ( .DIN1(n13428), .DIN2(n13799), .Q(n13794) );
  nnd4s1 U14069 ( .DIN1(n13800), .DIN2(n13801), .DIN3(n13802), .DIN4(n13803), 
        .Q(n13755) );
  nnd2s1 U14070 ( .DIN1(n13429), .DIN2(n13804), .Q(n13803) );
  nnd2s1 U14071 ( .DIN1(n13805), .DIN2(n13806), .Q(n13804) );
  nnd2s1 U14072 ( .DIN1(n13807), .DIN2(n13808), .Q(n13802) );
  nnd2s1 U14073 ( .DIN1(n13438), .DIN2(n13444), .Q(n13808) );
  nnd2s1 U14074 ( .DIN1(n13426), .DIN2(n13809), .Q(n13801) );
  nnd2s1 U14075 ( .DIN1(n13660), .DIN2(n13810), .Q(n13800) );
  or3s1 U14076 ( .DIN1(n13811), .DIN2(n13812), .DIN3(n13813), .Q(n5043) );
  nnd4s1 U14077 ( .DIN1(n13814), .DIN2(n13815), .DIN3(n13816), .DIN4(n13817), 
        .Q(n13813) );
  and3s1 U14078 ( .DIN1(n13818), .DIN2(n13819), .DIN3(n13820), .Q(n13817) );
  nnd2s1 U14079 ( .DIN1(n13181), .DIN2(n13247), .Q(n13815) );
  nnd2s1 U14080 ( .DIN1(n13261), .DIN2(n13579), .Q(n13814) );
  nnd3s1 U14081 ( .DIN1(n13821), .DIN2(n13822), .DIN3(n13823), .Q(n13812) );
  or2s1 U14082 ( .DIN1(n13609), .DIN2(n13167), .Q(n13823) );
  or2s1 U14083 ( .DIN1(n13824), .DIN2(n13825), .Q(n13822) );
  nnd2s1 U14084 ( .DIN1(n13173), .DIN2(n13826), .Q(n13821) );
  nnd3s1 U14085 ( .DIN1(n13827), .DIN2(n13828), .DIN3(n13829), .Q(n13811) );
  nnd2s1 U14086 ( .DIN1(n13159), .DIN2(n13830), .Q(n13829) );
  nnd2s1 U14087 ( .DIN1(n13161), .DIN2(n13831), .Q(n13830) );
  nnd2s1 U14088 ( .DIN1(n13168), .DIN2(n13832), .Q(n13828) );
  nnd2s1 U14089 ( .DIN1(n13833), .DIN2(n13834), .Q(n13832) );
  nnd2s1 U14090 ( .DIN1(n13642), .DIN2(n13835), .Q(n13827) );
  nnd2s1 U14091 ( .DIN1(n13594), .DIN2(n13593), .Q(n13835) );
  nnd2s1 U14092 ( .DIN1(n13836), .DIN2(n13837), .Q(N103) );
  nnd2s1 U14093 ( .DIN1(n13838), .DIN2(n1638), .Q(n13837) );
  xor2s1 U14094 ( .DIN1(n13839), .DIN2(n13840), .Q(n13838) );
  xnr2s1 U14095 ( .DIN1(n5418), .DIN2(n12928), .Q(n13840) );
  xnr2s1 U14096 ( .DIN1(n13695), .DIN2(n5066), .Q(n12928) );
  nor3s1 U14097 ( .DIN1(n13841), .DIN2(n13842), .DIN3(n13843), .Q(n5066) );
  nnd4s1 U14098 ( .DIN1(n13844), .DIN2(n13845), .DIN3(n13738), .DIN4(n13846), 
        .Q(n13843) );
  and4s1 U14099 ( .DIN1(n13847), .DIN2(n13848), .DIN3(n13849), .DIN4(n13850), 
        .Q(n13846) );
  nnd2s1 U14100 ( .DIN1(n13291), .DIN2(n13480), .Q(n13850) );
  nnd2s1 U14101 ( .DIN1(n13290), .DIN2(n13553), .Q(n13849) );
  nnd2s1 U14102 ( .DIN1(n13283), .DIN2(n13279), .Q(n13848) );
  nor2s1 U14103 ( .DIN1(n13851), .DIN2(n13852), .Q(n13738) );
  nnd4s1 U14104 ( .DIN1(n13853), .DIN2(n13854), .DIN3(n13855), .DIN4(n13856), 
        .Q(n13852) );
  nnd2s1 U14105 ( .DIN1(n13548), .DIN2(n13857), .Q(n13856) );
  nnd3s1 U14106 ( .DIN1(n13504), .DIN2(n13557), .DIN3(n13559), .Q(n13857) );
  nnd2s1 U14107 ( .DIN1(n13539), .DIN2(n13341), .Q(n13855) );
  nnd2s1 U14108 ( .DIN1(n13301), .DIN2(n13290), .Q(n13854) );
  nnd2s1 U14109 ( .DIN1(n13500), .DIN2(n13342), .Q(n13853) );
  nnd4s1 U14110 ( .DIN1(n13858), .DIN2(n13859), .DIN3(n13860), .DIN4(n13861), 
        .Q(n13851) );
  nnd2s1 U14111 ( .DIN1(n13357), .DIN2(n13862), .Q(n13861) );
  nnd2s1 U14112 ( .DIN1(n13863), .DIN2(n13368), .Q(n13862) );
  nnd2s1 U14113 ( .DIN1(n13283), .DIN2(n13864), .Q(n13860) );
  nnd2s1 U14114 ( .DIN1(n13329), .DIN2(n13865), .Q(n13864) );
  nnd2s1 U14115 ( .DIN1(n13304), .DIN2(n13866), .Q(n13859) );
  nnd2s1 U14116 ( .DIN1(n13504), .DIN2(n13326), .Q(n13866) );
  nnd2s1 U14117 ( .DIN1(n13306), .DIN2(n13867), .Q(n13858) );
  nnd2s1 U14118 ( .DIN1(n13749), .DIN2(n13519), .Q(n13867) );
  nnd4s1 U14119 ( .DIN1(n13868), .DIN2(n13869), .DIN3(n13870), .DIN4(n13871), 
        .Q(n13842) );
  nnd2s1 U14120 ( .DIN1(n13371), .DIN2(n13872), .Q(n13871) );
  nnd2s1 U14121 ( .DIN1(n13293), .DIN2(n13304), .Q(n13870) );
  nnd2s1 U14122 ( .DIN1(n13353), .DIN2(n13341), .Q(n13869) );
  nnd2s1 U14123 ( .DIN1(n13342), .DIN2(n13490), .Q(n13868) );
  nnd4s1 U14124 ( .DIN1(n13873), .DIN2(n13874), .DIN3(n13875), .DIN4(n13876), 
        .Q(n13841) );
  nnd2s1 U14125 ( .DIN1(n13369), .DIN2(n13877), .Q(n13876) );
  nnd2s1 U14126 ( .DIN1(n13489), .DIN2(n13878), .Q(n13875) );
  nnd2s1 U14127 ( .DIN1(n13281), .DIN2(n13328), .Q(n13878) );
  nnd2s1 U14128 ( .DIN1(n13301), .DIN2(n13879), .Q(n13874) );
  nnd2s1 U14129 ( .DIN1(n13520), .DIN2(n13555), .Q(n13879) );
  nnd2s1 U14130 ( .DIN1(n13331), .DIN2(n13327), .Q(n13873) );
  or3s1 U14131 ( .DIN1(n13880), .DIN2(n13881), .DIN3(n13882), .Q(n13695) );
  nnd4s1 U14132 ( .DIN1(n13883), .DIN2(n13884), .DIN3(n13705), .DIN4(n13885), 
        .Q(n13882) );
  and4s1 U14133 ( .DIN1(n13886), .DIN2(n13887), .DIN3(n13888), .DIN4(n13889), 
        .Q(n13885) );
  nnd2s1 U14134 ( .DIN1(n13412), .DIN2(n13890), .Q(n13889) );
  nnd2s1 U14135 ( .DIN1(n13397), .DIN2(n13725), .Q(n13888) );
  nnd2s1 U14136 ( .DIN1(n13891), .DIN2(n13381), .Q(n13887) );
  nor2s1 U14137 ( .DIN1(n13892), .DIN2(n13893), .Q(n13705) );
  nnd4s1 U14138 ( .DIN1(n13894), .DIN2(n13895), .DIN3(n13896), .DIN4(n13897), 
        .Q(n13893) );
  nnd2s1 U14139 ( .DIN1(n13898), .DIN2(n13899), .Q(n13897) );
  nnd3s1 U14140 ( .DIN1(n13728), .DIN2(n13720), .DIN3(n13900), .Q(n13899) );
  nnd2s1 U14141 ( .DIN1(n13901), .DIN2(n13415), .Q(n13896) );
  nnd2s1 U14142 ( .DIN1(n13902), .DIN2(n13385), .Q(n13895) );
  nnd2s1 U14143 ( .DIN1(n13903), .DIN2(n13397), .Q(n13894) );
  nnd4s1 U14144 ( .DIN1(n13904), .DIN2(n13905), .DIN3(n13906), .DIN4(n13907), 
        .Q(n13892) );
  nnd2s1 U14145 ( .DIN1(n13908), .DIN2(n13909), .Q(n13907) );
  nnd2s1 U14146 ( .DIN1(n13910), .DIN2(n13911), .Q(n13909) );
  nnd2s1 U14147 ( .DIN1(n13912), .DIN2(n13913), .Q(n13906) );
  nnd2s1 U14148 ( .DIN1(n13914), .DIN2(n13728), .Q(n13913) );
  nnd2s1 U14149 ( .DIN1(n13381), .DIN2(n13915), .Q(n13905) );
  nnd2s1 U14150 ( .DIN1(n13402), .DIN2(n13916), .Q(n13915) );
  nnd2s1 U14151 ( .DIN1(n13413), .DIN2(n13917), .Q(n13904) );
  nnd2s1 U14152 ( .DIN1(n13918), .DIN2(n13724), .Q(n13917) );
  nnd4s1 U14153 ( .DIN1(n13919), .DIN2(n13920), .DIN3(n13921), .DIN4(n13922), 
        .Q(n13881) );
  nnd2s1 U14154 ( .DIN1(n13387), .DIN2(n13404), .Q(n13922) );
  nnd2s1 U14155 ( .DIN1(n13901), .DIN2(n13923), .Q(n13921) );
  nnd2s1 U14156 ( .DIN1(n13415), .DIN2(n13707), .Q(n13920) );
  nnd2s1 U14157 ( .DIN1(n13385), .DIN2(n13924), .Q(n13919) );
  nnd4s1 U14158 ( .DIN1(n13925), .DIN2(n13926), .DIN3(n13927), .DIN4(n13928), 
        .Q(n13880) );
  nnd2s1 U14159 ( .DIN1(n13386), .DIN2(n13929), .Q(n13928) );
  nnd2s1 U14160 ( .DIN1(n13930), .DIN2(n13931), .Q(n13929) );
  nnd2s1 U14161 ( .DIN1(n13932), .DIN2(n13933), .Q(n13927) );
  nnd2s1 U14162 ( .DIN1(n13395), .DIN2(n13401), .Q(n13933) );
  nnd2s1 U14163 ( .DIN1(n13383), .DIN2(n13934), .Q(n13926) );
  nnd2s1 U14164 ( .DIN1(n13706), .DIN2(n13935), .Q(n13925) );
  xor2s1 U14165 ( .DIN1(n13027), .DIN2(n13936), .Q(n13839) );
  xor2s1 U14166 ( .DIN1(n1462), .DIN2(n5018), .Q(n13936) );
  or3s1 U14167 ( .DIN1(n13937), .DIN2(n13938), .DIN3(n13939), .Q(n5018) );
  nnd4s1 U14168 ( .DIN1(n13940), .DIN2(n13941), .DIN3(n13942), .DIN4(n13943), 
        .Q(n13939) );
  and4s1 U14169 ( .DIN1(n13944), .DIN2(n13945), .DIN3(n13946), .DIN4(n13947), 
        .Q(n13943) );
  nnd2s1 U14170 ( .DIN1(n13659), .DIN2(n13948), .Q(n13947) );
  nnd2s1 U14171 ( .DIN1(n13442), .DIN2(n13949), .Q(n13948) );
  nnd2s1 U14172 ( .DIN1(n13950), .DIN2(n13951), .Q(n13946) );
  nnd2s1 U14173 ( .DIN1(n13438), .DIN2(n13789), .Q(n13951) );
  nnd2s1 U14174 ( .DIN1(n13678), .DIN2(n13952), .Q(n13945) );
  nnd2s1 U14175 ( .DIN1(n13953), .DIN2(n13677), .Q(n13952) );
  nnd2s1 U14176 ( .DIN1(n13954), .DIN2(n13955), .Q(n13944) );
  nnd2s1 U14177 ( .DIN1(n13956), .DIN2(n13957), .Q(n13955) );
  nnd2s1 U14178 ( .DIN1(n13428), .DIN2(n13958), .Q(n13942) );
  nnd2s1 U14179 ( .DIN1(n13660), .DIN2(n13447), .Q(n13941) );
  nnd2s1 U14180 ( .DIN1(n13789), .DIN2(n13677), .Q(n13447) );
  nnd2s1 U14181 ( .DIN1(n13424), .DIN2(n13798), .Q(n13940) );
  nnd3s1 U14182 ( .DIN1(n13758), .DIN2(n13959), .DIN3(n13656), .Q(n13938) );
  nor4s1 U14183 ( .DIN1(n13960), .DIN2(n13961), .DIN3(n13962), .DIN4(n13963), 
        .Q(n13656) );
  nnd4s1 U14184 ( .DIN1(n13964), .DIN2(n13965), .DIN3(n13966), .DIN4(n13967), 
        .Q(n13963) );
  nnd2s1 U14185 ( .DIN1(n13787), .DIN2(n13783), .Q(n13967) );
  nnd2s1 U14186 ( .DIN1(n13456), .DIN2(n13968), .Q(n13966) );
  nnd2s1 U14187 ( .DIN1(n13807), .DIN2(n13457), .Q(n13965) );
  nnd2s1 U14188 ( .DIN1(n13428), .DIN2(n13969), .Q(n13964) );
  nnd3s1 U14189 ( .DIN1(n13970), .DIN2(n13971), .DIN3(n13972), .Q(n13962) );
  nnd2s1 U14190 ( .DIN1(n13440), .DIN2(n13973), .Q(n13972) );
  nnd2s1 U14191 ( .DIN1(n13785), .DIN2(n13806), .Q(n13973) );
  nnd2s1 U14192 ( .DIN1(n13659), .DIN2(n13974), .Q(n13971) );
  nnd2s1 U14193 ( .DIN1(n13431), .DIN2(n13975), .Q(n13970) );
  nnd2s1 U14194 ( .DIN1(n13976), .DIN2(n13674), .Q(n13975) );
  nor2s1 U14195 ( .DIN1(n13977), .DIN2(n13443), .Q(n13961) );
  and2s1 U14196 ( .DIN1(n13778), .DIN2(n13978), .Q(n13960) );
  nnd3s1 U14197 ( .DIN1(n13681), .DIN2(n13953), .DIN3(n13438), .Q(n13978) );
  nor3s1 U14198 ( .DIN1(n13979), .DIN2(n13980), .DIN3(n13981), .Q(n13758) );
  nnd4s1 U14199 ( .DIN1(n13982), .DIN2(n13983), .DIN3(n13657), .DIN4(n13984), 
        .Q(n13981) );
  and3s1 U14200 ( .DIN1(n13985), .DIN2(n13986), .DIN3(n13987), .Q(n13984) );
  nnd2s1 U14201 ( .DIN1(n13440), .DIN2(n13458), .Q(n13986) );
  nnd2s1 U14202 ( .DIN1(n13424), .DIN2(n13807), .Q(n13985) );
  nor2s1 U14203 ( .DIN1(n13988), .DIN2(n13989), .Q(n13657) );
  nnd4s1 U14204 ( .DIN1(n13990), .DIN2(n13991), .DIN3(n13992), .DIN4(n13993), 
        .Q(n13989) );
  nnd2s1 U14205 ( .DIN1(n13766), .DIN2(n13994), .Q(n13993) );
  nnd2s1 U14206 ( .DIN1(n13429), .DIN2(n13995), .Q(n13992) );
  nnd2s1 U14207 ( .DIN1(n13950), .DIN2(n13958), .Q(n13991) );
  nnd2s1 U14208 ( .DIN1(n13773), .DIN2(n13783), .Q(n13990) );
  nnd4s1 U14209 ( .DIN1(n13996), .DIN2(n13997), .DIN3(n13998), .DIN4(n13999), 
        .Q(n13988) );
  nnd2s1 U14210 ( .DIN1(n13659), .DIN2(n13995), .Q(n13999) );
  nnd2s1 U14211 ( .DIN1(n13455), .DIN2(n14000), .Q(n13998) );
  nnd2s1 U14212 ( .DIN1(n13442), .DIN2(n13957), .Q(n14000) );
  nnd2s1 U14213 ( .DIN1(n13787), .DIN2(n14001), .Q(n13997) );
  nnd2s1 U14214 ( .DIN1(n13793), .DIN2(n13680), .Q(n14001) );
  nnd2s1 U14215 ( .DIN1(n13430), .DIN2(n14002), .Q(n13996) );
  nnd3s1 U14216 ( .DIN1(n14003), .DIN2(n13949), .DIN3(n14004), .Q(n14002) );
  nnd3s1 U14217 ( .DIN1(n14005), .DIN2(n14006), .DIN3(n14007), .Q(n13980) );
  nnd2s1 U14218 ( .DIN1(n13430), .DIN2(n13436), .Q(n14007) );
  nnd2s1 U14219 ( .DIN1(n13455), .DIN2(n14008), .Q(n14006) );
  nnd3s1 U14220 ( .DIN1(n13443), .DIN2(n13791), .DIN3(n13668), .Q(n14008) );
  nor2s1 U14221 ( .DIN1(n13436), .DIN2(n13426), .Q(n13668) );
  nnd2s1 U14222 ( .DIN1(n13446), .DIN2(n13776), .Q(n14005) );
  nnd3s1 U14223 ( .DIN1(n14009), .DIN2(n14010), .DIN3(n14011), .Q(n13979) );
  nnd2s1 U14224 ( .DIN1(n13766), .DIN2(n14012), .Q(n14011) );
  nnd2s1 U14225 ( .DIN1(n13977), .DIN2(n13680), .Q(n14012) );
  nnd2s1 U14226 ( .DIN1(n13431), .DIN2(n14013), .Q(n14010) );
  nnd2s1 U14227 ( .DIN1(n13439), .DIN2(n13444), .Q(n14013) );
  nnd2s1 U14228 ( .DIN1(n13660), .DIN2(n14014), .Q(n14009) );
  nnd2s1 U14229 ( .DIN1(n13793), .DIN2(n13439), .Q(n14014) );
  nnd3s1 U14230 ( .DIN1(n13454), .DIN2(n14015), .DIN3(n14016), .Q(n13937) );
  nnd2s1 U14231 ( .DIN1(n13765), .DIN2(n14017), .Q(n13454) );
  or3s1 U14232 ( .DIN1(n14018), .DIN2(n14019), .DIN3(n14020), .Q(n13027) );
  nnd4s1 U14233 ( .DIN1(n14021), .DIN2(n14022), .DIN3(n13820), .DIN4(n14023), 
        .Q(n14020) );
  and4s1 U14234 ( .DIN1(n14024), .DIN2(n14025), .DIN3(n14026), .DIN4(n14027), 
        .Q(n14023) );
  nnd2s1 U14235 ( .DIN1(n13171), .DIN2(n13569), .Q(n14027) );
  nnd2s1 U14236 ( .DIN1(n13170), .DIN2(n13642), .Q(n14026) );
  nnd2s1 U14237 ( .DIN1(n13163), .DIN2(n13159), .Q(n14025) );
  nor2s1 U14238 ( .DIN1(n14028), .DIN2(n14029), .Q(n13820) );
  nnd4s1 U14239 ( .DIN1(n14030), .DIN2(n14031), .DIN3(n14032), .DIN4(n14033), 
        .Q(n14029) );
  nnd2s1 U14240 ( .DIN1(n13637), .DIN2(n14034), .Q(n14033) );
  nnd3s1 U14241 ( .DIN1(n13593), .DIN2(n13646), .DIN3(n13648), .Q(n14034) );
  nnd2s1 U14242 ( .DIN1(n13628), .DIN2(n13231), .Q(n14032) );
  nnd2s1 U14243 ( .DIN1(n13181), .DIN2(n13170), .Q(n14031) );
  nnd2s1 U14244 ( .DIN1(n13589), .DIN2(n13232), .Q(n14030) );
  nnd4s1 U14245 ( .DIN1(n14035), .DIN2(n14036), .DIN3(n14037), .DIN4(n14038), 
        .Q(n14028) );
  nnd2s1 U14246 ( .DIN1(n13247), .DIN2(n14039), .Q(n14038) );
  nnd2s1 U14247 ( .DIN1(n14040), .DIN2(n13258), .Q(n14039) );
  nnd2s1 U14248 ( .DIN1(n13163), .DIN2(n14041), .Q(n14037) );
  nnd2s1 U14249 ( .DIN1(n13219), .DIN2(n14042), .Q(n14041) );
  nnd2s1 U14250 ( .DIN1(n13184), .DIN2(n14043), .Q(n14036) );
  nnd2s1 U14251 ( .DIN1(n13593), .DIN2(n13216), .Q(n14043) );
  nnd2s1 U14252 ( .DIN1(n13186), .DIN2(n14044), .Q(n14035) );
  nnd2s1 U14253 ( .DIN1(n13831), .DIN2(n13608), .Q(n14044) );
  nnd4s1 U14254 ( .DIN1(n14045), .DIN2(n14046), .DIN3(n14047), .DIN4(n14048), 
        .Q(n14019) );
  nnd2s1 U14255 ( .DIN1(n13261), .DIN2(n14049), .Q(n14048) );
  nnd2s1 U14256 ( .DIN1(n13173), .DIN2(n13184), .Q(n14047) );
  nnd2s1 U14257 ( .DIN1(n13243), .DIN2(n13231), .Q(n14046) );
  nnd2s1 U14258 ( .DIN1(n13232), .DIN2(n13579), .Q(n14045) );
  nnd4s1 U14259 ( .DIN1(n14050), .DIN2(n14051), .DIN3(n14052), .DIN4(n14053), 
        .Q(n14018) );
  nnd2s1 U14260 ( .DIN1(n13259), .DIN2(n14054), .Q(n14053) );
  nnd2s1 U14261 ( .DIN1(n13578), .DIN2(n14055), .Q(n14052) );
  nnd2s1 U14262 ( .DIN1(n13161), .DIN2(n13218), .Q(n14055) );
  nnd2s1 U14263 ( .DIN1(n13181), .DIN2(n14056), .Q(n14051) );
  nnd2s1 U14264 ( .DIN1(n13609), .DIN2(n13644), .Q(n14056) );
  nnd2s1 U14265 ( .DIN1(n13221), .DIN2(n13217), .Q(n14050) );
  nnd2s1 U14266 ( .DIN1(n14057), .DIN2(n1601), .Q(n13836) );
  xor2s1 U14267 ( .DIN1(w2[5]), .DIN2(text_in_r[37]), .Q(n14057) );
  nnd2s1 U14268 ( .DIN1(n14058), .DIN2(n14059), .Q(N102) );
  nnd2s1 U14269 ( .DIN1(n14060), .DIN2(n1637), .Q(n14059) );
  xor2s1 U14270 ( .DIN1(n14061), .DIN2(n14062), .Q(n14060) );
  xor2s1 U14271 ( .DIN1(n12936), .DIN2(n14063), .Q(n14062) );
  xor2s1 U14272 ( .DIN1(n5417), .DIN2(n4739), .Q(n14063) );
  xnr2s1 U14273 ( .DIN1(n5418), .DIN2(n5065), .Q(n12936) );
  hi1s1 U14274 ( .DIN(n13044), .Q(n5065) );
  or3s1 U14275 ( .DIN1(n14064), .DIN2(n14065), .DIN3(n14066), .Q(n13044) );
  nnd4s1 U14276 ( .DIN1(n14067), .DIN2(n14068), .DIN3(n14069), .DIN4(n14070), 
        .Q(n14066) );
  and4s1 U14277 ( .DIN1(n14071), .DIN2(n14072), .DIN3(n14073), .DIN4(n14074), 
        .Q(n14070) );
  nnd2s1 U14278 ( .DIN1(n13359), .DIN2(n14075), .Q(n14074) );
  nnd2s1 U14279 ( .DIN1(n13281), .DIN2(n13326), .Q(n14075) );
  nnd2s1 U14280 ( .DIN1(n13490), .DIN2(n14076), .Q(n14073) );
  nnd2s1 U14281 ( .DIN1(n13502), .DIN2(n13277), .Q(n14076) );
  nnd2s1 U14282 ( .DIN1(n13275), .DIN2(n14077), .Q(n14072) );
  nnd2s1 U14283 ( .DIN1(n14078), .DIN2(n13286), .Q(n14077) );
  nnd2s1 U14284 ( .DIN1(n13553), .DIN2(n14079), .Q(n14071) );
  nnd2s1 U14285 ( .DIN1(n13749), .DIN2(n14080), .Q(n14079) );
  nnd2s1 U14286 ( .DIN1(n13341), .DIN2(n13372), .Q(n14069) );
  nnd2s1 U14287 ( .DIN1(n13371), .DIN2(n13327), .Q(n14068) );
  nnd2s1 U14288 ( .DIN1(n13749), .DIN2(n13326), .Q(n13327) );
  or2s1 U14289 ( .DIN1(n13499), .DIN2(n14081), .Q(n14067) );
  nnd3s1 U14290 ( .DIN1(n13844), .DIN2(n14082), .DIN3(n13736), .Q(n14065) );
  nor4s1 U14291 ( .DIN1(n14083), .DIN2(n14084), .DIN3(n14085), .DIN4(n14086), 
        .Q(n13736) );
  nnd4s1 U14292 ( .DIN1(n14087), .DIN2(n14088), .DIN3(n14089), .DIN4(n14090), 
        .Q(n14086) );
  nnd2s1 U14293 ( .DIN1(n13302), .DIN2(n13341), .Q(n14090) );
  nnd2s1 U14294 ( .DIN1(n13290), .DIN2(n13288), .Q(n14089) );
  nnd2s1 U14295 ( .DIN1(n13306), .DIN2(n13303), .Q(n14088) );
  nnd2s1 U14296 ( .DIN1(n13305), .DIN2(n13489), .Q(n14087) );
  nnd3s1 U14297 ( .DIN1(n14091), .DIN2(n14092), .DIN3(n14093), .Q(n14085) );
  nnd2s1 U14298 ( .DIN1(n13304), .DIN2(n14094), .Q(n14093) );
  nnd2s1 U14299 ( .DIN1(n13282), .DIN2(n13324), .Q(n14094) );
  nnd2s1 U14300 ( .DIN1(n13331), .DIN2(n14095), .Q(n14092) );
  nnd2s1 U14301 ( .DIN1(n14096), .DIN2(n13499), .Q(n14095) );
  nnd2s1 U14302 ( .DIN1(n13548), .DIN2(n14097), .Q(n14091) );
  nnd2s1 U14303 ( .DIN1(n14098), .DIN2(n13328), .Q(n14097) );
  nor2s1 U14304 ( .DIN1(n13558), .DIN2(n13328), .Q(n14084) );
  and2s1 U14305 ( .DIN1(n13301), .DIN2(n14099), .Q(n14083) );
  nnd3s1 U14306 ( .DIN1(n13281), .DIN2(n14080), .DIN3(n13504), .Q(n14099) );
  nor3s1 U14307 ( .DIN1(n14100), .DIN2(n14101), .DIN3(n14102), .Q(n13844) );
  nnd4s1 U14308 ( .DIN1(n14103), .DIN2(n14104), .DIN3(n13737), .DIN4(n14105), 
        .Q(n14102) );
  and3s1 U14309 ( .DIN1(n14106), .DIN2(n14107), .DIN3(n13477), .Q(n14105) );
  nnd2s1 U14310 ( .DIN1(n13539), .DIN2(n13306), .Q(n13477) );
  nnd2s1 U14311 ( .DIN1(n13330), .DIN2(n13288), .Q(n14107) );
  nnd2s1 U14312 ( .DIN1(n13489), .DIN2(n13283), .Q(n14106) );
  nor2s1 U14313 ( .DIN1(n14108), .DIN2(n14109), .Q(n13737) );
  nnd4s1 U14314 ( .DIN1(n14110), .DIN2(n14111), .DIN3(n14112), .DIN4(n14113), 
        .Q(n14109) );
  nnd2s1 U14315 ( .DIN1(n13279), .DIN2(n13537), .Q(n14113) );
  nnd2s1 U14316 ( .DIN1(n13326), .DIN2(n13324), .Q(n13537) );
  nnd2s1 U14317 ( .DIN1(n13293), .DIN2(n13512), .Q(n14112) );
  nnd2s1 U14318 ( .DIN1(n13359), .DIN2(n13372), .Q(n14111) );
  nnd2s1 U14319 ( .DIN1(n13749), .DIN2(n13520), .Q(n13372) );
  nnd2s1 U14320 ( .DIN1(n13548), .DIN2(n13357), .Q(n14110) );
  nnd4s1 U14321 ( .DIN1(n14114), .DIN2(n14115), .DIN3(n14116), .DIN4(n14117), 
        .Q(n14108) );
  nnd2s1 U14322 ( .DIN1(n13490), .DIN2(n13512), .Q(n14117) );
  nnd2s1 U14323 ( .DIN1(n13480), .DIN2(n14118), .Q(n14116) );
  nnd2s1 U14324 ( .DIN1(n13502), .DIN2(n13286), .Q(n14118) );
  nnd2s1 U14325 ( .DIN1(n13304), .DIN2(n14119), .Q(n14115) );
  nnd2s1 U14326 ( .DIN1(n13505), .DIN2(n13519), .Q(n14119) );
  nnd2s1 U14327 ( .DIN1(n13330), .DIN2(n14120), .Q(n14114) );
  nnd3s1 U14328 ( .DIN1(n13277), .DIN2(n13558), .DIN3(n13285), .Q(n14120) );
  nnd3s1 U14329 ( .DIN1(n14121), .DIN2(n14122), .DIN3(n14123), .Q(n14101) );
  nnd2s1 U14330 ( .DIN1(n13290), .DIN2(n13342), .Q(n14123) );
  nnd2s1 U14331 ( .DIN1(n13480), .DIN2(n14124), .Q(n14122) );
  nnd3s1 U14332 ( .DIN1(n13366), .DIN2(n13865), .DIN3(n13743), .Q(n14124) );
  nor2s1 U14333 ( .DIN1(n13369), .DIN2(n13288), .Q(n13743) );
  nnd2s1 U14334 ( .DIN1(n13292), .DIN2(n13500), .Q(n14121) );
  nnd3s1 U14335 ( .DIN1(n14125), .DIN2(n14126), .DIN3(n14127), .Q(n14100) );
  nnd2s1 U14336 ( .DIN1(n13279), .DIN2(n14128), .Q(n14127) );
  nnd2s1 U14337 ( .DIN1(n14129), .DIN2(n13742), .Q(n14128) );
  nnd2s1 U14338 ( .DIN1(n13331), .DIN2(n14130), .Q(n14126) );
  nnd2s1 U14339 ( .DIN1(n13328), .DIN2(n13324), .Q(n14130) );
  nnd2s1 U14340 ( .DIN1(n13371), .DIN2(n14131), .Q(n14125) );
  nnd2s1 U14341 ( .DIN1(n13519), .DIN2(n13324), .Q(n14131) );
  nnd3s1 U14342 ( .DIN1(n13267), .DIN2(n14132), .DIN3(n14133), .Q(n14064) );
  nnd2s1 U14343 ( .DIN1(n13333), .DIN2(n13291), .Q(n14132) );
  nnd2s1 U14344 ( .DIN1(n13500), .DIN2(n13331), .Q(n13267) );
  or3s1 U14345 ( .DIN1(n14134), .DIN2(n14135), .DIN3(n14136), .Q(n5418) );
  nnd4s1 U14346 ( .DIN1(n14137), .DIN2(n14138), .DIN3(n14139), .DIN4(n14140), 
        .Q(n14136) );
  and4s1 U14347 ( .DIN1(n14141), .DIN2(n14142), .DIN3(n14143), .DIN4(n14144), 
        .Q(n14140) );
  nnd2s1 U14348 ( .DIN1(n13707), .DIN2(n14145), .Q(n14144) );
  nnd2s1 U14349 ( .DIN1(n13399), .DIN2(n14146), .Q(n14145) );
  nnd2s1 U14350 ( .DIN1(n14147), .DIN2(n14148), .Q(n14143) );
  nnd2s1 U14351 ( .DIN1(n13395), .DIN2(n13914), .Q(n14148) );
  nnd2s1 U14352 ( .DIN1(n13725), .DIN2(n14149), .Q(n14142) );
  nnd2s1 U14353 ( .DIN1(n14150), .DIN2(n13724), .Q(n14149) );
  nnd2s1 U14354 ( .DIN1(n14151), .DIN2(n14152), .Q(n14141) );
  nnd2s1 U14355 ( .DIN1(n14153), .DIN2(n14154), .Q(n14152) );
  nnd2s1 U14356 ( .DIN1(n13385), .DIN2(n14155), .Q(n14139) );
  nnd2s1 U14357 ( .DIN1(n13706), .DIN2(n13404), .Q(n14138) );
  nnd2s1 U14358 ( .DIN1(n13914), .DIN2(n13724), .Q(n13404) );
  nnd2s1 U14359 ( .DIN1(n13381), .DIN2(n13923), .Q(n14137) );
  nnd3s1 U14360 ( .DIN1(n13883), .DIN2(n14156), .DIN3(n13703), .Q(n14135) );
  nor4s1 U14361 ( .DIN1(n14157), .DIN2(n14158), .DIN3(n14159), .DIN4(n14160), 
        .Q(n13703) );
  nnd4s1 U14362 ( .DIN1(n14161), .DIN2(n14162), .DIN3(n14163), .DIN4(n14164), 
        .Q(n14160) );
  nnd2s1 U14363 ( .DIN1(n13908), .DIN2(n13912), .Q(n14164) );
  nnd2s1 U14364 ( .DIN1(n13413), .DIN2(n14165), .Q(n14163) );
  nnd2s1 U14365 ( .DIN1(n13414), .DIN2(n13932), .Q(n14162) );
  nnd2s1 U14366 ( .DIN1(n14166), .DIN2(n13385), .Q(n14161) );
  nnd3s1 U14367 ( .DIN1(n14167), .DIN2(n14168), .DIN3(n14169), .Q(n14159) );
  nnd2s1 U14368 ( .DIN1(n13397), .DIN2(n14170), .Q(n14169) );
  nnd2s1 U14369 ( .DIN1(n13910), .DIN2(n13931), .Q(n14170) );
  nnd2s1 U14370 ( .DIN1(n13707), .DIN2(n14171), .Q(n14168) );
  nnd2s1 U14371 ( .DIN1(n13387), .DIN2(n14172), .Q(n14167) );
  nnd2s1 U14372 ( .DIN1(n14173), .DIN2(n13721), .Q(n14172) );
  nor2s1 U14373 ( .DIN1(n14174), .DIN2(n13400), .Q(n14158) );
  and2s1 U14374 ( .DIN1(n13903), .DIN2(n14175), .Q(n14157) );
  nnd3s1 U14375 ( .DIN1(n14150), .DIN2(n13395), .DIN3(n13728), .Q(n14175) );
  nor3s1 U14376 ( .DIN1(n14176), .DIN2(n14177), .DIN3(n14178), .Q(n13883) );
  nnd4s1 U14377 ( .DIN1(n14179), .DIN2(n14180), .DIN3(n13704), .DIN4(n14181), 
        .Q(n14178) );
  and3s1 U14378 ( .DIN1(n14182), .DIN2(n14183), .DIN3(n14184), .Q(n14181) );
  nnd2s1 U14379 ( .DIN1(n13397), .DIN2(n13415), .Q(n14183) );
  nnd2s1 U14380 ( .DIN1(n13932), .DIN2(n13381), .Q(n14182) );
  nor2s1 U14381 ( .DIN1(n14185), .DIN2(n14186), .Q(n13704) );
  nnd4s1 U14382 ( .DIN1(n14187), .DIN2(n14188), .DIN3(n14189), .DIN4(n14190), 
        .Q(n14186) );
  nnd2s1 U14383 ( .DIN1(n13891), .DIN2(n14191), .Q(n14190) );
  nnd2s1 U14384 ( .DIN1(n13386), .DIN2(n14192), .Q(n14189) );
  nnd2s1 U14385 ( .DIN1(n14147), .DIN2(n14155), .Q(n14188) );
  nnd2s1 U14386 ( .DIN1(n13898), .DIN2(n13908), .Q(n14187) );
  nnd4s1 U14387 ( .DIN1(n14193), .DIN2(n14194), .DIN3(n14195), .DIN4(n14196), 
        .Q(n14185) );
  nnd2s1 U14388 ( .DIN1(n13707), .DIN2(n14192), .Q(n14196) );
  nnd2s1 U14389 ( .DIN1(n13412), .DIN2(n14197), .Q(n14195) );
  nnd2s1 U14390 ( .DIN1(n13399), .DIN2(n14154), .Q(n14197) );
  nnd2s1 U14391 ( .DIN1(n13912), .DIN2(n14198), .Q(n14194) );
  nnd2s1 U14392 ( .DIN1(n13918), .DIN2(n13727), .Q(n14198) );
  nnd2s1 U14393 ( .DIN1(n13388), .DIN2(n14199), .Q(n14193) );
  nnd3s1 U14394 ( .DIN1(n14200), .DIN2(n14201), .DIN3(n14146), .Q(n14199) );
  nnd3s1 U14395 ( .DIN1(n14202), .DIN2(n14203), .DIN3(n14204), .Q(n14177) );
  nnd2s1 U14396 ( .DIN1(n13393), .DIN2(n13388), .Q(n14204) );
  nnd2s1 U14397 ( .DIN1(n13412), .DIN2(n14205), .Q(n14203) );
  nnd3s1 U14398 ( .DIN1(n13916), .DIN2(n13400), .DIN3(n13715), .Q(n14205) );
  nor2s1 U14399 ( .DIN1(n13393), .DIN2(n13383), .Q(n13715) );
  nnd2s1 U14400 ( .DIN1(n13403), .DIN2(n13901), .Q(n14202) );
  nnd3s1 U14401 ( .DIN1(n14206), .DIN2(n14207), .DIN3(n14208), .Q(n14176) );
  nnd2s1 U14402 ( .DIN1(n13891), .DIN2(n14209), .Q(n14208) );
  nnd2s1 U14403 ( .DIN1(n14174), .DIN2(n13727), .Q(n14209) );
  nnd2s1 U14404 ( .DIN1(n13387), .DIN2(n14210), .Q(n14207) );
  nnd2s1 U14405 ( .DIN1(n13396), .DIN2(n13401), .Q(n14210) );
  nnd2s1 U14406 ( .DIN1(n13706), .DIN2(n14211), .Q(n14206) );
  nnd2s1 U14407 ( .DIN1(n13918), .DIN2(n13396), .Q(n14211) );
  nnd3s1 U14408 ( .DIN1(n13411), .DIN2(n14212), .DIN3(n14213), .Q(n14134) );
  nnd2s1 U14409 ( .DIN1(n13890), .DIN2(n14214), .Q(n13411) );
  xor2s1 U14410 ( .DIN1(n13115), .DIN2(n14215), .Q(n14061) );
  xor2s1 U14411 ( .DIN1(n1478), .DIN2(n5017), .Q(n14215) );
  or3s1 U14412 ( .DIN1(n14216), .DIN2(n14217), .DIN3(n14218), .Q(n5017) );
  nnd4s1 U14413 ( .DIN1(n14219), .DIN2(n14220), .DIN3(n13654), .DIN4(n14221), 
        .Q(n14218) );
  and3s1 U14414 ( .DIN1(n13759), .DIN2(n13982), .DIN3(n13959), .Q(n14221) );
  nor4s1 U14415 ( .DIN1(n14222), .DIN2(n14223), .DIN3(n14224), .DIN4(n14225), 
        .Q(n13959) );
  nnd4s1 U14416 ( .DIN1(n14226), .DIN2(n14227), .DIN3(n14228), .DIN4(n14229), 
        .Q(n14225) );
  nor2s1 U14417 ( .DIN1(n14230), .DIN2(n14231), .Q(n14229) );
  nor2s1 U14418 ( .DIN1(n14232), .DIN2(n13664), .Q(n14231) );
  nor2s1 U14419 ( .DIN1(n14233), .DIN2(n14234), .Q(n14230) );
  nnd2s1 U14420 ( .DIN1(n13426), .DIN2(n13810), .Q(n14228) );
  nnd2s1 U14421 ( .DIN1(n13446), .DIN2(n14235), .Q(n14227) );
  nnd3s1 U14422 ( .DIN1(n13439), .DIN2(n13667), .DIN3(n13677), .Q(n14235) );
  nnd2s1 U14423 ( .DIN1(n14017), .DIN2(n14236), .Q(n14226) );
  nnd3s1 U14424 ( .DIN1(n14237), .DIN2(n13785), .DIN3(n14003), .Q(n14236) );
  nnd3s1 U14425 ( .DIN1(n14238), .DIN2(n14239), .DIN3(n14240), .Q(n14224) );
  nnd2s1 U14426 ( .DIN1(n13950), .DIN2(n13783), .Q(n14240) );
  nnd2s1 U14427 ( .DIN1(n13456), .DIN2(n13429), .Q(n14239) );
  nnd2s1 U14428 ( .DIN1(n13659), .DIN2(n13428), .Q(n14238) );
  nor2s1 U14429 ( .DIN1(n13438), .DIN2(n14237), .Q(n14223) );
  nor2s1 U14430 ( .DIN1(n13957), .DIN2(n13680), .Q(n14222) );
  nor4s1 U14431 ( .DIN1(n14241), .DIN2(n14242), .DIN3(n14243), .DIN4(n14244), 
        .Q(n13982) );
  nnd4s1 U14432 ( .DIN1(n14245), .DIN2(n14246), .DIN3(n14247), .DIN4(n14248), 
        .Q(n14244) );
  nor2s1 U14433 ( .DIN1(n14249), .DIN2(n14250), .Q(n14248) );
  nor2s1 U14434 ( .DIN1(n14003), .DIN2(n13674), .Q(n14250) );
  nor2s1 U14435 ( .DIN1(n13439), .DIN2(n14251), .Q(n14249) );
  nnd2s1 U14436 ( .DIN1(n13773), .DIN2(n13799), .Q(n14246) );
  nnd3s1 U14437 ( .DIN1(n14252), .DIN2(n14253), .DIN3(n14254), .Q(n14243) );
  nnd2s1 U14438 ( .DIN1(n13458), .DIN2(n14255), .Q(n14254) );
  nnd2s1 U14439 ( .DIN1(n14256), .DIN2(n13439), .Q(n14255) );
  nnd2s1 U14440 ( .DIN1(n13659), .DIN2(n13676), .Q(n14253) );
  nnd2s1 U14441 ( .DIN1(n13787), .DIN2(n13809), .Q(n14252) );
  nnd2s1 U14442 ( .DIN1(n14257), .DIN2(n13673), .Q(n13809) );
  nor2s1 U14443 ( .DIN1(n14258), .DIN2(n13805), .Q(n14242) );
  nor2s1 U14444 ( .DIN1(n13799), .DIN2(n13968), .Q(n14258) );
  nor2s1 U14445 ( .DIN1(n14259), .DIN2(n13438), .Q(n14241) );
  nor2s1 U14446 ( .DIN1(n13446), .DIN2(n13426), .Q(n14259) );
  nor4s1 U14447 ( .DIN1(n14260), .DIN2(n14261), .DIN3(n14262), .DIN4(n14263), 
        .Q(n13759) );
  nnd4s1 U14448 ( .DIN1(n14264), .DIN2(n14265), .DIN3(n14266), .DIN4(n14267), 
        .Q(n14263) );
  nor2s1 U14449 ( .DIN1(n14268), .DIN2(n14269), .Q(n14266) );
  nor2s1 U14450 ( .DIN1(n13786), .DIN2(n13680), .Q(n14269) );
  nor2s1 U14451 ( .DIN1(n13667), .DIN2(n14004), .Q(n14268) );
  nnd2s1 U14452 ( .DIN1(n13428), .DIN2(n13954), .Q(n14265) );
  nnd2s1 U14453 ( .DIN1(n13440), .DIN2(n13456), .Q(n14264) );
  nnd3s1 U14454 ( .DIN1(n14270), .DIN2(n14271), .DIN3(n14272), .Q(n14262) );
  nnd2s1 U14455 ( .DIN1(n13660), .DIN2(n14273), .Q(n14272) );
  nnd2s1 U14456 ( .DIN1(n13458), .DIN2(n14274), .Q(n14271) );
  nnd2s1 U14457 ( .DIN1(n13446), .DIN2(n14275), .Q(n14270) );
  nnd3s1 U14458 ( .DIN1(n13953), .DIN2(n14234), .DIN3(n14276), .Q(n14275) );
  nor2s1 U14459 ( .DIN1(n14277), .DIN2(n13785), .Q(n14261) );
  nor2s1 U14460 ( .DIN1(n14278), .DIN2(n13806), .Q(n14260) );
  and4s1 U14461 ( .DIN1(n13983), .DIN2(n14016), .DIN3(n14279), .DIN4(n14280), 
        .Q(n13654) );
  and4s1 U14462 ( .DIN1(n14281), .DIN2(n14282), .DIN3(n14283), .DIN4(n14284), 
        .Q(n14280) );
  and3s1 U14463 ( .DIN1(n14285), .DIN2(n14286), .DIN3(n14287), .Q(n14284) );
  nnd2s1 U14464 ( .DIN1(n13426), .DIN2(n14288), .Q(n14287) );
  nnd2s1 U14465 ( .DIN1(n13674), .DIN2(n13439), .Q(n14288) );
  nnd2s1 U14466 ( .DIN1(n13773), .DIN2(n14289), .Q(n14286) );
  nnd2s1 U14467 ( .DIN1(n13677), .DIN2(n14277), .Q(n14289) );
  nnd2s1 U14468 ( .DIN1(n13660), .DIN2(n14290), .Q(n14285) );
  nnd2s1 U14469 ( .DIN1(n13673), .DIN2(n14277), .Q(n14290) );
  or2s1 U14470 ( .DIN1(n13793), .DIN2(n14291), .Q(n14283) );
  nnd2s1 U14471 ( .DIN1(n13456), .DIN2(n14292), .Q(n14282) );
  or2s1 U14472 ( .DIN1(n13810), .DIN2(n14017), .Q(n14292) );
  nnd2s1 U14473 ( .DIN1(n13680), .DIN2(n13664), .Q(n13810) );
  nnd2s1 U14474 ( .DIN1(n13457), .DIN2(n14293), .Q(n14281) );
  nnd3s1 U14475 ( .DIN1(n14004), .DIN2(n14237), .DIN3(n14294), .Q(n14293) );
  and3s1 U14476 ( .DIN1(n14295), .DIN2(n14296), .DIN3(n13761), .Q(n14279) );
  nor4s1 U14477 ( .DIN1(n14297), .DIN2(n14298), .DIN3(n14299), .DIN4(n14300), 
        .Q(n13761) );
  nnd4s1 U14478 ( .DIN1(n14301), .DIN2(n14302), .DIN3(n14303), .DIN4(n14304), 
        .Q(n14300) );
  nnd2s1 U14479 ( .DIN1(n13426), .DIN2(n14017), .Q(n14304) );
  nnd2s1 U14480 ( .DIN1(n13954), .DIN2(n13431), .Q(n14303) );
  nnd2s1 U14481 ( .DIN1(n13678), .DIN2(n13777), .Q(n14302) );
  nnd2s1 U14482 ( .DIN1(n13807), .DIN2(n13968), .Q(n14301) );
  nnd3s1 U14483 ( .DIN1(n14305), .DIN2(n14306), .DIN3(n14307), .Q(n14299) );
  nnd2s1 U14484 ( .DIN1(n13436), .DIN2(n14308), .Q(n14307) );
  nnd3s1 U14485 ( .DIN1(n13793), .DIN2(n14257), .DIN3(n13680), .Q(n14308) );
  nnd2s1 U14486 ( .DIN1(n13428), .DIN2(n14309), .Q(n14306) );
  nnd2s1 U14487 ( .DIN1(n14234), .DIN2(n13681), .Q(n14309) );
  nnd2s1 U14488 ( .DIN1(n13765), .DIN2(n14310), .Q(n14305) );
  nnd2s1 U14489 ( .DIN1(n14256), .DIN2(n13793), .Q(n14310) );
  nor2s1 U14490 ( .DIN1(n13457), .DIN2(n14311), .Q(n14256) );
  nor2s1 U14491 ( .DIN1(n13956), .DIN2(n13681), .Q(n14298) );
  nor2s1 U14492 ( .DIN1(n13775), .DIN2(n13957), .Q(n14297) );
  hi1s1 U14493 ( .DIN(n13427), .Q(n13775) );
  nnd2s1 U14494 ( .DIN1(n13455), .DIN2(n13678), .Q(n14296) );
  nnd2s1 U14495 ( .DIN1(n13428), .DIN2(n13968), .Q(n14295) );
  nor4s1 U14496 ( .DIN1(n14312), .DIN2(n14313), .DIN3(n14314), .DIN4(n14315), 
        .Q(n14016) );
  nnd4s1 U14497 ( .DIN1(n14316), .DIN2(n14317), .DIN3(n14318), .DIN4(n14319), 
        .Q(n14315) );
  nnd2s1 U14498 ( .DIN1(n13457), .DIN2(n13995), .Q(n14319) );
  nor2s1 U14499 ( .DIN1(n14320), .DIN2(n14321), .Q(n14318) );
  nor2s1 U14500 ( .DIN1(n14322), .DIN2(n14323), .Q(n14321) );
  nor2s1 U14501 ( .DIN1(n13429), .DIN2(n14017), .Q(n14322) );
  nor2s1 U14502 ( .DIN1(n14324), .DIN2(n13805), .Q(n14320) );
  nor2s1 U14503 ( .DIN1(n13455), .DIN2(n14325), .Q(n14324) );
  nnd2s1 U14504 ( .DIN1(n13954), .DIN2(n14326), .Q(n14317) );
  nnd3s1 U14505 ( .DIN1(n13442), .DIN2(n13786), .DIN3(n14004), .Q(n14326) );
  nnd2s1 U14506 ( .DIN1(n13659), .DIN2(n13787), .Q(n14316) );
  nnd3s1 U14507 ( .DIN1(n14327), .DIN2(n14328), .DIN3(n14329), .Q(n14314) );
  nnd2s1 U14508 ( .DIN1(n13950), .DIN2(n14017), .Q(n14328) );
  nnd2s1 U14509 ( .DIN1(n13426), .DIN2(n14311), .Q(n14327) );
  nor2s1 U14510 ( .DIN1(n13956), .DIN2(n14234), .Q(n14313) );
  nor2s1 U14511 ( .DIN1(n14232), .DIN2(n13674), .Q(n14312) );
  nor2s1 U14512 ( .DIN1(n14330), .DIN2(n14331), .Q(n13983) );
  nnd4s1 U14513 ( .DIN1(n14332), .DIN2(n14333), .DIN3(n14334), .DIN4(n14335), 
        .Q(n14331) );
  nnd2s1 U14514 ( .DIN1(n13968), .DIN2(n14336), .Q(n14335) );
  nnd3s1 U14515 ( .DIN1(n13957), .DIN2(n13786), .DIN3(n14237), .Q(n14336) );
  nnd2s1 U14516 ( .DIN1(n13950), .DIN2(n13424), .Q(n14334) );
  nnd4s1 U14517 ( .DIN1(n14337), .DIN2(n14338), .DIN3(n14339), .DIN4(n14340), 
        .Q(n14330) );
  nnd2s1 U14518 ( .DIN1(n13429), .DIN2(n14341), .Q(n14340) );
  nnd2s1 U14519 ( .DIN1(n13786), .DIN2(n13949), .Q(n14341) );
  nnd2s1 U14520 ( .DIN1(n13430), .DIN2(n14342), .Q(n14339) );
  nnd2s1 U14521 ( .DIN1(n13665), .DIN2(n13442), .Q(n14342) );
  nnd2s1 U14522 ( .DIN1(n13807), .DIN2(n14343), .Q(n14338) );
  nnd2s1 U14523 ( .DIN1(n14344), .DIN2(n13680), .Q(n14343) );
  nnd2s1 U14524 ( .DIN1(n13778), .DIN2(n14345), .Q(n14337) );
  nnd2s1 U14525 ( .DIN1(n13783), .DIN2(n13678), .Q(n14219) );
  nnd3s1 U14526 ( .DIN1(n14346), .DIN2(n14347), .DIN3(n14348), .Q(n14217) );
  nnd2s1 U14527 ( .DIN1(n14311), .DIN2(n13807), .Q(n14348) );
  nnd2s1 U14528 ( .DIN1(n13969), .DIN2(n13425), .Q(n14347) );
  nnd2s1 U14529 ( .DIN1(n13440), .DIN2(n13773), .Q(n14346) );
  nnd4s1 U14530 ( .DIN1(n14349), .DIN2(n14350), .DIN3(n14351), .DIN4(n14352), 
        .Q(n14216) );
  nnd2s1 U14531 ( .DIN1(n13799), .DIN2(n14353), .Q(n14352) );
  nnd2s1 U14532 ( .DIN1(n14004), .DIN2(n13791), .Q(n14353) );
  nnd2s1 U14533 ( .DIN1(n13777), .DIN2(n14354), .Q(n14351) );
  nnd2s1 U14534 ( .DIN1(n13445), .DIN2(n14003), .Q(n14354) );
  nor2s1 U14535 ( .DIN1(n13458), .DIN2(n13773), .Q(n13445) );
  nnd2s1 U14536 ( .DIN1(n13765), .DIN2(n14355), .Q(n14350) );
  nnd2s1 U14537 ( .DIN1(n14278), .DIN2(n13444), .Q(n14355) );
  nor2s1 U14538 ( .DIN1(n13777), .DIN2(n13424), .Q(n14278) );
  nnd2s1 U14539 ( .DIN1(n13954), .DIN2(n13995), .Q(n14349) );
  or3s1 U14540 ( .DIN1(n14356), .DIN2(n14357), .DIN3(n14358), .Q(n13115) );
  nnd4s1 U14541 ( .DIN1(n14359), .DIN2(n14360), .DIN3(n14361), .DIN4(n14362), 
        .Q(n14358) );
  and4s1 U14542 ( .DIN1(n14363), .DIN2(n14364), .DIN3(n14365), .DIN4(n14366), 
        .Q(n14362) );
  nnd2s1 U14543 ( .DIN1(n13249), .DIN2(n14367), .Q(n14366) );
  nnd2s1 U14544 ( .DIN1(n13161), .DIN2(n13216), .Q(n14367) );
  nnd2s1 U14545 ( .DIN1(n13579), .DIN2(n14368), .Q(n14365) );
  nnd2s1 U14546 ( .DIN1(n13591), .DIN2(n13157), .Q(n14368) );
  nnd2s1 U14547 ( .DIN1(n13155), .DIN2(n14369), .Q(n14364) );
  nnd2s1 U14548 ( .DIN1(n14370), .DIN2(n13166), .Q(n14369) );
  nnd2s1 U14549 ( .DIN1(n13642), .DIN2(n14371), .Q(n14363) );
  nnd2s1 U14550 ( .DIN1(n13831), .DIN2(n14372), .Q(n14371) );
  nnd2s1 U14551 ( .DIN1(n13231), .DIN2(n13262), .Q(n14361) );
  nnd2s1 U14552 ( .DIN1(n13261), .DIN2(n13217), .Q(n14360) );
  nnd2s1 U14553 ( .DIN1(n13831), .DIN2(n13216), .Q(n13217) );
  or2s1 U14554 ( .DIN1(n13588), .DIN2(n14373), .Q(n14359) );
  nnd3s1 U14555 ( .DIN1(n14021), .DIN2(n14374), .DIN3(n13818), .Q(n14357) );
  nor4s1 U14556 ( .DIN1(n14375), .DIN2(n14376), .DIN3(n14377), .DIN4(n14378), 
        .Q(n13818) );
  nnd4s1 U14557 ( .DIN1(n14379), .DIN2(n14380), .DIN3(n14381), .DIN4(n14382), 
        .Q(n14378) );
  nnd2s1 U14558 ( .DIN1(n13182), .DIN2(n13231), .Q(n14382) );
  nnd2s1 U14559 ( .DIN1(n13170), .DIN2(n13168), .Q(n14381) );
  nnd2s1 U14560 ( .DIN1(n13186), .DIN2(n13183), .Q(n14380) );
  nnd2s1 U14561 ( .DIN1(n13185), .DIN2(n13578), .Q(n14379) );
  nnd3s1 U14562 ( .DIN1(n14383), .DIN2(n14384), .DIN3(n14385), .Q(n14377) );
  nnd2s1 U14563 ( .DIN1(n13184), .DIN2(n14386), .Q(n14385) );
  nnd2s1 U14564 ( .DIN1(n13162), .DIN2(n13214), .Q(n14386) );
  nnd2s1 U14565 ( .DIN1(n13221), .DIN2(n14387), .Q(n14384) );
  nnd2s1 U14566 ( .DIN1(n14388), .DIN2(n13588), .Q(n14387) );
  nnd2s1 U14567 ( .DIN1(n13637), .DIN2(n14389), .Q(n14383) );
  nnd2s1 U14568 ( .DIN1(n14390), .DIN2(n13218), .Q(n14389) );
  nor2s1 U14569 ( .DIN1(n13647), .DIN2(n13218), .Q(n14376) );
  and2s1 U14570 ( .DIN1(n13181), .DIN2(n14391), .Q(n14375) );
  nnd3s1 U14571 ( .DIN1(n13161), .DIN2(n14372), .DIN3(n13593), .Q(n14391) );
  nor3s1 U14572 ( .DIN1(n14392), .DIN2(n14393), .DIN3(n14394), .Q(n14021) );
  nnd4s1 U14573 ( .DIN1(n14395), .DIN2(n14396), .DIN3(n13819), .DIN4(n14397), 
        .Q(n14394) );
  and3s1 U14574 ( .DIN1(n14398), .DIN2(n14399), .DIN3(n13566), .Q(n14397) );
  nnd2s1 U14575 ( .DIN1(n13628), .DIN2(n13186), .Q(n13566) );
  nnd2s1 U14576 ( .DIN1(n13220), .DIN2(n13168), .Q(n14399) );
  nnd2s1 U14577 ( .DIN1(n13578), .DIN2(n13163), .Q(n14398) );
  nor2s1 U14578 ( .DIN1(n14400), .DIN2(n14401), .Q(n13819) );
  nnd4s1 U14579 ( .DIN1(n14402), .DIN2(n14403), .DIN3(n14404), .DIN4(n14405), 
        .Q(n14401) );
  nnd2s1 U14580 ( .DIN1(n13159), .DIN2(n13626), .Q(n14405) );
  nnd2s1 U14581 ( .DIN1(n13216), .DIN2(n13214), .Q(n13626) );
  nnd2s1 U14582 ( .DIN1(n13173), .DIN2(n13601), .Q(n14404) );
  nnd2s1 U14583 ( .DIN1(n13249), .DIN2(n13262), .Q(n14403) );
  nnd2s1 U14584 ( .DIN1(n13831), .DIN2(n13609), .Q(n13262) );
  nnd2s1 U14585 ( .DIN1(n13637), .DIN2(n13247), .Q(n14402) );
  nnd4s1 U14586 ( .DIN1(n14406), .DIN2(n14407), .DIN3(n14408), .DIN4(n14409), 
        .Q(n14400) );
  nnd2s1 U14587 ( .DIN1(n13579), .DIN2(n13601), .Q(n14409) );
  nnd2s1 U14588 ( .DIN1(n13569), .DIN2(n14410), .Q(n14408) );
  nnd2s1 U14589 ( .DIN1(n13591), .DIN2(n13166), .Q(n14410) );
  nnd2s1 U14590 ( .DIN1(n13184), .DIN2(n14411), .Q(n14407) );
  nnd2s1 U14591 ( .DIN1(n13594), .DIN2(n13608), .Q(n14411) );
  nnd2s1 U14592 ( .DIN1(n13220), .DIN2(n14412), .Q(n14406) );
  nnd3s1 U14593 ( .DIN1(n13157), .DIN2(n13647), .DIN3(n13165), .Q(n14412) );
  nnd3s1 U14594 ( .DIN1(n14413), .DIN2(n14414), .DIN3(n14415), .Q(n14393) );
  nnd2s1 U14595 ( .DIN1(n13170), .DIN2(n13232), .Q(n14415) );
  nnd2s1 U14596 ( .DIN1(n13569), .DIN2(n14416), .Q(n14414) );
  nnd3s1 U14597 ( .DIN1(n13256), .DIN2(n14042), .DIN3(n13825), .Q(n14416) );
  nor2s1 U14598 ( .DIN1(n13259), .DIN2(n13168), .Q(n13825) );
  nnd2s1 U14599 ( .DIN1(n13172), .DIN2(n13589), .Q(n14413) );
  nnd3s1 U14600 ( .DIN1(n14417), .DIN2(n14418), .DIN3(n14419), .Q(n14392) );
  nnd2s1 U14601 ( .DIN1(n13159), .DIN2(n14420), .Q(n14419) );
  nnd2s1 U14602 ( .DIN1(n14421), .DIN2(n13824), .Q(n14420) );
  nnd2s1 U14603 ( .DIN1(n13221), .DIN2(n14422), .Q(n14418) );
  nnd2s1 U14604 ( .DIN1(n13218), .DIN2(n13214), .Q(n14422) );
  nnd2s1 U14605 ( .DIN1(n13261), .DIN2(n14423), .Q(n14417) );
  nnd2s1 U14606 ( .DIN1(n13608), .DIN2(n13214), .Q(n14423) );
  nnd3s1 U14607 ( .DIN1(n13147), .DIN2(n14424), .DIN3(n14425), .Q(n14356) );
  nnd2s1 U14608 ( .DIN1(n13223), .DIN2(n13171), .Q(n14424) );
  nnd2s1 U14609 ( .DIN1(n13589), .DIN2(n13221), .Q(n13147) );
  nnd2s1 U14610 ( .DIN1(n14426), .DIN2(n1599), .Q(n14058) );
  xor2s1 U14611 ( .DIN1(w2[4]), .DIN2(text_in_r[36]), .Q(n14426) );
  nnd2s1 U14612 ( .DIN1(n14427), .DIN2(n14428), .Q(N101) );
  nnd2s1 U14613 ( .DIN1(n14429), .DIN2(n1638), .Q(n14428) );
  xor2s1 U14614 ( .DIN1(n14430), .DIN2(n14431), .Q(n14429) );
  xor2s1 U14615 ( .DIN1(n12950), .DIN2(n14432), .Q(n14431) );
  xor2s1 U14616 ( .DIN1(n13070), .DIN2(n4739), .Q(n14432) );
  hi1s1 U14617 ( .DIN(n4752), .Q(n4739) );
  xor2s1 U14618 ( .DIN1(n5021), .DIN2(n5421), .Q(n4752) );
  hi1s1 U14619 ( .DIN(n13009), .Q(n5421) );
  or3s1 U14620 ( .DIN1(n14433), .DIN2(n14434), .DIN3(n14435), .Q(n13009) );
  nnd4s1 U14621 ( .DIN1(n13407), .DIN2(n14436), .DIN3(n14437), .DIN4(n14438), 
        .Q(n14435) );
  and4s1 U14622 ( .DIN1(n14439), .DIN2(n14184), .DIN3(n14440), .DIN4(n14441), 
        .Q(n14438) );
  nnd2s1 U14623 ( .DIN1(n14214), .DIN2(n13706), .Q(n14441) );
  nnd2s1 U14624 ( .DIN1(n13903), .DIN2(n13412), .Q(n14440) );
  nnd2s1 U14625 ( .DIN1(n13902), .DIN2(n13413), .Q(n14184) );
  nor4s1 U14626 ( .DIN1(n14442), .DIN2(n14443), .DIN3(n14444), .DIN4(n14445), 
        .Q(n13407) );
  nnd4s1 U14627 ( .DIN1(n14446), .DIN2(n14447), .DIN3(n13699), .DIN4(n14448), 
        .Q(n14445) );
  nor2s1 U14628 ( .DIN1(n14449), .DIN2(n14450), .Q(n14448) );
  nor2s1 U14629 ( .DIN1(n13721), .DIN2(n13399), .Q(n14450) );
  nor2s1 U14630 ( .DIN1(n14451), .DIN2(n13720), .Q(n14449) );
  nnd2s1 U14631 ( .DIN1(n13903), .DIN2(n13908), .Q(n13699) );
  nnd2s1 U14632 ( .DIN1(n13387), .DIN2(n14165), .Q(n14447) );
  nnd3s1 U14633 ( .DIN1(n14452), .DIN2(n14453), .DIN3(n14454), .Q(n14444) );
  nnd2s1 U14634 ( .DIN1(n13415), .DIN2(n14191), .Q(n14454) );
  nnd2s1 U14635 ( .DIN1(n13396), .DIN2(n13914), .Q(n14191) );
  nnd2s1 U14636 ( .DIN1(n14214), .DIN2(n14455), .Q(n14453) );
  nnd3s1 U14637 ( .DIN1(n14154), .DIN2(n13400), .DIN3(n14456), .Q(n14455) );
  nnd2s1 U14638 ( .DIN1(n13902), .DIN2(n14457), .Q(n14452) );
  nnd3s1 U14639 ( .DIN1(n14451), .DIN2(n14201), .DIN3(n14458), .Q(n14457) );
  nor2s1 U14640 ( .DIN1(n14459), .DIN2(n14201), .Q(n14443) );
  nor2s1 U14641 ( .DIN1(n14460), .DIN2(n14461), .Q(n14442) );
  nnd4s1 U14642 ( .DIN1(n14462), .DIN2(n14463), .DIN3(n14464), .DIN4(n14465), 
        .Q(n14434) );
  nnd2s1 U14643 ( .DIN1(n13912), .DIN2(n13901), .Q(n14465) );
  nnd2s1 U14644 ( .DIN1(n13898), .DIN2(n13381), .Q(n14464) );
  nnd2s1 U14645 ( .DIN1(n14147), .DIN2(n13386), .Q(n14463) );
  nnd2s1 U14646 ( .DIN1(n13393), .DIN2(n13924), .Q(n14462) );
  nnd4s1 U14647 ( .DIN1(n14466), .DIN2(n14467), .DIN3(n14468), .DIN4(n14469), 
        .Q(n14433) );
  nnd2s1 U14648 ( .DIN1(n13725), .DIN2(n14470), .Q(n14469) );
  nnd2s1 U14649 ( .DIN1(n14471), .DIN2(n14459), .Q(n14470) );
  nnd2s1 U14650 ( .DIN1(n14165), .DIN2(n14171), .Q(n14468) );
  nnd2s1 U14651 ( .DIN1(n14151), .DIN2(n14472), .Q(n14467) );
  nnd2s1 U14652 ( .DIN1(n14473), .DIN2(n13931), .Q(n14472) );
  nnd2s1 U14653 ( .DIN1(n13932), .DIN2(n13384), .Q(n14466) );
  nor3s1 U14654 ( .DIN1(n14474), .DIN2(n14475), .DIN3(n14476), .Q(n5021) );
  nnd4s1 U14655 ( .DIN1(n14477), .DIN2(n13450), .DIN3(n14478), .DIN4(n14479), 
        .Q(n14476) );
  and4s1 U14656 ( .DIN1(n14480), .DIN2(n13987), .DIN3(n14481), .DIN4(n14482), 
        .Q(n14479) );
  nnd2s1 U14657 ( .DIN1(n13660), .DIN2(n14017), .Q(n14482) );
  nnd2s1 U14658 ( .DIN1(n13455), .DIN2(n13778), .Q(n14481) );
  nnd2s1 U14659 ( .DIN1(n13456), .DIN2(n13777), .Q(n13987) );
  nor4s1 U14660 ( .DIN1(n14483), .DIN2(n14484), .DIN3(n14485), .DIN4(n14486), 
        .Q(n13450) );
  nnd4s1 U14661 ( .DIN1(n14267), .DIN2(n14487), .DIN3(n13652), .DIN4(n14488), 
        .Q(n14486) );
  nor2s1 U14662 ( .DIN1(n14489), .DIN2(n14490), .Q(n14488) );
  nor2s1 U14663 ( .DIN1(n13674), .DIN2(n13442), .Q(n14490) );
  nor2s1 U14664 ( .DIN1(n14251), .DIN2(n13673), .Q(n14489) );
  nnd2s1 U14665 ( .DIN1(n13778), .DIN2(n13783), .Q(n13652) );
  nnd2s1 U14666 ( .DIN1(n13431), .DIN2(n13968), .Q(n14487) );
  nnd2s1 U14667 ( .DIN1(n13969), .DIN2(n13678), .Q(n14267) );
  nnd3s1 U14668 ( .DIN1(n14491), .DIN2(n14492), .DIN3(n14493), .Q(n14485) );
  nnd2s1 U14669 ( .DIN1(n13458), .DIN2(n13994), .Q(n14493) );
  nnd2s1 U14670 ( .DIN1(n13439), .DIN2(n13789), .Q(n13994) );
  nnd2s1 U14671 ( .DIN1(n14017), .DIN2(n14494), .Q(n14492) );
  nnd3s1 U14672 ( .DIN1(n13957), .DIN2(n14323), .DIN3(n13443), .Q(n14494) );
  nnd2s1 U14673 ( .DIN1(n13777), .DIN2(n14495), .Q(n14491) );
  nnd3s1 U14674 ( .DIN1(n14003), .DIN2(n14237), .DIN3(n14251), .Q(n14495) );
  nor2s1 U14675 ( .DIN1(n14003), .DIN2(n14277), .Q(n14484) );
  nor2s1 U14676 ( .DIN1(n14291), .DIN2(n14257), .Q(n14483) );
  nnd4s1 U14677 ( .DIN1(n14496), .DIN2(n14497), .DIN3(n14498), .DIN4(n14499), 
        .Q(n14475) );
  nnd2s1 U14678 ( .DIN1(n13787), .DIN2(n13776), .Q(n14499) );
  nnd2s1 U14679 ( .DIN1(n13773), .DIN2(n13424), .Q(n14498) );
  nnd2s1 U14680 ( .DIN1(n13950), .DIN2(n13429), .Q(n14497) );
  nnd2s1 U14681 ( .DIN1(n13436), .DIN2(n13799), .Q(n14496) );
  nnd4s1 U14682 ( .DIN1(n14500), .DIN2(n14501), .DIN3(n14502), .DIN4(n14503), 
        .Q(n14474) );
  nnd2s1 U14683 ( .DIN1(n13678), .DIN2(n14504), .Q(n14503) );
  nnd2s1 U14684 ( .DIN1(n14234), .DIN2(n14277), .Q(n14504) );
  nnd2s1 U14685 ( .DIN1(n13968), .DIN2(n13974), .Q(n14502) );
  nnd2s1 U14686 ( .DIN1(n13954), .DIN2(n14505), .Q(n14501) );
  nnd2s1 U14687 ( .DIN1(n14506), .DIN2(n13806), .Q(n14505) );
  nnd2s1 U14688 ( .DIN1(n13807), .DIN2(n13427), .Q(n14500) );
  hi1s1 U14689 ( .DIN(n12943), .Q(n12950) );
  xor2s1 U14690 ( .DIN1(n5064), .DIN2(n14507), .Q(n12943) );
  hi1s1 U14691 ( .DIN(n5417), .Q(n14507) );
  or3s1 U14692 ( .DIN1(n14508), .DIN2(n14509), .DIN3(n14510), .Q(n5417) );
  nnd4s1 U14693 ( .DIN1(n14511), .DIN2(n14512), .DIN3(n13701), .DIN4(n14513), 
        .Q(n14510) );
  and3s1 U14694 ( .DIN1(n13884), .DIN2(n14179), .DIN3(n14156), .Q(n14513) );
  nor4s1 U14695 ( .DIN1(n14514), .DIN2(n14515), .DIN3(n14516), .DIN4(n14517), 
        .Q(n14156) );
  nnd4s1 U14696 ( .DIN1(n14518), .DIN2(n14519), .DIN3(n14520), .DIN4(n14521), 
        .Q(n14517) );
  nor2s1 U14697 ( .DIN1(n14522), .DIN2(n14523), .Q(n14521) );
  nor2s1 U14698 ( .DIN1(n14458), .DIN2(n13395), .Q(n14523) );
  nor2s1 U14699 ( .DIN1(n13727), .DIN2(n14154), .Q(n14522) );
  nnd2s1 U14700 ( .DIN1(n14147), .DIN2(n13908), .Q(n14520) );
  nnd2s1 U14701 ( .DIN1(n13413), .DIN2(n13386), .Q(n14519) );
  nnd2s1 U14702 ( .DIN1(n13385), .DIN2(n13707), .Q(n14518) );
  nnd3s1 U14703 ( .DIN1(n14524), .DIN2(n14525), .DIN3(n14526), .Q(n14516) );
  nnd2s1 U14704 ( .DIN1(n13383), .DIN2(n13935), .Q(n14526) );
  nnd2s1 U14705 ( .DIN1(n13403), .DIN2(n14527), .Q(n14525) );
  nnd3s1 U14706 ( .DIN1(n13396), .DIN2(n13714), .DIN3(n13724), .Q(n14527) );
  nnd2s1 U14707 ( .DIN1(n14214), .DIN2(n14528), .Q(n14524) );
  nnd3s1 U14708 ( .DIN1(n14201), .DIN2(n13910), .DIN3(n14458), .Q(n14528) );
  nor2s1 U14709 ( .DIN1(n13711), .DIN2(n14529), .Q(n14515) );
  nor2s1 U14710 ( .DIN1(n14530), .DIN2(n14471), .Q(n14514) );
  nor4s1 U14711 ( .DIN1(n14531), .DIN2(n14532), .DIN3(n14533), .DIN4(n14534), 
        .Q(n14179) );
  nnd4s1 U14712 ( .DIN1(n14535), .DIN2(n14536), .DIN3(n14537), .DIN4(n14538), 
        .Q(n14534) );
  nor2s1 U14713 ( .DIN1(n14539), .DIN2(n14540), .Q(n14538) );
  nor2s1 U14714 ( .DIN1(n14201), .DIN2(n13721), .Q(n14540) );
  nor2s1 U14715 ( .DIN1(n13396), .DIN2(n14451), .Q(n14539) );
  nnd2s1 U14716 ( .DIN1(n13898), .DIN2(n13924), .Q(n14536) );
  nnd3s1 U14717 ( .DIN1(n14541), .DIN2(n14542), .DIN3(n14543), .Q(n14533) );
  nnd2s1 U14718 ( .DIN1(n13415), .DIN2(n14544), .Q(n14543) );
  nnd2s1 U14719 ( .DIN1(n14545), .DIN2(n13396), .Q(n14544) );
  nnd2s1 U14720 ( .DIN1(n13707), .DIN2(n13723), .Q(n14542) );
  nnd2s1 U14721 ( .DIN1(n13912), .DIN2(n13934), .Q(n14541) );
  nnd2s1 U14722 ( .DIN1(n14461), .DIN2(n13720), .Q(n13934) );
  nor2s1 U14723 ( .DIN1(n14546), .DIN2(n13930), .Q(n14532) );
  nor2s1 U14724 ( .DIN1(n13924), .DIN2(n14165), .Q(n14546) );
  nor2s1 U14725 ( .DIN1(n14547), .DIN2(n13395), .Q(n14531) );
  nor2s1 U14726 ( .DIN1(n13403), .DIN2(n13383), .Q(n14547) );
  nor4s1 U14727 ( .DIN1(n14548), .DIN2(n14549), .DIN3(n14550), .DIN4(n14551), 
        .Q(n13884) );
  nnd4s1 U14728 ( .DIN1(n14552), .DIN2(n14553), .DIN3(n14554), .DIN4(n14446), 
        .Q(n14551) );
  nnd2s1 U14729 ( .DIN1(n13725), .DIN2(n14166), .Q(n14446) );
  nor2s1 U14730 ( .DIN1(n14555), .DIN2(n14556), .Q(n14554) );
  nor2s1 U14731 ( .DIN1(n13727), .DIN2(n13911), .Q(n14556) );
  nor2s1 U14732 ( .DIN1(n13714), .DIN2(n14200), .Q(n14555) );
  nnd2s1 U14733 ( .DIN1(n14151), .DIN2(n13385), .Q(n14553) );
  nnd2s1 U14734 ( .DIN1(n13397), .DIN2(n13413), .Q(n14552) );
  nnd3s1 U14735 ( .DIN1(n14557), .DIN2(n14558), .DIN3(n14559), .Q(n14550) );
  nnd2s1 U14736 ( .DIN1(n13706), .DIN2(n14560), .Q(n14559) );
  nnd2s1 U14737 ( .DIN1(n13415), .DIN2(n14561), .Q(n14558) );
  nnd2s1 U14738 ( .DIN1(n13403), .DIN2(n14562), .Q(n14557) );
  nnd3s1 U14739 ( .DIN1(n14471), .DIN2(n14150), .DIN3(n14563), .Q(n14562) );
  nor2s1 U14740 ( .DIN1(n14459), .DIN2(n13910), .Q(n14549) );
  nor2s1 U14741 ( .DIN1(n14564), .DIN2(n13931), .Q(n14548) );
  and4s1 U14742 ( .DIN1(n14180), .DIN2(n14213), .DIN3(n14565), .DIN4(n14566), 
        .Q(n13701) );
  and4s1 U14743 ( .DIN1(n14567), .DIN2(n14568), .DIN3(n14569), .DIN4(n14570), 
        .Q(n14566) );
  and3s1 U14744 ( .DIN1(n14571), .DIN2(n14572), .DIN3(n14573), .Q(n14570) );
  nnd2s1 U14745 ( .DIN1(n13383), .DIN2(n14574), .Q(n14573) );
  nnd2s1 U14746 ( .DIN1(n13721), .DIN2(n13396), .Q(n14574) );
  nnd2s1 U14747 ( .DIN1(n13898), .DIN2(n14575), .Q(n14572) );
  nnd2s1 U14748 ( .DIN1(n13724), .DIN2(n14459), .Q(n14575) );
  nnd2s1 U14749 ( .DIN1(n13706), .DIN2(n14576), .Q(n14571) );
  nnd2s1 U14750 ( .DIN1(n13720), .DIN2(n14459), .Q(n14576) );
  or2s1 U14751 ( .DIN1(n13918), .DIN2(n14460), .Q(n14569) );
  nnd2s1 U14752 ( .DIN1(n13413), .DIN2(n14577), .Q(n14568) );
  or2s1 U14753 ( .DIN1(n13935), .DIN2(n14214), .Q(n14577) );
  nnd2s1 U14754 ( .DIN1(n13727), .DIN2(n13711), .Q(n13935) );
  nnd2s1 U14755 ( .DIN1(n13414), .DIN2(n14578), .Q(n14567) );
  nnd3s1 U14756 ( .DIN1(n14458), .DIN2(n14200), .DIN3(n14579), .Q(n14578) );
  and3s1 U14757 ( .DIN1(n14580), .DIN2(n14581), .DIN3(n13886), .Q(n14565) );
  nor4s1 U14758 ( .DIN1(n14582), .DIN2(n14583), .DIN3(n14584), .DIN4(n14585), 
        .Q(n13886) );
  nnd4s1 U14759 ( .DIN1(n14586), .DIN2(n14587), .DIN3(n14588), .DIN4(n14589), 
        .Q(n14585) );
  nnd2s1 U14760 ( .DIN1(n14214), .DIN2(n13383), .Q(n14589) );
  nnd2s1 U14761 ( .DIN1(n14151), .DIN2(n13387), .Q(n14588) );
  nnd2s1 U14762 ( .DIN1(n13902), .DIN2(n13725), .Q(n14587) );
  nnd2s1 U14763 ( .DIN1(n13932), .DIN2(n14165), .Q(n14586) );
  nnd3s1 U14764 ( .DIN1(n14590), .DIN2(n14591), .DIN3(n14592), .Q(n14584) );
  nnd2s1 U14765 ( .DIN1(n13393), .DIN2(n14593), .Q(n14592) );
  nnd3s1 U14766 ( .DIN1(n14461), .DIN2(n13727), .DIN3(n13918), .Q(n14593) );
  nnd2s1 U14767 ( .DIN1(n13385), .DIN2(n14594), .Q(n14591) );
  nnd2s1 U14768 ( .DIN1(n14471), .DIN2(n13728), .Q(n14594) );
  nnd2s1 U14769 ( .DIN1(n13890), .DIN2(n14595), .Q(n14590) );
  nnd2s1 U14770 ( .DIN1(n14545), .DIN2(n13918), .Q(n14595) );
  nor2s1 U14771 ( .DIN1(n13414), .DIN2(n14596), .Q(n14545) );
  nor2s1 U14772 ( .DIN1(n13728), .DIN2(n14153), .Q(n14583) );
  nor2s1 U14773 ( .DIN1(n13900), .DIN2(n14154), .Q(n14582) );
  hi1s1 U14774 ( .DIN(n13384), .Q(n13900) );
  nnd2s1 U14775 ( .DIN1(n13412), .DIN2(n13725), .Q(n14581) );
  nnd2s1 U14776 ( .DIN1(n13385), .DIN2(n14165), .Q(n14580) );
  nor4s1 U14777 ( .DIN1(n14597), .DIN2(n14598), .DIN3(n14599), .DIN4(n14600), 
        .Q(n14213) );
  nnd4s1 U14778 ( .DIN1(n14601), .DIN2(n14602), .DIN3(n14603), .DIN4(n14604), 
        .Q(n14600) );
  nnd2s1 U14779 ( .DIN1(n13414), .DIN2(n14192), .Q(n14604) );
  nor2s1 U14780 ( .DIN1(n14605), .DIN2(n14606), .Q(n14603) );
  nor2s1 U14781 ( .DIN1(n14607), .DIN2(n14456), .Q(n14606) );
  nor2s1 U14782 ( .DIN1(n13386), .DIN2(n14214), .Q(n14607) );
  nor2s1 U14783 ( .DIN1(n14608), .DIN2(n13930), .Q(n14605) );
  nor2s1 U14784 ( .DIN1(n13412), .DIN2(n14609), .Q(n14608) );
  nnd2s1 U14785 ( .DIN1(n14151), .DIN2(n14610), .Q(n14602) );
  nnd3s1 U14786 ( .DIN1(n14200), .DIN2(n13399), .DIN3(n13911), .Q(n14610) );
  nnd2s1 U14787 ( .DIN1(n13912), .DIN2(n13707), .Q(n14601) );
  nnd3s1 U14788 ( .DIN1(n14611), .DIN2(n14612), .DIN3(n14613), .Q(n14599) );
  nnd2s1 U14789 ( .DIN1(n14147), .DIN2(n14214), .Q(n14612) );
  nnd2s1 U14790 ( .DIN1(n14596), .DIN2(n13383), .Q(n14611) );
  nor2s1 U14791 ( .DIN1(n14153), .DIN2(n14471), .Q(n14598) );
  nor2s1 U14792 ( .DIN1(n13721), .DIN2(n14529), .Q(n14597) );
  nor2s1 U14793 ( .DIN1(n14614), .DIN2(n14615), .Q(n14180) );
  nnd4s1 U14794 ( .DIN1(n14616), .DIN2(n14617), .DIN3(n14618), .DIN4(n14619), 
        .Q(n14615) );
  nnd2s1 U14795 ( .DIN1(n14165), .DIN2(n14620), .Q(n14619) );
  nnd3s1 U14796 ( .DIN1(n14458), .DIN2(n14154), .DIN3(n13911), .Q(n14620) );
  nnd2s1 U14797 ( .DIN1(n14147), .DIN2(n13381), .Q(n14618) );
  nnd4s1 U14798 ( .DIN1(n14621), .DIN2(n14622), .DIN3(n14623), .DIN4(n14624), 
        .Q(n14614) );
  nnd2s1 U14799 ( .DIN1(n13386), .DIN2(n14625), .Q(n14624) );
  nnd2s1 U14800 ( .DIN1(n13911), .DIN2(n14146), .Q(n14625) );
  nnd2s1 U14801 ( .DIN1(n13388), .DIN2(n14626), .Q(n14623) );
  nnd2s1 U14802 ( .DIN1(n13712), .DIN2(n13399), .Q(n14626) );
  nnd2s1 U14803 ( .DIN1(n13932), .DIN2(n14627), .Q(n14622) );
  nnd2s1 U14804 ( .DIN1(n14628), .DIN2(n13727), .Q(n14627) );
  nnd2s1 U14805 ( .DIN1(n13903), .DIN2(n14629), .Q(n14621) );
  nnd2s1 U14806 ( .DIN1(n13725), .DIN2(n13908), .Q(n14511) );
  nnd3s1 U14807 ( .DIN1(n14630), .DIN2(n14631), .DIN3(n14632), .Q(n14509) );
  nnd2s1 U14808 ( .DIN1(n14596), .DIN2(n13932), .Q(n14632) );
  nnd2s1 U14809 ( .DIN1(n14166), .DIN2(n13382), .Q(n14631) );
  nnd2s1 U14810 ( .DIN1(n13898), .DIN2(n13397), .Q(n14630) );
  nnd4s1 U14811 ( .DIN1(n14633), .DIN2(n14634), .DIN3(n14635), .DIN4(n14636), 
        .Q(n14508) );
  nnd2s1 U14812 ( .DIN1(n13924), .DIN2(n14637), .Q(n14636) );
  nnd2s1 U14813 ( .DIN1(n14200), .DIN2(n13916), .Q(n14637) );
  nnd2s1 U14814 ( .DIN1(n13902), .DIN2(n14638), .Q(n14635) );
  nnd2s1 U14815 ( .DIN1(n13402), .DIN2(n14201), .Q(n14638) );
  nor2s1 U14816 ( .DIN1(n13415), .DIN2(n13898), .Q(n13402) );
  nnd2s1 U14817 ( .DIN1(n13890), .DIN2(n14639), .Q(n14634) );
  nnd2s1 U14818 ( .DIN1(n14564), .DIN2(n13401), .Q(n14639) );
  nor2s1 U14819 ( .DIN1(n13902), .DIN2(n13381), .Q(n14564) );
  nnd2s1 U14820 ( .DIN1(n14151), .DIN2(n14192), .Q(n14633) );
  or3s1 U14821 ( .DIN1(n14640), .DIN2(n14641), .DIN3(n14642), .Q(n5064) );
  nnd4s1 U14822 ( .DIN1(n14643), .DIN2(n13339), .DIN3(n13734), .DIN4(n14644), 
        .Q(n14642) );
  and3s1 U14823 ( .DIN1(n13845), .DIN2(n14103), .DIN3(n14082), .Q(n14644) );
  nor4s1 U14824 ( .DIN1(n14645), .DIN2(n14646), .DIN3(n14647), .DIN4(n14648), 
        .Q(n14082) );
  nnd4s1 U14825 ( .DIN1(n14649), .DIN2(n14650), .DIN3(n14651), .DIN4(n14652), 
        .Q(n14648) );
  nor2s1 U14826 ( .DIN1(n14653), .DIN2(n14654), .Q(n14652) );
  nor2s1 U14827 ( .DIN1(n13505), .DIN2(n13286), .Q(n14654) );
  nor2s1 U14828 ( .DIN1(n13520), .DIN2(n13365), .Q(n14653) );
  nnd2s1 U14829 ( .DIN1(n13539), .DIN2(n13331), .Q(n14650) );
  nnd2s1 U14830 ( .DIN1(n13306), .DIN2(n13293), .Q(n14649) );
  nnd3s1 U14831 ( .DIN1(n14655), .DIN2(n14656), .DIN3(n14657), .Q(n14647) );
  nnd2s1 U14832 ( .DIN1(n13369), .DIN2(n13872), .Q(n14657) );
  nnd2s1 U14833 ( .DIN1(n13505), .DIN2(n13520), .Q(n13872) );
  nnd2s1 U14834 ( .DIN1(n13333), .DIN2(n14658), .Q(n14656) );
  nnd3s1 U14835 ( .DIN1(n13541), .DIN2(n13863), .DIN3(n13285), .Q(n14658) );
  nnd2s1 U14836 ( .DIN1(n13292), .DIN2(n14659), .Q(n14655) );
  nnd3s1 U14837 ( .DIN1(n13749), .DIN2(n13742), .DIN3(n13324), .Q(n14659) );
  nor2s1 U14838 ( .DIN1(n13324), .DIN2(n13558), .Q(n14646) );
  and2s1 U14839 ( .DIN1(n13334), .DIN2(n13290), .Q(n14645) );
  nor4s1 U14840 ( .DIN1(n14660), .DIN2(n14661), .DIN3(n14662), .DIN4(n14663), 
        .Q(n14103) );
  nnd4s1 U14841 ( .DIN1(n14664), .DIN2(n14665), .DIN3(n14666), .DIN4(n14667), 
        .Q(n14663) );
  nor2s1 U14842 ( .DIN1(n14668), .DIN2(n14669), .Q(n14666) );
  nor2s1 U14843 ( .DIN1(n13541), .DIN2(n13282), .Q(n14669) );
  nor2s1 U14844 ( .DIN1(n13324), .DIN2(n13495), .Q(n14668) );
  nnd2s1 U14845 ( .DIN1(n13283), .DIN2(n13371), .Q(n14665) );
  nnd2s1 U14846 ( .DIN1(n13548), .DIN2(n13353), .Q(n14664) );
  nnd3s1 U14847 ( .DIN1(n14670), .DIN2(n14671), .DIN3(n14672), .Q(n14662) );
  nnd2s1 U14848 ( .DIN1(n13304), .DIN2(n13877), .Q(n14672) );
  nnd2s1 U14849 ( .DIN1(n13498), .DIN2(n13557), .Q(n13877) );
  nnd2s1 U14850 ( .DIN1(n13490), .DIN2(n14673), .Q(n14671) );
  nnd2s1 U14851 ( .DIN1(n14078), .DIN2(n13863), .Q(n14673) );
  nnd2s1 U14852 ( .DIN1(n13342), .DIN2(n14674), .Q(n14670) );
  nnd2s1 U14853 ( .DIN1(n14675), .DIN2(n13324), .Q(n14674) );
  nor2s1 U14854 ( .DIN1(n14676), .DIN2(n13496), .Q(n14661) );
  nor2s1 U14855 ( .DIN1(n13353), .DIN2(n13303), .Q(n14676) );
  nor2s1 U14856 ( .DIN1(n14677), .DIN2(n13281), .Q(n14660) );
  nor2s1 U14857 ( .DIN1(n13292), .DIN2(n13369), .Q(n14677) );
  nor4s1 U14858 ( .DIN1(n14678), .DIN2(n14679), .DIN3(n14680), .DIN4(n14681), 
        .Q(n13845) );
  nnd4s1 U14859 ( .DIN1(n14682), .DIN2(n14683), .DIN3(n14684), .DIN4(n14685), 
        .Q(n14681) );
  nor2s1 U14860 ( .DIN1(n14686), .DIN2(n14687), .Q(n14684) );
  nor2s1 U14861 ( .DIN1(n13278), .DIN2(n13557), .Q(n14687) );
  nor2s1 U14862 ( .DIN1(n13555), .DIN2(n13863), .Q(n14686) );
  nnd2s1 U14863 ( .DIN1(n13290), .DIN2(n13306), .Q(n14683) );
  nnd2s1 U14864 ( .DIN1(n13553), .DIN2(n13302), .Q(n14682) );
  nnd3s1 U14865 ( .DIN1(n14688), .DIN2(n14689), .DIN3(n14690), .Q(n14680) );
  nnd2s1 U14866 ( .DIN1(n13371), .DIN2(n13370), .Q(n14690) );
  nnd2s1 U14867 ( .DIN1(n13742), .DIN2(n13282), .Q(n13370) );
  nnd2s1 U14868 ( .DIN1(n13342), .DIN2(n14691), .Q(n14689) );
  nnd2s1 U14869 ( .DIN1(n13292), .DIN2(n14692), .Q(n14688) );
  nnd3s1 U14870 ( .DIN1(n14080), .DIN2(n13282), .DIN3(n14693), .Q(n14692) );
  nor2s1 U14871 ( .DIN1(n13558), .DIN2(n13742), .Q(n14679) );
  nor2s1 U14872 ( .DIN1(n13751), .DIN2(n14694), .Q(n14678) );
  and4s1 U14873 ( .DIN1(n14104), .DIN2(n13847), .DIN3(n14695), .DIN4(n14696), 
        .Q(n13734) );
  and4s1 U14874 ( .DIN1(n14697), .DIN2(n14698), .DIN3(n14699), .DIN4(n14700), 
        .Q(n14696) );
  and3s1 U14875 ( .DIN1(n14701), .DIN2(n14702), .DIN3(n14703), .Q(n14700) );
  nnd2s1 U14876 ( .DIN1(n13369), .DIN2(n14704), .Q(n14703) );
  nnd2s1 U14877 ( .DIN1(n13499), .DIN2(n13324), .Q(n14704) );
  nnd2s1 U14878 ( .DIN1(n13371), .DIN2(n14705), .Q(n14702) );
  nnd2s1 U14879 ( .DIN1(n13557), .DIN2(n13555), .Q(n14705) );
  nnd2s1 U14880 ( .DIN1(n13548), .DIN2(n14706), .Q(n14701) );
  nnd2s1 U14881 ( .DIN1(n13749), .DIN2(n13555), .Q(n14706) );
  or2s1 U14882 ( .DIN1(n13519), .DIN2(n13542), .Q(n14699) );
  nnd2s1 U14883 ( .DIN1(n13306), .DIN2(n14707), .Q(n14698) );
  nnd2s1 U14884 ( .DIN1(n13505), .DIN2(n14080), .Q(n14707) );
  nnd2s1 U14885 ( .DIN1(n13305), .DIN2(n14708), .Q(n14697) );
  nnd3s1 U14886 ( .DIN1(n13558), .DIN2(n13541), .DIN3(n14081), .Q(n14708) );
  and3s1 U14887 ( .DIN1(n14709), .DIN2(n14710), .DIN3(n14133), .Q(n14695) );
  nor4s1 U14888 ( .DIN1(n14711), .DIN2(n14712), .DIN3(n14713), .DIN4(n14714), 
        .Q(n14133) );
  nnd4s1 U14889 ( .DIN1(n14715), .DIN2(n14716), .DIN3(n14717), .DIN4(n14718), 
        .Q(n14714) );
  nnd2s1 U14890 ( .DIN1(n13301), .DIN2(n14719), .Q(n14718) );
  nnd2s1 U14891 ( .DIN1(n13752), .DIN2(n13326), .Q(n14719) );
  nor2s1 U14892 ( .DIN1(n14720), .DIN2(n14721), .Q(n14717) );
  nor2s1 U14893 ( .DIN1(n14722), .DIN2(n13498), .Q(n14721) );
  nor2s1 U14894 ( .DIN1(n13292), .DIN2(n13553), .Q(n14722) );
  nor2s1 U14895 ( .DIN1(n14723), .DIN2(n13278), .Q(n14720) );
  nor2s1 U14896 ( .DIN1(n13333), .DIN2(n13293), .Q(n14723) );
  nnd2s1 U14897 ( .DIN1(n13275), .DIN2(n14724), .Q(n14716) );
  nnd3s1 U14898 ( .DIN1(n13368), .DIN2(n13502), .DIN3(n13558), .Q(n14724) );
  nnd2s1 U14899 ( .DIN1(n13333), .DIN2(n13359), .Q(n14715) );
  nnd3s1 U14900 ( .DIN1(n14725), .DIN2(n14726), .DIN3(n14727), .Q(n14713) );
  nnd2s1 U14901 ( .DIN1(n13290), .DIN2(n13279), .Q(n14727) );
  nnd2s1 U14902 ( .DIN1(n13490), .DIN2(n13304), .Q(n14725) );
  nor2s1 U14903 ( .DIN1(n13749), .DIN2(n13277), .Q(n14712) );
  nor2s1 U14904 ( .DIN1(n13499), .DIN2(n13365), .Q(n14711) );
  nnd2s1 U14905 ( .DIN1(n13303), .DIN2(n13341), .Q(n14710) );
  nnd2s1 U14906 ( .DIN1(n13553), .DIN2(n13480), .Q(n14709) );
  nor4s1 U14907 ( .DIN1(n14728), .DIN2(n14729), .DIN3(n14730), .DIN4(n14731), 
        .Q(n13847) );
  nnd4s1 U14908 ( .DIN1(n14732), .DIN2(n14733), .DIN3(n14734), .DIN4(n14735), 
        .Q(n14731) );
  nor2s1 U14909 ( .DIN1(n14736), .DIN2(n14737), .Q(n14735) );
  nor2s1 U14910 ( .DIN1(n13277), .DIN2(n14080), .Q(n14737) );
  nor2s1 U14911 ( .DIN1(n13559), .DIN2(n13286), .Q(n14736) );
  nnd2s1 U14912 ( .DIN1(n13330), .DIN2(n14738), .Q(n14734) );
  nnd2s1 U14913 ( .DIN1(n14078), .DIN2(n13278), .Q(n14738) );
  nnd2s1 U14914 ( .DIN1(n13291), .DIN2(n14739), .Q(n14733) );
  nnd2s1 U14915 ( .DIN1(n14675), .DIN2(n13519), .Q(n14739) );
  nor2s1 U14916 ( .DIN1(n13305), .DIN2(n13358), .Q(n14675) );
  nnd2s1 U14917 ( .DIN1(n13288), .DIN2(n14740), .Q(n14732) );
  nnd2s1 U14918 ( .DIN1(n14129), .DIN2(n13519), .Q(n14740) );
  nor2s1 U14919 ( .DIN1(n13305), .DIN2(n13353), .Q(n14129) );
  nnd3s1 U14920 ( .DIN1(n14741), .DIN2(n14742), .DIN3(n14743), .Q(n14730) );
  nnd2s1 U14921 ( .DIN1(n13306), .DIN2(n13500), .Q(n14743) );
  nnd2s1 U14922 ( .DIN1(n13331), .DIN2(n13275), .Q(n14742) );
  nnd2s1 U14923 ( .DIN1(n13290), .DIN2(n13341), .Q(n14741) );
  nor2s1 U14924 ( .DIN1(n13742), .DIN2(n13495), .Q(n14729) );
  nor2s1 U14925 ( .DIN1(n13365), .DIN2(n13281), .Q(n14728) );
  nor2s1 U14926 ( .DIN1(n14744), .DIN2(n14745), .Q(n14104) );
  nnd4s1 U14927 ( .DIN1(n14746), .DIN2(n14747), .DIN3(n14748), .DIN4(n14749), 
        .Q(n14745) );
  nnd2s1 U14928 ( .DIN1(n13303), .DIN2(n14750), .Q(n14749) );
  nnd3s1 U14929 ( .DIN1(n13541), .DIN2(n13368), .DIN3(n13286), .Q(n14750) );
  nnd2s1 U14930 ( .DIN1(n13283), .DIN2(n13359), .Q(n14748) );
  nnd4s1 U14931 ( .DIN1(n14751), .DIN2(n14752), .DIN3(n14753), .DIN4(n14754), 
        .Q(n14744) );
  nnd2s1 U14932 ( .DIN1(n13293), .DIN2(n13334), .Q(n14754) );
  nnd2s1 U14933 ( .DIN1(n13330), .DIN2(n14755), .Q(n14753) );
  nnd2s1 U14934 ( .DIN1(n13287), .DIN2(n13502), .Q(n14755) );
  nnd2s1 U14935 ( .DIN1(n13489), .DIN2(n14756), .Q(n14752) );
  nnd2s1 U14936 ( .DIN1(n14757), .DIN2(n13505), .Q(n14756) );
  nnd2s1 U14937 ( .DIN1(n13301), .DIN2(n14758), .Q(n14751) );
  nnd2s1 U14938 ( .DIN1(n13519), .DIN2(n13328), .Q(n14758) );
  nnd2s1 U14939 ( .DIN1(n13548), .DIN2(n13290), .Q(n13339) );
  nnd2s1 U14940 ( .DIN1(n13489), .DIN2(n13358), .Q(n14643) );
  nnd3s1 U14941 ( .DIN1(n14759), .DIN2(n14760), .DIN3(n14761), .Q(n14641) );
  nnd2s1 U14942 ( .DIN1(n13302), .DIN2(n13332), .Q(n14760) );
  nnd2s1 U14943 ( .DIN1(n13277), .DIN2(n13558), .Q(n13332) );
  nnd2s1 U14944 ( .DIN1(n13553), .DIN2(n13357), .Q(n14759) );
  nnd4s1 U14945 ( .DIN1(n14762), .DIN2(n14763), .DIN3(n14764), .DIN4(n14765), 
        .Q(n14640) );
  nnd2s1 U14946 ( .DIN1(n13291), .DIN2(n14766), .Q(n14765) );
  nnd2s1 U14947 ( .DIN1(n13751), .DIN2(n13328), .Q(n14766) );
  nor2s1 U14948 ( .DIN1(n13539), .DIN2(n13283), .Q(n13751) );
  nnd2s1 U14949 ( .DIN1(n13353), .DIN2(n14767), .Q(n14764) );
  nnd2s1 U14950 ( .DIN1(n13865), .DIN2(n13558), .Q(n14767) );
  nnd2s1 U14951 ( .DIN1(n13539), .DIN2(n14768), .Q(n14763) );
  nnd2s1 U14952 ( .DIN1(n13329), .DIN2(n13285), .Q(n14768) );
  nor2s1 U14953 ( .DIN1(n13342), .DIN2(n13548), .Q(n13329) );
  nnd2s1 U14954 ( .DIN1(n13275), .DIN2(n13512), .Q(n14762) );
  nnd2s1 U14955 ( .DIN1(n13365), .DIN2(n13865), .Q(n13512) );
  xor2s1 U14956 ( .DIN1(n5040), .DIN2(n14769), .Q(n14430) );
  xor2s1 U14957 ( .DIN1(n1484), .DIN2(n5016), .Q(n14769) );
  or3s1 U14958 ( .DIN1(n14770), .DIN2(n14771), .DIN3(n14772), .Q(n5016) );
  nnd4s1 U14959 ( .DIN1(n14477), .DIN2(n13448), .DIN3(n14773), .DIN4(n14774), 
        .Q(n14772) );
  and3s1 U14960 ( .DIN1(n14775), .DIN2(n14776), .DIN3(n14777), .Q(n14774) );
  nnd2s1 U14961 ( .DIN1(n13954), .DIN2(n13458), .Q(n14776) );
  nnd2s1 U14962 ( .DIN1(n13440), .DIN2(n13660), .Q(n14775) );
  nor4s1 U14963 ( .DIN1(n14778), .DIN2(n14779), .DIN3(n14780), .DIN4(n14781), 
        .Q(n13448) );
  nnd4s1 U14964 ( .DIN1(n14782), .DIN2(n14783), .DIN3(n14784), .DIN4(n14785), 
        .Q(n14781) );
  nor2s1 U14965 ( .DIN1(n14786), .DIN2(n14787), .Q(n14785) );
  nor2s1 U14966 ( .DIN1(n14788), .DIN2(n13786), .Q(n14787) );
  and2s1 U14967 ( .DIN1(n13438), .DIN2(n13976), .Q(n14788) );
  nor2s1 U14968 ( .DIN1(n13969), .DIN2(n13429), .Q(n13976) );
  nor2s1 U14969 ( .DIN1(n14789), .DIN2(n13805), .Q(n14786) );
  nor2s1 U14970 ( .DIN1(n14311), .DIN2(n14017), .Q(n14789) );
  nnd2s1 U14971 ( .DIN1(n13968), .DIN2(n14790), .Q(n14784) );
  nnd2s1 U14972 ( .DIN1(n13785), .DIN2(n14323), .Q(n14790) );
  nnd2s1 U14973 ( .DIN1(n13950), .DIN2(n14791), .Q(n14783) );
  nnd2s1 U14974 ( .DIN1(n13789), .DIN2(n13664), .Q(n14791) );
  nnd2s1 U14975 ( .DIN1(n13783), .DIN2(n14792), .Q(n14782) );
  nnd2s1 U14976 ( .DIN1(n14237), .DIN2(n13791), .Q(n14792) );
  nnd3s1 U14977 ( .DIN1(n14793), .DIN2(n14794), .DIN3(n14795), .Q(n14780) );
  nnd2s1 U14978 ( .DIN1(n13799), .DIN2(n13660), .Q(n14795) );
  nnd2s1 U14979 ( .DIN1(n13766), .DIN2(n13776), .Q(n14794) );
  nnd2s1 U14980 ( .DIN1(n14311), .DIN2(n13458), .Q(n14793) );
  nor2s1 U14981 ( .DIN1(n13793), .DIN2(n13442), .Q(n14779) );
  nor2s1 U14982 ( .DIN1(n13438), .DIN2(n13806), .Q(n14778) );
  nor3s1 U14983 ( .DIN1(n14796), .DIN2(n14797), .DIN3(n14798), .Q(n14477) );
  nnd4s1 U14984 ( .DIN1(n13449), .DIN2(n14799), .DIN3(n14800), .DIN4(n14801), 
        .Q(n14798) );
  and3s1 U14985 ( .DIN1(n14802), .DIN2(n14803), .DIN3(n14332), .Q(n14801) );
  nnd2s1 U14986 ( .DIN1(n13428), .DIN2(n13457), .Q(n14332) );
  nnd2s1 U14987 ( .DIN1(n13440), .DIN2(n13950), .Q(n14803) );
  nnd2s1 U14988 ( .DIN1(n13799), .DIN2(n13766), .Q(n14802) );
  nor4s1 U14989 ( .DIN1(n14804), .DIN2(n14805), .DIN3(n14806), .DIN4(n14807), 
        .Q(n13449) );
  nnd4s1 U14990 ( .DIN1(n14808), .DIN2(n14809), .DIN3(n14329), .DIN4(n14810), 
        .Q(n14807) );
  nnd2s1 U14991 ( .DIN1(n13436), .DIN2(n13429), .Q(n14810) );
  nnd2s1 U14992 ( .DIN1(n13799), .DIN2(n13431), .Q(n14329) );
  nnd2s1 U14993 ( .DIN1(n13783), .DIN2(n13660), .Q(n14809) );
  nnd2s1 U14994 ( .DIN1(n13765), .DIN2(n13457), .Q(n14808) );
  nnd3s1 U14995 ( .DIN1(n14811), .DIN2(n14812), .DIN3(n14813), .Q(n14806) );
  nnd2s1 U14996 ( .DIN1(n13428), .DIN2(n14345), .Q(n14813) );
  nnd2s1 U14997 ( .DIN1(n13793), .DIN2(n13444), .Q(n14345) );
  nnd2s1 U14998 ( .DIN1(n13455), .DIN2(n14814), .Q(n14812) );
  nnd2s1 U14999 ( .DIN1(n14815), .DIN2(n14237), .Q(n14814) );
  nnd2s1 U15000 ( .DIN1(n13778), .DIN2(n14816), .Q(n14811) );
  nnd2s1 U15001 ( .DIN1(n13674), .DIN2(n13680), .Q(n14816) );
  nor2s1 U15002 ( .DIN1(n13677), .DIN2(n13443), .Q(n14805) );
  and2s1 U15003 ( .DIN1(n13678), .DIN2(n14817), .Q(n14804) );
  nnd3s1 U15004 ( .DIN1(n13444), .DIN2(n13681), .DIN3(n13667), .Q(n14817) );
  nnd3s1 U15005 ( .DIN1(n14818), .DIN2(n14819), .DIN3(n14820), .Q(n14797) );
  nnd2s1 U15006 ( .DIN1(n13773), .DIN2(n13777), .Q(n14820) );
  or2s1 U15007 ( .DIN1(n14232), .DIN2(n14344), .Q(n14819) );
  nor2s1 U15008 ( .DIN1(n13455), .DIN2(n14017), .Q(n14344) );
  nnd2s1 U15009 ( .DIN1(n13765), .DIN2(n14325), .Q(n14818) );
  nnd2s1 U15010 ( .DIN1(n13673), .DIN2(n13677), .Q(n14325) );
  nnd4s1 U15011 ( .DIN1(n14821), .DIN2(n14822), .DIN3(n14823), .DIN4(n14824), 
        .Q(n14796) );
  nnd2s1 U15012 ( .DIN1(n13429), .DIN2(n14825), .Q(n14824) );
  nnd2s1 U15013 ( .DIN1(n14294), .DIN2(n14237), .Q(n14825) );
  hi1s1 U15014 ( .DIN(n13798), .Q(n14294) );
  nnd2s1 U15015 ( .DIN1(n13442), .DIN2(n13805), .Q(n13798) );
  nnd2s1 U15016 ( .DIN1(n13424), .DIN2(n14826), .Q(n14823) );
  nnd2s1 U15017 ( .DIN1(n13806), .DIN2(n13791), .Q(n14826) );
  nnd2s1 U15018 ( .DIN1(n13969), .DIN2(n14827), .Q(n14822) );
  nnd2s1 U15019 ( .DIN1(n13436), .DIN2(n14828), .Q(n14821) );
  nnd2s1 U15020 ( .DIN1(n13677), .DIN2(n13444), .Q(n14828) );
  nnd3s1 U15021 ( .DIN1(n14829), .DIN2(n14830), .DIN3(n14831), .Q(n14771) );
  nnd2s1 U15022 ( .DIN1(n13430), .DIN2(n13807), .Q(n14831) );
  or2s1 U15023 ( .DIN1(n13674), .DIN2(n14506), .Q(n14830) );
  nor2s1 U15024 ( .DIN1(n13766), .DIN2(n13678), .Q(n14506) );
  nnd2s1 U15025 ( .DIN1(n13773), .DIN2(n13776), .Q(n14829) );
  nnd4s1 U15026 ( .DIN1(n14832), .DIN2(n14833), .DIN3(n14834), .DIN4(n14835), 
        .Q(n14770) );
  nnd2s1 U15027 ( .DIN1(n14311), .DIN2(n14836), .Q(n14835) );
  nnd2s1 U15028 ( .DIN1(n14291), .DIN2(n13442), .Q(n14836) );
  nor2s1 U15029 ( .DIN1(n13766), .DIN2(n13807), .Q(n14291) );
  nnd2s1 U15030 ( .DIN1(n13799), .DIN2(n14827), .Q(n14834) );
  nnd2s1 U15031 ( .DIN1(n13949), .DIN2(n13806), .Q(n14827) );
  nnd2s1 U15032 ( .DIN1(n13778), .DIN2(n14837), .Q(n14833) );
  nnd2s1 U15033 ( .DIN1(n13977), .DIN2(n13438), .Q(n14837) );
  nor2s1 U15034 ( .DIN1(n13457), .DIN2(n13968), .Q(n13977) );
  nnd2s1 U15035 ( .DIN1(n13436), .DIN2(n14838), .Q(n14832) );
  nnd2s1 U15036 ( .DIN1(n13793), .DIN2(n13789), .Q(n14838) );
  or3s1 U15037 ( .DIN1(n14839), .DIN2(n14840), .DIN3(n14841), .Q(n5040) );
  nnd4s1 U15038 ( .DIN1(n14842), .DIN2(n13229), .DIN3(n13816), .DIN4(n14843), 
        .Q(n14841) );
  and3s1 U15039 ( .DIN1(n14022), .DIN2(n14395), .DIN3(n14374), .Q(n14843) );
  nor4s1 U15040 ( .DIN1(n14844), .DIN2(n14845), .DIN3(n14846), .DIN4(n14847), 
        .Q(n14374) );
  nnd4s1 U15041 ( .DIN1(n14848), .DIN2(n14849), .DIN3(n14850), .DIN4(n14851), 
        .Q(n14847) );
  nor2s1 U15042 ( .DIN1(n14852), .DIN2(n14853), .Q(n14851) );
  nor2s1 U15043 ( .DIN1(n13594), .DIN2(n13166), .Q(n14853) );
  nor2s1 U15044 ( .DIN1(n13609), .DIN2(n13255), .Q(n14852) );
  nnd2s1 U15045 ( .DIN1(n13628), .DIN2(n13221), .Q(n14849) );
  nnd2s1 U15046 ( .DIN1(n13186), .DIN2(n13173), .Q(n14848) );
  nnd3s1 U15047 ( .DIN1(n14854), .DIN2(n14855), .DIN3(n14856), .Q(n14846) );
  nnd2s1 U15048 ( .DIN1(n13259), .DIN2(n14049), .Q(n14856) );
  nnd2s1 U15049 ( .DIN1(n13594), .DIN2(n13609), .Q(n14049) );
  nnd2s1 U15050 ( .DIN1(n13223), .DIN2(n14857), .Q(n14855) );
  nnd3s1 U15051 ( .DIN1(n13630), .DIN2(n14040), .DIN3(n13165), .Q(n14857) );
  nnd2s1 U15052 ( .DIN1(n13172), .DIN2(n14858), .Q(n14854) );
  nnd3s1 U15053 ( .DIN1(n13831), .DIN2(n13824), .DIN3(n13214), .Q(n14858) );
  nor2s1 U15054 ( .DIN1(n13214), .DIN2(n13647), .Q(n14845) );
  and2s1 U15055 ( .DIN1(n13224), .DIN2(n13170), .Q(n14844) );
  nor4s1 U15056 ( .DIN1(n14859), .DIN2(n14860), .DIN3(n14861), .DIN4(n14862), 
        .Q(n14395) );
  nnd4s1 U15057 ( .DIN1(n14863), .DIN2(n14864), .DIN3(n14865), .DIN4(n14866), 
        .Q(n14862) );
  nor2s1 U15058 ( .DIN1(n14867), .DIN2(n14868), .Q(n14865) );
  nor2s1 U15059 ( .DIN1(n13630), .DIN2(n13162), .Q(n14868) );
  nor2s1 U15060 ( .DIN1(n13214), .DIN2(n13584), .Q(n14867) );
  nnd2s1 U15061 ( .DIN1(n13163), .DIN2(n13261), .Q(n14864) );
  nnd2s1 U15062 ( .DIN1(n13637), .DIN2(n13243), .Q(n14863) );
  nnd3s1 U15063 ( .DIN1(n14869), .DIN2(n14870), .DIN3(n14871), .Q(n14861) );
  nnd2s1 U15064 ( .DIN1(n13184), .DIN2(n14054), .Q(n14871) );
  nnd2s1 U15065 ( .DIN1(n13587), .DIN2(n13646), .Q(n14054) );
  nnd2s1 U15066 ( .DIN1(n13579), .DIN2(n14872), .Q(n14870) );
  nnd2s1 U15067 ( .DIN1(n14370), .DIN2(n14040), .Q(n14872) );
  nnd2s1 U15068 ( .DIN1(n13232), .DIN2(n14873), .Q(n14869) );
  nnd2s1 U15069 ( .DIN1(n14874), .DIN2(n13214), .Q(n14873) );
  nor2s1 U15070 ( .DIN1(n14875), .DIN2(n13585), .Q(n14860) );
  nor2s1 U15071 ( .DIN1(n13243), .DIN2(n13183), .Q(n14875) );
  nor2s1 U15072 ( .DIN1(n14876), .DIN2(n13161), .Q(n14859) );
  nor2s1 U15073 ( .DIN1(n13172), .DIN2(n13259), .Q(n14876) );
  nor4s1 U15074 ( .DIN1(n14877), .DIN2(n14878), .DIN3(n14879), .DIN4(n14880), 
        .Q(n14022) );
  nnd4s1 U15075 ( .DIN1(n14881), .DIN2(n14882), .DIN3(n14883), .DIN4(n14884), 
        .Q(n14880) );
  nor2s1 U15076 ( .DIN1(n14885), .DIN2(n14886), .Q(n14883) );
  nor2s1 U15077 ( .DIN1(n13158), .DIN2(n13646), .Q(n14886) );
  nor2s1 U15078 ( .DIN1(n13644), .DIN2(n14040), .Q(n14885) );
  nnd2s1 U15079 ( .DIN1(n13170), .DIN2(n13186), .Q(n14882) );
  nnd2s1 U15080 ( .DIN1(n13642), .DIN2(n13182), .Q(n14881) );
  nnd3s1 U15081 ( .DIN1(n14887), .DIN2(n14888), .DIN3(n14889), .Q(n14879) );
  nnd2s1 U15082 ( .DIN1(n13261), .DIN2(n13260), .Q(n14889) );
  nnd2s1 U15083 ( .DIN1(n13824), .DIN2(n13162), .Q(n13260) );
  nnd2s1 U15084 ( .DIN1(n13232), .DIN2(n14890), .Q(n14888) );
  nnd2s1 U15085 ( .DIN1(n13172), .DIN2(n14891), .Q(n14887) );
  nnd3s1 U15086 ( .DIN1(n14372), .DIN2(n13162), .DIN3(n14892), .Q(n14891) );
  nor2s1 U15087 ( .DIN1(n13647), .DIN2(n13824), .Q(n14878) );
  nor2s1 U15088 ( .DIN1(n13833), .DIN2(n14893), .Q(n14877) );
  and4s1 U15089 ( .DIN1(n14396), .DIN2(n14024), .DIN3(n14894), .DIN4(n14895), 
        .Q(n13816) );
  and4s1 U15090 ( .DIN1(n14896), .DIN2(n14897), .DIN3(n14898), .DIN4(n14899), 
        .Q(n14895) );
  and3s1 U15091 ( .DIN1(n14900), .DIN2(n14901), .DIN3(n14902), .Q(n14899) );
  nnd2s1 U15092 ( .DIN1(n13259), .DIN2(n14903), .Q(n14902) );
  nnd2s1 U15093 ( .DIN1(n13588), .DIN2(n13214), .Q(n14903) );
  nnd2s1 U15094 ( .DIN1(n13261), .DIN2(n14904), .Q(n14901) );
  nnd2s1 U15095 ( .DIN1(n13646), .DIN2(n13644), .Q(n14904) );
  nnd2s1 U15096 ( .DIN1(n13637), .DIN2(n14905), .Q(n14900) );
  nnd2s1 U15097 ( .DIN1(n13831), .DIN2(n13644), .Q(n14905) );
  or2s1 U15098 ( .DIN1(n13608), .DIN2(n13631), .Q(n14898) );
  nnd2s1 U15099 ( .DIN1(n13186), .DIN2(n14906), .Q(n14897) );
  nnd2s1 U15100 ( .DIN1(n13594), .DIN2(n14372), .Q(n14906) );
  nnd2s1 U15101 ( .DIN1(n13185), .DIN2(n14907), .Q(n14896) );
  nnd3s1 U15102 ( .DIN1(n13647), .DIN2(n13630), .DIN3(n14373), .Q(n14907) );
  and3s1 U15103 ( .DIN1(n14908), .DIN2(n14909), .DIN3(n14425), .Q(n14894) );
  nor4s1 U15104 ( .DIN1(n14910), .DIN2(n14911), .DIN3(n14912), .DIN4(n14913), 
        .Q(n14425) );
  nnd4s1 U15105 ( .DIN1(n14914), .DIN2(n14915), .DIN3(n14916), .DIN4(n14917), 
        .Q(n14913) );
  nnd2s1 U15106 ( .DIN1(n13181), .DIN2(n14918), .Q(n14917) );
  nnd2s1 U15107 ( .DIN1(n13834), .DIN2(n13216), .Q(n14918) );
  nor2s1 U15108 ( .DIN1(n14919), .DIN2(n14920), .Q(n14916) );
  nor2s1 U15109 ( .DIN1(n14921), .DIN2(n13587), .Q(n14920) );
  nor2s1 U15110 ( .DIN1(n13172), .DIN2(n13642), .Q(n14921) );
  nor2s1 U15111 ( .DIN1(n14922), .DIN2(n13158), .Q(n14919) );
  nor2s1 U15112 ( .DIN1(n13223), .DIN2(n13173), .Q(n14922) );
  nnd2s1 U15113 ( .DIN1(n13155), .DIN2(n14923), .Q(n14915) );
  nnd3s1 U15114 ( .DIN1(n13258), .DIN2(n13591), .DIN3(n13647), .Q(n14923) );
  nnd2s1 U15115 ( .DIN1(n13223), .DIN2(n13249), .Q(n14914) );
  nnd3s1 U15116 ( .DIN1(n14924), .DIN2(n14925), .DIN3(n14926), .Q(n14912) );
  nnd2s1 U15117 ( .DIN1(n13170), .DIN2(n13159), .Q(n14926) );
  nnd2s1 U15118 ( .DIN1(n13579), .DIN2(n13184), .Q(n14924) );
  nor2s1 U15119 ( .DIN1(n13831), .DIN2(n13157), .Q(n14911) );
  nor2s1 U15120 ( .DIN1(n13588), .DIN2(n13255), .Q(n14910) );
  nnd2s1 U15121 ( .DIN1(n13183), .DIN2(n13231), .Q(n14909) );
  nnd2s1 U15122 ( .DIN1(n13642), .DIN2(n13569), .Q(n14908) );
  nor4s1 U15123 ( .DIN1(n14927), .DIN2(n14928), .DIN3(n14929), .DIN4(n14930), 
        .Q(n14024) );
  nnd4s1 U15124 ( .DIN1(n14931), .DIN2(n14932), .DIN3(n14933), .DIN4(n14934), 
        .Q(n14930) );
  nor2s1 U15125 ( .DIN1(n14935), .DIN2(n14936), .Q(n14934) );
  nor2s1 U15126 ( .DIN1(n13157), .DIN2(n14372), .Q(n14936) );
  nor2s1 U15127 ( .DIN1(n13648), .DIN2(n13166), .Q(n14935) );
  nnd2s1 U15128 ( .DIN1(n13220), .DIN2(n14937), .Q(n14933) );
  nnd2s1 U15129 ( .DIN1(n14370), .DIN2(n13158), .Q(n14937) );
  nnd2s1 U15130 ( .DIN1(n13171), .DIN2(n14938), .Q(n14932) );
  nnd2s1 U15131 ( .DIN1(n14874), .DIN2(n13608), .Q(n14938) );
  nor2s1 U15132 ( .DIN1(n13185), .DIN2(n13248), .Q(n14874) );
  nnd2s1 U15133 ( .DIN1(n13168), .DIN2(n14939), .Q(n14931) );
  nnd2s1 U15134 ( .DIN1(n14421), .DIN2(n13608), .Q(n14939) );
  nor2s1 U15135 ( .DIN1(n13185), .DIN2(n13243), .Q(n14421) );
  nnd3s1 U15136 ( .DIN1(n14940), .DIN2(n14941), .DIN3(n14942), .Q(n14929) );
  nnd2s1 U15137 ( .DIN1(n13186), .DIN2(n13589), .Q(n14942) );
  nnd2s1 U15138 ( .DIN1(n13221), .DIN2(n13155), .Q(n14941) );
  nnd2s1 U15139 ( .DIN1(n13170), .DIN2(n13231), .Q(n14940) );
  nor2s1 U15140 ( .DIN1(n13824), .DIN2(n13584), .Q(n14928) );
  nor2s1 U15141 ( .DIN1(n13255), .DIN2(n13161), .Q(n14927) );
  nor2s1 U15142 ( .DIN1(n14943), .DIN2(n14944), .Q(n14396) );
  nnd4s1 U15143 ( .DIN1(n14945), .DIN2(n14946), .DIN3(n14947), .DIN4(n14948), 
        .Q(n14944) );
  nnd2s1 U15144 ( .DIN1(n13183), .DIN2(n14949), .Q(n14948) );
  nnd3s1 U15145 ( .DIN1(n13630), .DIN2(n13258), .DIN3(n13166), .Q(n14949) );
  nnd2s1 U15146 ( .DIN1(n13163), .DIN2(n13249), .Q(n14947) );
  nnd4s1 U15147 ( .DIN1(n14950), .DIN2(n14951), .DIN3(n14952), .DIN4(n14953), 
        .Q(n14943) );
  nnd2s1 U15148 ( .DIN1(n13173), .DIN2(n13224), .Q(n14953) );
  nnd2s1 U15149 ( .DIN1(n13220), .DIN2(n14954), .Q(n14952) );
  nnd2s1 U15150 ( .DIN1(n13167), .DIN2(n13591), .Q(n14954) );
  nnd2s1 U15151 ( .DIN1(n13578), .DIN2(n14955), .Q(n14951) );
  nnd2s1 U15152 ( .DIN1(n14956), .DIN2(n13594), .Q(n14955) );
  nnd2s1 U15153 ( .DIN1(n13181), .DIN2(n14957), .Q(n14950) );
  nnd2s1 U15154 ( .DIN1(n13608), .DIN2(n13218), .Q(n14957) );
  nnd2s1 U15155 ( .DIN1(n13637), .DIN2(n13170), .Q(n13229) );
  nnd2s1 U15156 ( .DIN1(n13578), .DIN2(n13248), .Q(n14842) );
  nnd3s1 U15157 ( .DIN1(n14958), .DIN2(n14959), .DIN3(n14960), .Q(n14840) );
  nnd2s1 U15158 ( .DIN1(n13182), .DIN2(n13222), .Q(n14959) );
  nnd2s1 U15159 ( .DIN1(n13157), .DIN2(n13647), .Q(n13222) );
  nnd2s1 U15160 ( .DIN1(n13642), .DIN2(n13247), .Q(n14958) );
  nnd4s1 U15161 ( .DIN1(n14961), .DIN2(n14962), .DIN3(n14963), .DIN4(n14964), 
        .Q(n14839) );
  nnd2s1 U15162 ( .DIN1(n13171), .DIN2(n14965), .Q(n14964) );
  nnd2s1 U15163 ( .DIN1(n13833), .DIN2(n13218), .Q(n14965) );
  nor2s1 U15164 ( .DIN1(n13628), .DIN2(n13163), .Q(n13833) );
  nnd2s1 U15165 ( .DIN1(n13243), .DIN2(n14966), .Q(n14963) );
  nnd2s1 U15166 ( .DIN1(n14042), .DIN2(n13647), .Q(n14966) );
  nnd2s1 U15167 ( .DIN1(n13628), .DIN2(n14967), .Q(n14962) );
  nnd2s1 U15168 ( .DIN1(n13219), .DIN2(n13165), .Q(n14967) );
  nor2s1 U15169 ( .DIN1(n13232), .DIN2(n13637), .Q(n13219) );
  nnd2s1 U15170 ( .DIN1(n13155), .DIN2(n13601), .Q(n14961) );
  nnd2s1 U15171 ( .DIN1(n13255), .DIN2(n14042), .Q(n13601) );
  nnd2s1 U15172 ( .DIN1(n14968), .DIN2(n1601), .Q(n14427) );
  xor2s1 U15173 ( .DIN1(w2[3]), .DIN2(text_in_r[35]), .Q(n14968) );
  nnd3s1 U15174 ( .DIN1(n14969), .DIN2(n14970), .DIN3(n14971), .Q(N100) );
  nnd2s1 U15175 ( .DIN1(n1596), .DIN2(n14972), .Q(n14971) );
  xor2s1 U15176 ( .DIN1(w2[2]), .DIN2(text_in_r[34]), .Q(n14972) );
  nnd2s1 U15177 ( .DIN1(n14973), .DIN2(n14974), .Q(n14970) );
  nnd2s1 U15178 ( .DIN1(n14975), .DIN2(n14976), .Q(n14973) );
  nnd2s1 U15179 ( .DIN1(n12964), .DIN2(n5225), .Q(n14976) );
  nnd2s1 U15180 ( .DIN1(n13089), .DIN2(n12966), .Q(n14975) );
  nnd2s1 U15181 ( .DIN1(n14977), .DIN2(n14978), .Q(n14969) );
  nnd2s1 U15182 ( .DIN1(n14979), .DIN2(n14980), .Q(n14978) );
  nnd2s1 U15183 ( .DIN1(n12966), .DIN2(n5225), .Q(n14980) );
  and2s1 U15184 ( .DIN1(n13143), .DIN2(n1543), .Q(n12966) );
  nnd2s1 U15185 ( .DIN1(n13089), .DIN2(n12964), .Q(n14979) );
  nor2s1 U15186 ( .DIN1(n13143), .DIN2(n1595), .Q(n12964) );
  xor2s1 U15187 ( .DIN1(n13070), .DIN2(n5063), .Q(n13143) );
  or3s1 U15188 ( .DIN1(n14981), .DIN2(n14982), .DIN3(n14983), .Q(n5063) );
  nnd4s1 U15189 ( .DIN1(n13336), .DIN2(n13296), .DIN3(n13475), .DIN4(n14984), 
        .Q(n14983) );
  and3s1 U15190 ( .DIN1(n14985), .DIN2(n14986), .DIN3(n13348), .Q(n14984) );
  nor2s1 U15191 ( .DIN1(n14987), .DIN2(n14988), .Q(n13348) );
  nnd4s1 U15192 ( .DIN1(n14667), .DIN2(n14989), .DIN3(n14990), .DIN4(n14991), 
        .Q(n14988) );
  nnd2s1 U15193 ( .DIN1(n13358), .DIN2(n14992), .Q(n14991) );
  nnd2s1 U15194 ( .DIN1(n13277), .DIN2(n13365), .Q(n14992) );
  nnd2s1 U15195 ( .DIN1(n13342), .DIN2(n14993), .Q(n14990) );
  nnd3s1 U15196 ( .DIN1(n13505), .DIN2(n13742), .DIN3(n13281), .Q(n14993) );
  nnd2s1 U15197 ( .DIN1(n13290), .DIN2(n13292), .Q(n14989) );
  nnd2s1 U15198 ( .DIN1(n13480), .DIN2(n13341), .Q(n14667) );
  nnd4s1 U15199 ( .DIN1(n14994), .DIN2(n14995), .DIN3(n14996), .DIN4(n14997), 
        .Q(n14987) );
  nnd2s1 U15200 ( .DIN1(n13371), .DIN2(n14998), .Q(n14997) );
  nnd2s1 U15201 ( .DIN1(n14693), .DIN2(n13557), .Q(n14998) );
  nor2s1 U15202 ( .DIN1(n13330), .DIN2(n13302), .Q(n14693) );
  nnd2s1 U15203 ( .DIN1(n13500), .DIN2(n14999), .Q(n14996) );
  nnd2s1 U15204 ( .DIN1(n13496), .DIN2(n13863), .Q(n14999) );
  nnd2s1 U15205 ( .DIN1(n13304), .DIN2(n15000), .Q(n14995) );
  nnd2s1 U15206 ( .DIN1(n13504), .DIN2(n13324), .Q(n15000) );
  nnd2s1 U15207 ( .DIN1(n13279), .DIN2(n14691), .Q(n14994) );
  nnd2s1 U15208 ( .DIN1(n13504), .DIN2(n13555), .Q(n14691) );
  nnd2s1 U15209 ( .DIN1(n13342), .DIN2(n13275), .Q(n14986) );
  nnd2s1 U15210 ( .DIN1(n13489), .DIN2(n13330), .Q(n14985) );
  hi1s1 U15211 ( .DIN(n13504), .Q(n13330) );
  nor3s1 U15212 ( .DIN1(n15001), .DIN2(n15002), .DIN3(n15003), .Q(n13475) );
  nnd4s1 U15213 ( .DIN1(n13295), .DIN2(n13347), .DIN3(n13335), .DIN4(n15004), 
        .Q(n15003) );
  and3s1 U15214 ( .DIN1(n15005), .DIN2(n14747), .DIN3(n15006), .Q(n15004) );
  nnd2s1 U15215 ( .DIN1(n13279), .DIN2(n13353), .Q(n15006) );
  nnd2s1 U15216 ( .DIN1(n13305), .DIN2(n13341), .Q(n14747) );
  nnd2s1 U15217 ( .DIN1(n13539), .DIN2(n13548), .Q(n15005) );
  nor4s1 U15218 ( .DIN1(n15007), .DIN2(n15008), .DIN3(n15009), .DIN4(n15010), 
        .Q(n13335) );
  nnd4s1 U15219 ( .DIN1(n15011), .DIN2(n15012), .DIN3(n15013), .DIN4(n15014), 
        .Q(n15010) );
  nnd2s1 U15220 ( .DIN1(n13301), .DIN2(n15015), .Q(n15014) );
  nnd2s1 U15221 ( .DIN1(n13505), .DIN2(n13499), .Q(n15015) );
  nor2s1 U15222 ( .DIN1(n15016), .DIN2(n15017), .Q(n15013) );
  nor2s1 U15223 ( .DIN1(n15018), .DIN2(n13326), .Q(n15017) );
  and2s1 U15224 ( .DIN1(n13541), .DIN2(n13523), .Q(n15018) );
  nor2s1 U15225 ( .DIN1(n13489), .DIN2(n13304), .Q(n13523) );
  nor2s1 U15226 ( .DIN1(n15019), .DIN2(n13519), .Q(n15016) );
  nor2s1 U15227 ( .DIN1(n13341), .DIN2(n13369), .Q(n15019) );
  hi1s1 U15228 ( .DIN(n13277), .Q(n13369) );
  nnd2s1 U15229 ( .DIN1(n13553), .DIN2(n15020), .Q(n15012) );
  nnd3s1 U15230 ( .DIN1(n13504), .DIN2(n13742), .DIN3(n13328), .Q(n15020) );
  nnd2s1 U15231 ( .DIN1(n13371), .DIN2(n13357), .Q(n15011) );
  nnd3s1 U15232 ( .DIN1(n15021), .DIN2(n14726), .DIN3(n14651), .Q(n15009) );
  nnd2s1 U15233 ( .DIN1(n13490), .DIN2(n13341), .Q(n14651) );
  nnd2s1 U15234 ( .DIN1(n13353), .DIN2(n13331), .Q(n14726) );
  nnd2s1 U15235 ( .DIN1(n13288), .DIN2(n13293), .Q(n15021) );
  nor2s1 U15236 ( .DIN1(n13749), .DIN2(n13366), .Q(n15008) );
  nor2s1 U15237 ( .DIN1(n13368), .DIN2(n13498), .Q(n15007) );
  nor4s1 U15238 ( .DIN1(n15022), .DIN2(n15023), .DIN3(n15024), .DIN4(n15025), 
        .Q(n13347) );
  nnd4s1 U15239 ( .DIN1(n15026), .DIN2(n15027), .DIN3(n15028), .DIN4(n15029), 
        .Q(n15025) );
  and3s1 U15240 ( .DIN1(n15030), .DIN2(n15031), .DIN3(n15032), .Q(n15029) );
  nnd2s1 U15241 ( .DIN1(n13305), .DIN2(n13359), .Q(n15032) );
  nnd2s1 U15242 ( .DIN1(n13303), .DIN2(n15033), .Q(n15031) );
  nnd2s1 U15243 ( .DIN1(n13495), .DIN2(n13865), .Q(n15033) );
  nnd2s1 U15244 ( .DIN1(n13301), .DIN2(n15034), .Q(n15030) );
  nnd2s1 U15245 ( .DIN1(n13504), .DIN2(n13328), .Q(n15034) );
  nnd2s1 U15246 ( .DIN1(n13358), .DIN2(n15035), .Q(n15028) );
  nnd2s1 U15247 ( .DIN1(n13278), .DIN2(n13541), .Q(n15035) );
  nnd2s1 U15248 ( .DIN1(n13333), .DIN2(n15036), .Q(n15027) );
  nnd2s1 U15249 ( .DIN1(n14694), .DIN2(n13558), .Q(n15036) );
  nnd2s1 U15250 ( .DIN1(n13480), .DIN2(n15037), .Q(n15026) );
  nnd2s1 U15251 ( .DIN1(n14078), .DIN2(n13366), .Q(n15037) );
  nnd3s1 U15252 ( .DIN1(n15038), .DIN2(n15039), .DIN3(n15040), .Q(n15024) );
  nnd2s1 U15253 ( .DIN1(n13548), .DIN2(n13302), .Q(n15040) );
  nnd2s1 U15254 ( .DIN1(n13293), .DIN2(n13342), .Q(n15039) );
  hi1s1 U15255 ( .DIN(n13286), .Q(n13342) );
  nnd2s1 U15256 ( .DIN1(n13490), .DIN2(n13291), .Q(n15038) );
  hi1s1 U15257 ( .DIN(n13328), .Q(n13490) );
  nor2s1 U15258 ( .DIN1(n13277), .DIN2(n13281), .Q(n15023) );
  nor2s1 U15259 ( .DIN1(n13520), .DIN2(n13495), .Q(n15022) );
  nor2s1 U15260 ( .DIN1(n15041), .DIN2(n15042), .Q(n13295) );
  nnd4s1 U15261 ( .DIN1(n15043), .DIN2(n15044), .DIN3(n14761), .DIN4(n15045), 
        .Q(n15042) );
  nnd2s1 U15262 ( .DIN1(n13304), .DIN2(n13289), .Q(n15045) );
  nnd2s1 U15263 ( .DIN1(n13498), .DIN2(n13282), .Q(n13289) );
  nnd2s1 U15264 ( .DIN1(n13333), .DIN2(n13279), .Q(n14761) );
  nnd2s1 U15265 ( .DIN1(n13292), .DIN2(n13302), .Q(n15044) );
  nnd2s1 U15266 ( .DIN1(n13553), .DIN2(n13353), .Q(n15043) );
  hi1s1 U15267 ( .DIN(n13365), .Q(n13553) );
  nnd4s1 U15268 ( .DIN1(n15046), .DIN2(n15047), .DIN3(n15048), .DIN4(n15049), 
        .Q(n15041) );
  nnd2s1 U15269 ( .DIN1(n13331), .DIN2(n15050), .Q(n15049) );
  nnd2s1 U15270 ( .DIN1(n13557), .DIN2(n13328), .Q(n15050) );
  hi1s1 U15271 ( .DIN(n13541), .Q(n13331) );
  nnd2s1 U15272 ( .DIN1(n13341), .DIN2(n15051), .Q(n15048) );
  nnd3s1 U15273 ( .DIN1(n13505), .DIN2(n13520), .DIN3(n13281), .Q(n15051) );
  nnd2s1 U15274 ( .DIN1(n13306), .DIN2(n15052), .Q(n15047) );
  nnd4s1 U15275 ( .DIN1(n13504), .DIN2(n14080), .DIN3(n13324), .DIN4(n13557), 
        .Q(n15052) );
  nnd2s1 U15276 ( .DIN1(n13357), .DIN2(n13744), .Q(n15046) );
  nnd3s1 U15277 ( .DIN1(n15053), .DIN2(n15054), .DIN3(n15055), .Q(n15002) );
  nnd2s1 U15278 ( .DIN1(n13292), .DIN2(n13283), .Q(n15055) );
  hi1s1 U15279 ( .DIN(n13865), .Q(n13292) );
  or2s1 U15280 ( .DIN1(n13368), .DIN2(n13752), .Q(n15054) );
  nor2s1 U15281 ( .DIN1(n13358), .DIN2(n13275), .Q(n13752) );
  hi1s1 U15282 ( .DIN(n13557), .Q(n13275) );
  nnd2s1 U15283 ( .DIN1(n13290), .DIN2(n13359), .Q(n15053) );
  nnd4s1 U15284 ( .DIN1(n15056), .DIN2(n15057), .DIN3(n15058), .DIN4(n15059), 
        .Q(n15001) );
  nnd2s1 U15285 ( .DIN1(n13293), .DIN2(n15060), .Q(n15059) );
  nnd2s1 U15286 ( .DIN1(n14081), .DIN2(n13541), .Q(n15060) );
  nor2s1 U15287 ( .DIN1(n13301), .DIN2(n13306), .Q(n14081) );
  hi1s1 U15288 ( .DIN(n13502), .Q(n13306) );
  nnd2s1 U15289 ( .DIN1(n13288), .DIN2(n15061), .Q(n15058) );
  nnd2s1 U15290 ( .DIN1(n13749), .DIN2(n13328), .Q(n15061) );
  nnd3s1 U15291 ( .DIN1(sa13[5]), .DIN2(sa13[4]), .DIN3(n15062), .Q(n13328) );
  nnd2s1 U15292 ( .DIN1(n13304), .DIN2(n15063), .Q(n15057) );
  nnd2s1 U15293 ( .DIN1(n13499), .DIN2(n13519), .Q(n15063) );
  or2s1 U15294 ( .DIN1(n13365), .DIN2(n14757), .Q(n15056) );
  nor2s1 U15295 ( .DIN1(n13480), .DIN2(n13333), .Q(n14757) );
  nor4s1 U15296 ( .DIN1(n15064), .DIN2(n15065), .DIN3(n15066), .DIN4(n15067), 
        .Q(n13296) );
  nnd4s1 U15297 ( .DIN1(n14746), .DIN2(n15068), .DIN3(n14685), .DIN4(n15069), 
        .Q(n15067) );
  nnd2s1 U15298 ( .DIN1(n13480), .DIN2(n13334), .Q(n15069) );
  nnd2s1 U15299 ( .DIN1(n13277), .DIN2(n13368), .Q(n13334) );
  nnd2s1 U15300 ( .DIN1(n13291), .DIN2(n13353), .Q(n14685) );
  nnd2s1 U15301 ( .DIN1(n13279), .DIN2(n13302), .Q(n15068) );
  nnd2s1 U15302 ( .DIN1(n13304), .DIN2(n13358), .Q(n14746) );
  hi1s1 U15303 ( .DIN(n14694), .Q(n13304) );
  nnd3s1 U15304 ( .DIN1(n15070), .DIN2(n15071), .DIN3(n15072), .Q(n15066) );
  nnd2s1 U15305 ( .DIN1(n13341), .DIN2(n15073), .Q(n15072) );
  nnd2s1 U15306 ( .DIN1(n13499), .DIN2(n13282), .Q(n15073) );
  nnd2s1 U15307 ( .DIN1(n13357), .DIN2(n15074), .Q(n15071) );
  nnd2s1 U15308 ( .DIN1(n13287), .DIN2(n13365), .Q(n15074) );
  nor2s1 U15309 ( .DIN1(n13489), .DIN2(n13291), .Q(n13287) );
  hi1s1 U15310 ( .DIN(n13368), .Q(n13291) );
  nnd2s1 U15311 ( .DIN1(n13359), .DIN2(n15075), .Q(n15070) );
  nnd2s1 U15312 ( .DIN1(n13281), .DIN2(n13504), .Q(n15075) );
  nnd3s1 U15313 ( .DIN1(n1370), .DIN2(n1422), .DIN3(n15076), .Q(n13504) );
  nor2s1 U15314 ( .DIN1(n13559), .DIN2(n13541), .Q(n15065) );
  nor2s1 U15315 ( .DIN1(n13302), .DIN2(n13333), .Q(n13559) );
  nor2s1 U15316 ( .DIN1(n15077), .DIN2(n13557), .Q(n15064) );
  nnd3s1 U15317 ( .DIN1(sa13[7]), .DIN2(n1384), .DIN3(n15078), .Q(n13557) );
  nor2s1 U15318 ( .DIN1(n13288), .DIN2(n13301), .Q(n15077) );
  nor4s1 U15319 ( .DIN1(n15079), .DIN2(n15080), .DIN3(n15081), .DIN4(n15082), 
        .Q(n13336) );
  nnd4s1 U15320 ( .DIN1(n15083), .DIN2(n15084), .DIN3(n15085), .DIN4(n15086), 
        .Q(n15082) );
  nor2s1 U15321 ( .DIN1(n15087), .DIN2(n15088), .Q(n15086) );
  nor2s1 U15322 ( .DIN1(n13519), .DIN2(n13502), .Q(n15088) );
  nor2s1 U15323 ( .DIN1(n13749), .DIN2(n13286), .Q(n15087) );
  nnd3s1 U15324 ( .DIN1(n15089), .DIN2(sa13[0]), .DIN3(sa13[3]), .Q(n13286) );
  nnd2s1 U15325 ( .DIN1(n13371), .DIN2(n13353), .Q(n15085) );
  or2s1 U15326 ( .DIN1(n13368), .DIN2(n14096), .Q(n15084) );
  nor2s1 U15327 ( .DIN1(n13302), .DIN2(n13293), .Q(n14096) );
  hi1s1 U15328 ( .DIN(n13555), .Q(n13293) );
  nnd3s1 U15329 ( .DIN1(n1384), .DIN2(n1422), .DIN3(n15078), .Q(n13555) );
  hi1s1 U15330 ( .DIN(n13519), .Q(n13302) );
  nnd2s1 U15331 ( .DIN1(n13480), .DIN2(n13359), .Q(n15083) );
  hi1s1 U15332 ( .DIN(n13558), .Q(n13359) );
  hi1s1 U15333 ( .DIN(n13326), .Q(n13480) );
  nnd3s1 U15334 ( .DIN1(n15090), .DIN2(n15091), .DIN3(n15092), .Q(n15081) );
  nnd2s1 U15335 ( .DIN1(n13539), .DIN2(n15093), .Q(n15092) );
  nnd2s1 U15336 ( .DIN1(n14694), .DIN2(n13368), .Q(n15093) );
  nnd3s1 U15337 ( .DIN1(sa13[0]), .DIN2(n1436), .DIN3(n15089), .Q(n13368) );
  hi1s1 U15338 ( .DIN(n13281), .Q(n13539) );
  nnd2s1 U15339 ( .DIN1(n13357), .DIN2(n15094), .Q(n15091) );
  nnd2s1 U15340 ( .DIN1(n13541), .DIN2(n13865), .Q(n15094) );
  nnd3s1 U15341 ( .DIN1(n15095), .DIN2(n1358), .DIN3(sa13[3]), .Q(n13865) );
  nnd3s1 U15342 ( .DIN1(sa13[0]), .DIN2(n1386), .DIN3(n15096), .Q(n13541) );
  hi1s1 U15343 ( .DIN(n13324), .Q(n13357) );
  nnd3s1 U15344 ( .DIN1(n15097), .DIN2(n1384), .DIN3(sa13[4]), .Q(n13324) );
  nnd2s1 U15345 ( .DIN1(n13500), .DIN2(n13744), .Q(n15090) );
  nnd2s1 U15346 ( .DIN1(n14078), .DIN2(n13558), .Q(n13744) );
  nnd3s1 U15347 ( .DIN1(sa13[0]), .DIN2(n15095), .DIN3(sa13[3]), .Q(n13558) );
  nor2s1 U15348 ( .DIN1(n15098), .DIN2(n13496), .Q(n15080) );
  nor2s1 U15349 ( .DIN1(n13333), .DIN2(n13358), .Q(n15098) );
  hi1s1 U15350 ( .DIN(n14080), .Q(n13333) );
  nnd2s1 U15351 ( .DIN1(n15099), .DIN2(n15097), .Q(n14080) );
  nor2s1 U15352 ( .DIN1(n15100), .DIN2(n13742), .Q(n15079) );
  nor2s1 U15353 ( .DIN1(n13341), .DIN2(n13288), .Q(n15100) );
  hi1s1 U15354 ( .DIN(n13278), .Q(n13341) );
  nnd3s1 U15355 ( .DIN1(sa13[0]), .DIN2(sa13[2]), .DIN3(n15101), .Q(n13278) );
  nnd3s1 U15356 ( .DIN1(n15102), .DIN2(n15103), .DIN3(n15104), .Q(n14982) );
  nnd2s1 U15357 ( .DIN1(n13548), .DIN2(n13500), .Q(n15104) );
  hi1s1 U15358 ( .DIN(n13520), .Q(n13500) );
  nnd3s1 U15359 ( .DIN1(sa13[5]), .DIN2(n1422), .DIN3(n15078), .Q(n13520) );
  hi1s1 U15360 ( .DIN(n13366), .Q(n13548) );
  nnd3s1 U15361 ( .DIN1(n1358), .DIN2(n1386), .DIN3(n15101), .Q(n13366) );
  nnd2s1 U15362 ( .DIN1(n13283), .DIN2(n13547), .Q(n15103) );
  nnd2s1 U15363 ( .DIN1(n14078), .DIN2(n13365), .Q(n13547) );
  nnd3s1 U15364 ( .DIN1(n15095), .DIN2(n1436), .DIN3(sa13[0]), .Q(n13365) );
  hi1s1 U15365 ( .DIN(n13499), .Q(n13283) );
  nnd3s1 U15366 ( .DIN1(sa13[7]), .DIN2(n1370), .DIN3(n15099), .Q(n13499) );
  nnd2s1 U15367 ( .DIN1(n13290), .DIN2(n13371), .Q(n15102) );
  hi1s1 U15368 ( .DIN(n13285), .Q(n13371) );
  nnd3s1 U15369 ( .DIN1(n1358), .DIN2(n1436), .DIN3(n15089), .Q(n13285) );
  hi1s1 U15370 ( .DIN(n13282), .Q(n13290) );
  nnd2s1 U15371 ( .DIN1(n15062), .DIN2(n15076), .Q(n13282) );
  nnd4s1 U15372 ( .DIN1(n15105), .DIN2(n15106), .DIN3(n15107), .DIN4(n15108), 
        .Q(n14981) );
  nnd2s1 U15373 ( .DIN1(n13288), .DIN2(n15109), .Q(n15108) );
  nnd2s1 U15374 ( .DIN1(n13326), .DIN2(n13519), .Q(n15109) );
  nnd3s1 U15375 ( .DIN1(sa13[5]), .DIN2(sa13[7]), .DIN3(n15078), .Q(n13519) );
  and2s1 U15376 ( .DIN1(sa13[4]), .DIN2(n1370), .Q(n15078) );
  nnd3s1 U15377 ( .DIN1(n1370), .DIN2(n1422), .DIN3(n15099), .Q(n13326) );
  hi1s1 U15378 ( .DIN(n13863), .Q(n13288) );
  nnd3s1 U15379 ( .DIN1(n1358), .DIN2(n1386), .DIN3(n15096), .Q(n13863) );
  nnd2s1 U15380 ( .DIN1(n13353), .DIN2(n15110), .Q(n15107) );
  nnd2s1 U15381 ( .DIN1(n13277), .DIN2(n14694), .Q(n15110) );
  nnd3s1 U15382 ( .DIN1(n15089), .DIN2(n1358), .DIN3(sa13[3]), .Q(n14694) );
  nor2s1 U15383 ( .DIN1(n1506), .DIN2(sa13[2]), .Q(n15089) );
  nnd3s1 U15384 ( .DIN1(sa13[2]), .DIN2(n1358), .DIN3(n15101), .Q(n13277) );
  hi1s1 U15385 ( .DIN(n13505), .Q(n13353) );
  nnd2s1 U15386 ( .DIN1(n15076), .DIN2(n15097), .Q(n13505) );
  nnd2s1 U15387 ( .DIN1(n13358), .DIN2(n15111), .Q(n15106) );
  nnd2s1 U15388 ( .DIN1(n13542), .DIN2(n13502), .Q(n15111) );
  nnd3s1 U15389 ( .DIN1(sa13[2]), .DIN2(n1358), .DIN3(n15096), .Q(n13502) );
  nor2s1 U15390 ( .DIN1(n13489), .DIN2(n13279), .Q(n13542) );
  hi1s1 U15391 ( .DIN(n14078), .Q(n13279) );
  nnd3s1 U15392 ( .DIN1(n1358), .DIN2(n1436), .DIN3(n15095), .Q(n14078) );
  nor2s1 U15393 ( .DIN1(n1386), .DIN2(n1506), .Q(n15095) );
  hi1s1 U15394 ( .DIN(n13495), .Q(n13489) );
  nnd3s1 U15395 ( .DIN1(sa13[0]), .DIN2(n1386), .DIN3(n15101), .Q(n13495) );
  nor2s1 U15396 ( .DIN1(sa13[3]), .DIN2(sa13[1]), .Q(n15101) );
  hi1s1 U15397 ( .DIN(n13749), .Q(n13358) );
  nnd3s1 U15398 ( .DIN1(sa13[7]), .DIN2(n1370), .DIN3(n15076), .Q(n13749) );
  nor2s1 U15399 ( .DIN1(sa13[5]), .DIN2(sa13[4]), .Q(n15076) );
  nnd2s1 U15400 ( .DIN1(n13301), .DIN2(n15112), .Q(n15105) );
  nnd2s1 U15401 ( .DIN1(n14098), .DIN2(n13281), .Q(n15112) );
  nnd3s1 U15402 ( .DIN1(sa13[4]), .DIN2(n15097), .DIN3(sa13[5]), .Q(n13281) );
  nor2s1 U15403 ( .DIN1(n1422), .DIN2(n1370), .Q(n15097) );
  nor2s1 U15404 ( .DIN1(n13305), .DIN2(n13303), .Q(n14098) );
  hi1s1 U15405 ( .DIN(n13742), .Q(n13303) );
  nnd2s1 U15406 ( .DIN1(n15099), .DIN2(n15062), .Q(n13742) );
  nor2s1 U15407 ( .DIN1(n1384), .DIN2(sa13[4]), .Q(n15099) );
  hi1s1 U15408 ( .DIN(n13498), .Q(n13305) );
  nnd3s1 U15409 ( .DIN1(sa13[4]), .DIN2(n1384), .DIN3(n15062), .Q(n13498) );
  nor2s1 U15410 ( .DIN1(n1370), .DIN2(sa13[7]), .Q(n15062) );
  hi1s1 U15411 ( .DIN(n13496), .Q(n13301) );
  nnd3s1 U15412 ( .DIN1(sa13[0]), .DIN2(sa13[2]), .DIN3(n15096), .Q(n13496) );
  nor2s1 U15413 ( .DIN1(n1436), .DIN2(sa13[1]), .Q(n15096) );
  or3s1 U15414 ( .DIN1(n15113), .DIN2(n15114), .DIN3(n15115), .Q(n13070) );
  nnd4s1 U15415 ( .DIN1(n13406), .DIN2(n15116), .DIN3(n14437), .DIN4(n15117), 
        .Q(n15115) );
  and3s1 U15416 ( .DIN1(n15118), .DIN2(n15119), .DIN3(n15120), .Q(n15117) );
  nnd2s1 U15417 ( .DIN1(n14151), .DIN2(n13415), .Q(n15119) );
  nnd2s1 U15418 ( .DIN1(n13397), .DIN2(n13706), .Q(n15118) );
  nor3s1 U15419 ( .DIN1(n15121), .DIN2(n15122), .DIN3(n15123), .Q(n14437) );
  nnd4s1 U15420 ( .DIN1(n15124), .DIN2(n15125), .DIN3(n13405), .DIN4(n15126), 
        .Q(n15123) );
  and3s1 U15421 ( .DIN1(n15127), .DIN2(n15128), .DIN3(n14616), .Q(n15126) );
  nnd2s1 U15422 ( .DIN1(n13414), .DIN2(n13385), .Q(n14616) );
  nnd2s1 U15423 ( .DIN1(n14147), .DIN2(n13397), .Q(n15128) );
  nnd2s1 U15424 ( .DIN1(n13891), .DIN2(n13924), .Q(n15127) );
  nor4s1 U15425 ( .DIN1(n15129), .DIN2(n15130), .DIN3(n15131), .DIN4(n15132), 
        .Q(n13405) );
  nnd4s1 U15426 ( .DIN1(n15133), .DIN2(n15134), .DIN3(n14613), .DIN4(n15135), 
        .Q(n15132) );
  nnd2s1 U15427 ( .DIN1(n13393), .DIN2(n13386), .Q(n15135) );
  nnd2s1 U15428 ( .DIN1(n13387), .DIN2(n13924), .Q(n14613) );
  nnd2s1 U15429 ( .DIN1(n13908), .DIN2(n13706), .Q(n15134) );
  nnd2s1 U15430 ( .DIN1(n13414), .DIN2(n13890), .Q(n15133) );
  nnd3s1 U15431 ( .DIN1(n15136), .DIN2(n15137), .DIN3(n15138), .Q(n15131) );
  nnd2s1 U15432 ( .DIN1(n13385), .DIN2(n14629), .Q(n15138) );
  nnd2s1 U15433 ( .DIN1(n13918), .DIN2(n13401), .Q(n14629) );
  nnd2s1 U15434 ( .DIN1(n13412), .DIN2(n15139), .Q(n15137) );
  nnd2s1 U15435 ( .DIN1(n15140), .DIN2(n14458), .Q(n15139) );
  nnd2s1 U15436 ( .DIN1(n13903), .DIN2(n15141), .Q(n15136) );
  nnd2s1 U15437 ( .DIN1(n13721), .DIN2(n13727), .Q(n15141) );
  nor2s1 U15438 ( .DIN1(n13724), .DIN2(n13400), .Q(n15130) );
  and2s1 U15439 ( .DIN1(n13725), .DIN2(n15142), .Q(n15129) );
  nnd3s1 U15440 ( .DIN1(n13728), .DIN2(n13714), .DIN3(n13401), .Q(n15142) );
  nnd3s1 U15441 ( .DIN1(n15143), .DIN2(n15144), .DIN3(n15145), .Q(n15122) );
  nnd2s1 U15442 ( .DIN1(n13902), .DIN2(n13898), .Q(n15145) );
  or2s1 U15443 ( .DIN1(n14529), .DIN2(n14628), .Q(n15144) );
  nor2s1 U15444 ( .DIN1(n13412), .DIN2(n14214), .Q(n14628) );
  nnd2s1 U15445 ( .DIN1(n13890), .DIN2(n14609), .Q(n15143) );
  nnd2s1 U15446 ( .DIN1(n13720), .DIN2(n13724), .Q(n14609) );
  nnd4s1 U15447 ( .DIN1(n15146), .DIN2(n15147), .DIN3(n15148), .DIN4(n15149), 
        .Q(n15121) );
  nnd2s1 U15448 ( .DIN1(n13386), .DIN2(n15150), .Q(n15149) );
  nnd2s1 U15449 ( .DIN1(n14579), .DIN2(n14458), .Q(n15150) );
  hi1s1 U15450 ( .DIN(n13923), .Q(n14579) );
  nnd2s1 U15451 ( .DIN1(n13399), .DIN2(n13930), .Q(n13923) );
  nnd2s1 U15452 ( .DIN1(n13381), .DIN2(n15151), .Q(n15148) );
  nnd2s1 U15453 ( .DIN1(n13931), .DIN2(n13916), .Q(n15151) );
  nnd2s1 U15454 ( .DIN1(n14166), .DIN2(n15152), .Q(n15147) );
  nnd2s1 U15455 ( .DIN1(n13393), .DIN2(n15153), .Q(n15146) );
  nnd2s1 U15456 ( .DIN1(n13724), .DIN2(n13401), .Q(n15153) );
  nor4s1 U15457 ( .DIN1(n15154), .DIN2(n15155), .DIN3(n15156), .DIN4(n15157), 
        .Q(n13406) );
  nnd4s1 U15458 ( .DIN1(n15158), .DIN2(n15159), .DIN3(n15160), .DIN4(n15161), 
        .Q(n15157) );
  nor2s1 U15459 ( .DIN1(n15162), .DIN2(n15163), .Q(n15161) );
  nor2s1 U15460 ( .DIN1(n15164), .DIN2(n13911), .Q(n15163) );
  and2s1 U15461 ( .DIN1(n13395), .DIN2(n14173), .Q(n15164) );
  nor2s1 U15462 ( .DIN1(n14166), .DIN2(n13386), .Q(n14173) );
  nor2s1 U15463 ( .DIN1(n15165), .DIN2(n13930), .Q(n15162) );
  nor2s1 U15464 ( .DIN1(n14596), .DIN2(n14214), .Q(n15165) );
  nnd2s1 U15465 ( .DIN1(n14165), .DIN2(n15166), .Q(n15160) );
  nnd2s1 U15466 ( .DIN1(n13910), .DIN2(n14456), .Q(n15166) );
  nnd2s1 U15467 ( .DIN1(n14147), .DIN2(n15167), .Q(n15159) );
  nnd2s1 U15468 ( .DIN1(n13914), .DIN2(n13711), .Q(n15167) );
  nnd2s1 U15469 ( .DIN1(n13908), .DIN2(n15168), .Q(n15158) );
  nnd2s1 U15470 ( .DIN1(n14458), .DIN2(n13916), .Q(n15168) );
  nnd3s1 U15471 ( .DIN1(n15169), .DIN2(n15170), .DIN3(n15171), .Q(n15156) );
  nnd2s1 U15472 ( .DIN1(n13706), .DIN2(n13924), .Q(n15171) );
  nnd2s1 U15473 ( .DIN1(n13891), .DIN2(n13901), .Q(n15170) );
  nnd2s1 U15474 ( .DIN1(n14596), .DIN2(n13415), .Q(n15169) );
  nor2s1 U15475 ( .DIN1(n13399), .DIN2(n13918), .Q(n15155) );
  nor2s1 U15476 ( .DIN1(n13931), .DIN2(n13395), .Q(n15154) );
  nnd3s1 U15477 ( .DIN1(n15172), .DIN2(n15173), .DIN3(n15174), .Q(n15114) );
  nnd2s1 U15478 ( .DIN1(n13932), .DIN2(n13388), .Q(n15174) );
  or2s1 U15479 ( .DIN1(n13721), .DIN2(n14473), .Q(n15173) );
  nor2s1 U15480 ( .DIN1(n13891), .DIN2(n13725), .Q(n14473) );
  nnd2s1 U15481 ( .DIN1(n13898), .DIN2(n13901), .Q(n15172) );
  nnd4s1 U15482 ( .DIN1(n15175), .DIN2(n15176), .DIN3(n15177), .DIN4(n15178), 
        .Q(n15113) );
  nnd2s1 U15483 ( .DIN1(n14596), .DIN2(n15179), .Q(n15178) );
  nnd2s1 U15484 ( .DIN1(n14460), .DIN2(n13399), .Q(n15179) );
  nor2s1 U15485 ( .DIN1(n13891), .DIN2(n13932), .Q(n14460) );
  nnd2s1 U15486 ( .DIN1(n13924), .DIN2(n15152), .Q(n15177) );
  nnd2s1 U15487 ( .DIN1(n14146), .DIN2(n13931), .Q(n15152) );
  nnd2s1 U15488 ( .DIN1(n13903), .DIN2(n15180), .Q(n15176) );
  nnd2s1 U15489 ( .DIN1(n14174), .DIN2(n13395), .Q(n15180) );
  nor2s1 U15490 ( .DIN1(n13414), .DIN2(n14165), .Q(n14174) );
  nnd2s1 U15491 ( .DIN1(n13393), .DIN2(n15181), .Q(n15175) );
  nnd2s1 U15492 ( .DIN1(n13918), .DIN2(n13914), .Q(n15181) );
  hi1s1 U15493 ( .DIN(n5225), .Q(n13089) );
  or3s1 U15494 ( .DIN1(n15182), .DIN2(n15183), .DIN3(n15184), .Q(n5225) );
  nnd4s1 U15495 ( .DIN1(n15124), .DIN2(n13408), .DIN3(n14436), .DIN4(n15185), 
        .Q(n15184) );
  and3s1 U15496 ( .DIN1(n15186), .DIN2(n15187), .DIN3(n15116), .Q(n15185) );
  nor4s1 U15497 ( .DIN1(n15188), .DIN2(n15189), .DIN3(n15190), .DIN4(n15191), 
        .Q(n15116) );
  nnd4s1 U15498 ( .DIN1(n15192), .DIN2(n15193), .DIN3(n14617), .DIN4(n15194), 
        .Q(n15191) );
  nnd2s1 U15499 ( .DIN1(n13387), .DIN2(n13384), .Q(n15194) );
  nnd2s1 U15500 ( .DIN1(n13918), .DIN2(n14150), .Q(n13384) );
  nnd2s1 U15501 ( .DIN1(n14596), .DIN2(n13912), .Q(n14617) );
  nnd2s1 U15502 ( .DIN1(n13890), .DIN2(n13924), .Q(n15193) );
  nnd2s1 U15503 ( .DIN1(n13891), .DIN2(n14166), .Q(n15192) );
  nnd3s1 U15504 ( .DIN1(n15195), .DIN2(n15196), .DIN3(n15197), .Q(n15190) );
  nnd2s1 U15505 ( .DIN1(n13385), .DIN2(n15198), .Q(n15197) );
  nnd2s1 U15506 ( .DIN1(n14471), .DIN2(n13721), .Q(n15198) );
  nnd2s1 U15507 ( .DIN1(n14147), .DIN2(n15199), .Q(n15196) );
  nnd2s1 U15508 ( .DIN1(n13395), .DIN2(n13728), .Q(n15199) );
  nnd2s1 U15509 ( .DIN1(n13908), .DIN2(n15200), .Q(n15195) );
  nnd2s1 U15510 ( .DIN1(n13712), .DIN2(n14529), .Q(n15200) );
  nor2s1 U15511 ( .DIN1(n14530), .DIN2(n13914), .Q(n15189) );
  nor2s1 U15512 ( .DIN1(n13890), .DIN2(n13383), .Q(n14530) );
  nor2s1 U15513 ( .DIN1(n15201), .DIN2(n13720), .Q(n15188) );
  nor2s1 U15514 ( .DIN1(n13903), .DIN2(n13393), .Q(n15201) );
  nnd2s1 U15515 ( .DIN1(n13902), .DIN2(n13891), .Q(n15187) );
  nnd2s1 U15516 ( .DIN1(n13903), .DIN2(n14166), .Q(n15186) );
  nor2s1 U15517 ( .DIN1(n15202), .DIN2(n15203), .Q(n14436) );
  nnd4s1 U15518 ( .DIN1(n15204), .DIN2(n15205), .DIN3(n15206), .DIN4(n15207), 
        .Q(n15203) );
  nnd2s1 U15519 ( .DIN1(n13901), .DIN2(n14192), .Q(n15207) );
  nnd2s1 U15520 ( .DIN1(n14529), .DIN2(n13916), .Q(n14192) );
  nnd2s1 U15521 ( .DIN1(n13383), .DIN2(n13388), .Q(n15206) );
  nnd2s1 U15522 ( .DIN1(n13706), .DIN2(n14165), .Q(n15205) );
  nnd2s1 U15523 ( .DIN1(n13393), .DIN2(n13381), .Q(n15204) );
  nnd4s1 U15524 ( .DIN1(n15208), .DIN2(n15209), .DIN3(n15210), .DIN4(n15211), 
        .Q(n15202) );
  nnd2s1 U15525 ( .DIN1(n13707), .DIN2(n15212), .Q(n15211) );
  or2s1 U15526 ( .DIN1(n13382), .DIN2(n13912), .Q(n15212) );
  nnd2s1 U15527 ( .DIN1(n14146), .DIN2(n14200), .Q(n13382) );
  nnd2s1 U15528 ( .DIN1(n13924), .DIN2(n14171), .Q(n15210) );
  nnd2s1 U15529 ( .DIN1(n14200), .DIN2(n13400), .Q(n14171) );
  nnd2s1 U15530 ( .DIN1(n13415), .DIN2(n15213), .Q(n15209) );
  nnd2s1 U15531 ( .DIN1(n13918), .DIN2(n13711), .Q(n15213) );
  nnd2s1 U15532 ( .DIN1(n13386), .DIN2(n15214), .Q(n15208) );
  nnd3s1 U15533 ( .DIN1(n14146), .DIN2(n13400), .DIN3(n15140), .Q(n15214) );
  nor2s1 U15534 ( .DIN1(n13932), .DIN2(n13912), .Q(n15140) );
  nor3s1 U15535 ( .DIN1(n15215), .DIN2(n15216), .DIN3(n15217), .Q(n13408) );
  nnd4s1 U15536 ( .DIN1(n15125), .DIN2(n15120), .DIN3(n14439), .DIN4(n15218), 
        .Q(n15217) );
  and3s1 U15537 ( .DIN1(n15219), .DIN2(n14535), .DIN3(n15220), .Q(n15218) );
  nnd2s1 U15538 ( .DIN1(n13891), .DIN2(n14165), .Q(n15220) );
  nnd2s1 U15539 ( .DIN1(n13397), .DIN2(n13387), .Q(n14535) );
  nnd2s1 U15540 ( .DIN1(n13908), .DIN2(n13385), .Q(n15219) );
  nor4s1 U15541 ( .DIN1(n15221), .DIN2(n15222), .DIN3(n15223), .DIN4(n15224), 
        .Q(n14439) );
  nnd4s1 U15542 ( .DIN1(n15225), .DIN2(n15226), .DIN3(n15227), .DIN4(n15228), 
        .Q(n15224) );
  nnd2s1 U15543 ( .DIN1(n13932), .DIN2(n13707), .Q(n15228) );
  nnd2s1 U15544 ( .DIN1(n14151), .DIN2(n14147), .Q(n15227) );
  nnd2s1 U15545 ( .DIN1(n14214), .DIN2(n13393), .Q(n15226) );
  hi1s1 U15546 ( .DIN(n13910), .Q(n13393) );
  nnd2s1 U15547 ( .DIN1(n13412), .DIN2(n13706), .Q(n15225) );
  nnd3s1 U15548 ( .DIN1(n15229), .DIN2(n15230), .DIN3(n15231), .Q(n15223) );
  nnd2s1 U15549 ( .DIN1(n13397), .DIN2(n15232), .Q(n15231) );
  nnd3s1 U15550 ( .DIN1(n14451), .DIN2(n13930), .DIN3(n14154), .Q(n15232) );
  nnd2s1 U15551 ( .DIN1(n13387), .DIN2(n15233), .Q(n15230) );
  nnd2s1 U15552 ( .DIN1(n14461), .DIN2(n13721), .Q(n15233) );
  nnd2s1 U15553 ( .DIN1(n13890), .DIN2(n15234), .Q(n15229) );
  nor2s1 U15554 ( .DIN1(n13711), .DIN2(n13399), .Q(n15222) );
  and2s1 U15555 ( .DIN1(n13403), .DIN2(n15235), .Q(n15221) );
  nnd4s1 U15556 ( .DIN1(n13401), .DIN2(n13728), .DIN3(n13727), .DIN4(n13395), 
        .Q(n15235) );
  nor2s1 U15557 ( .DIN1(n15236), .DIN2(n15237), .Q(n15120) );
  nnd4s1 U15558 ( .DIN1(n14537), .DIN2(n15238), .DIN3(n15239), .DIN4(n15240), 
        .Q(n15237) );
  nnd2s1 U15559 ( .DIN1(n13891), .DIN2(n14561), .Q(n15240) );
  nnd2s1 U15560 ( .DIN1(n13728), .DIN2(n14459), .Q(n14561) );
  nnd2s1 U15561 ( .DIN1(n13415), .DIN2(n15241), .Q(n15239) );
  nnd3s1 U15562 ( .DIN1(n13714), .DIN2(n13395), .DIN3(n13727), .Q(n15241) );
  nnd2s1 U15563 ( .DIN1(n13397), .DIN2(n13403), .Q(n15238) );
  nnd2s1 U15564 ( .DIN1(n13412), .DIN2(n13385), .Q(n14537) );
  hi1s1 U15565 ( .DIN(n13914), .Q(n13412) );
  nnd4s1 U15566 ( .DIN1(n15242), .DIN2(n15243), .DIN3(n15244), .DIN4(n15245), 
        .Q(n15236) );
  nnd2s1 U15567 ( .DIN1(n13901), .DIN2(n15246), .Q(n15245) );
  nnd2s1 U15568 ( .DIN1(n13910), .DIN2(n13930), .Q(n15246) );
  nnd2s1 U15569 ( .DIN1(n14596), .DIN2(n15247), .Q(n15244) );
  nnd2s1 U15570 ( .DIN1(n14146), .DIN2(n14529), .Q(n15247) );
  nnd2s1 U15571 ( .DIN1(n13912), .DIN2(n15248), .Q(n15243) );
  nnd2s1 U15572 ( .DIN1(n13396), .DIN2(n13728), .Q(n15248) );
  nnd2s1 U15573 ( .DIN1(n13706), .DIN2(n15249), .Q(n15242) );
  nnd2s1 U15574 ( .DIN1(n14563), .DIN2(n13720), .Q(n15249) );
  nor2s1 U15575 ( .DIN1(n14166), .DIN2(n13388), .Q(n14563) );
  and4s1 U15576 ( .DIN1(n15250), .DIN2(n15251), .DIN3(n15252), .DIN4(n15253), 
        .Q(n15125) );
  nor4s1 U15577 ( .DIN1(n15254), .DIN2(n15255), .DIN3(n15256), .DIN4(n15257), 
        .Q(n15253) );
  nor2s1 U15578 ( .DIN1(n15258), .DIN2(n14150), .Q(n15257) );
  nor2s1 U15579 ( .DIN1(n14147), .DIN2(n13912), .Q(n15258) );
  nor2s1 U15580 ( .DIN1(n15259), .DIN2(n13724), .Q(n15256) );
  nor2s1 U15581 ( .DIN1(n13387), .DIN2(n13385), .Q(n15259) );
  nor2s1 U15582 ( .DIN1(n15260), .DIN2(n13914), .Q(n15255) );
  nnd2s1 U15583 ( .DIN1(n15261), .DIN2(n15262), .Q(n13914) );
  nor2s1 U15584 ( .DIN1(n13898), .DIN2(n13891), .Q(n15260) );
  nnd3s1 U15585 ( .DIN1(n15263), .DIN2(n15264), .DIN3(n15265), .Q(n15254) );
  nnd2s1 U15586 ( .DIN1(n13403), .DIN2(n14165), .Q(n15265) );
  nnd2s1 U15587 ( .DIN1(n13932), .DIN2(n15234), .Q(n15264) );
  nnd2s1 U15588 ( .DIN1(n13714), .DIN2(n13711), .Q(n15234) );
  nnd2s1 U15589 ( .DIN1(n13903), .DIN2(n15266), .Q(n15263) );
  nnd2s1 U15590 ( .DIN1(n13728), .DIN2(n13401), .Q(n15266) );
  hi1s1 U15591 ( .DIN(n13930), .Q(n13903) );
  nnd2s1 U15592 ( .DIN1(n15267), .DIN2(n15268), .Q(n13930) );
  and3s1 U15593 ( .DIN1(n15269), .DIN2(n15270), .DIN3(n15271), .Q(n15252) );
  nnd2s1 U15594 ( .DIN1(n13890), .DIN2(n13707), .Q(n15271) );
  hi1s1 U15595 ( .DIN(n13401), .Q(n13707) );
  nnd2s1 U15596 ( .DIN1(n13898), .DIN2(n14166), .Q(n15270) );
  hi1s1 U15597 ( .DIN(n13400), .Q(n13898) );
  nnd2s1 U15598 ( .DIN1(n13386), .DIN2(n13415), .Q(n15269) );
  hi1s1 U15599 ( .DIN(n14154), .Q(n13415) );
  nnd2s1 U15600 ( .DIN1(n13414), .DIN2(n14147), .Q(n15251) );
  nnd2s1 U15601 ( .DIN1(n13902), .DIN2(n13383), .Q(n15250) );
  hi1s1 U15602 ( .DIN(n13395), .Q(n13902) );
  nnd3s1 U15603 ( .DIN1(n15272), .DIN2(n15273), .DIN3(n15274), .Q(n15216) );
  nnd2s1 U15604 ( .DIN1(n13413), .DIN2(n13924), .Q(n15274) );
  nnd2s1 U15605 ( .DIN1(n14151), .DIN2(n13403), .Q(n15273) );
  nnd2s1 U15606 ( .DIN1(n14596), .DIN2(n14147), .Q(n15272) );
  hi1s1 U15607 ( .DIN(n14200), .Q(n14147) );
  hi1s1 U15608 ( .DIN(n13724), .Q(n14596) );
  nnd4s1 U15609 ( .DIN1(n15275), .DIN2(n15276), .DIN3(n15277), .DIN4(n15278), 
        .Q(n15215) );
  nnd2s1 U15610 ( .DIN1(n13414), .DIN2(n15279), .Q(n15278) );
  nnd2s1 U15611 ( .DIN1(n14529), .DIN2(n13400), .Q(n15279) );
  nnd2s1 U15612 ( .DIN1(n13388), .DIN2(n15280), .Q(n15277) );
  nnd4s1 U15613 ( .DIN1(n13911), .DIN2(n14456), .DIN3(n14154), .DIN4(n13400), 
        .Q(n15280) );
  nnd3s1 U15614 ( .DIN1(n1380), .DIN2(n1420), .DIN3(n15281), .Q(n13400) );
  hi1s1 U15615 ( .DIN(n13728), .Q(n13388) );
  nnd2s1 U15616 ( .DIN1(n13383), .DIN2(n14560), .Q(n15276) );
  nnd2s1 U15617 ( .DIN1(n14471), .DIN2(n13714), .Q(n14560) );
  hi1s1 U15618 ( .DIN(n14146), .Q(n13383) );
  nnd2s1 U15619 ( .DIN1(n13706), .DIN2(n14155), .Q(n15275) );
  nnd2s1 U15620 ( .DIN1(n13724), .DIN2(n13711), .Q(n14155) );
  nnd2s1 U15621 ( .DIN1(n15282), .DIN2(n15283), .Q(n13724) );
  hi1s1 U15622 ( .DIN(n14201), .Q(n13706) );
  nor2s1 U15623 ( .DIN1(n15284), .DIN2(n15285), .Q(n15124) );
  nnd4s1 U15624 ( .DIN1(n14512), .DIN2(n15286), .DIN3(n15287), .DIN4(n15288), 
        .Q(n15285) );
  nnd2s1 U15625 ( .DIN1(n13908), .DIN2(n13713), .Q(n15288) );
  nnd2s1 U15626 ( .DIN1(n14153), .DIN2(n14200), .Q(n13713) );
  nnd2s1 U15627 ( .DIN1(n15268), .DIN2(n15289), .Q(n14200) );
  hi1s1 U15628 ( .DIN(n13396), .Q(n13908) );
  nnd2s1 U15629 ( .DIN1(n14166), .DIN2(n13403), .Q(n15287) );
  hi1s1 U15630 ( .DIN(n13918), .Q(n14166) );
  nnd2s1 U15631 ( .DIN1(n15282), .DIN2(n15290), .Q(n13918) );
  nnd2s1 U15632 ( .DIN1(n13725), .DIN2(n13924), .Q(n15286) );
  hi1s1 U15633 ( .DIN(n13727), .Q(n13924) );
  hi1s1 U15634 ( .DIN(n14529), .Q(n13725) );
  nnd3s1 U15635 ( .DIN1(sa02[1]), .DIN2(n1377), .DIN3(n15268), .Q(n14529) );
  nnd2s1 U15636 ( .DIN1(n14214), .DIN2(n13891), .Q(n14512) );
  hi1s1 U15637 ( .DIN(n14153), .Q(n13891) );
  hi1s1 U15638 ( .DIN(n14150), .Q(n14214) );
  nnd4s1 U15639 ( .DIN1(n15291), .DIN2(n15292), .DIN3(n15293), .DIN4(n15294), 
        .Q(n15284) );
  nnd2s1 U15640 ( .DIN1(n13387), .DIN2(n15295), .Q(n15294) );
  nnd2s1 U15641 ( .DIN1(n13720), .DIN2(n13401), .Q(n15295) );
  nnd2s1 U15642 ( .DIN1(n15290), .DIN2(n15296), .Q(n13401) );
  nnd2s1 U15643 ( .DIN1(n13912), .DIN2(n15297), .Q(n15293) );
  nnd2s1 U15644 ( .DIN1(n14471), .DIN2(n14461), .Q(n15297) );
  nnd2s1 U15645 ( .DIN1(n13385), .DIN2(n15298), .Q(n15292) );
  nnd3s1 U15646 ( .DIN1(n13727), .DIN2(n13395), .DIN3(n13711), .Q(n15298) );
  nnd2s1 U15647 ( .DIN1(n15299), .DIN2(n15290), .Q(n13395) );
  nnd2s1 U15648 ( .DIN1(n15299), .DIN2(n15283), .Q(n13727) );
  hi1s1 U15649 ( .DIN(n14456), .Q(n13385) );
  nnd2s1 U15650 ( .DIN1(n13413), .DIN2(n15300), .Q(n15291) );
  nnd4s1 U15651 ( .DIN1(n13728), .DIN2(n13396), .DIN3(n14150), .DIN4(n13720), 
        .Q(n15300) );
  nnd2s1 U15652 ( .DIN1(n15261), .DIN2(n15299), .Q(n14150) );
  nnd2s1 U15653 ( .DIN1(n15301), .DIN2(n15299), .Q(n13396) );
  nor2s1 U15654 ( .DIN1(n1524), .DIN2(n1407), .Q(n15299) );
  nnd2s1 U15655 ( .DIN1(n15262), .DIN2(n15283), .Q(n13728) );
  hi1s1 U15656 ( .DIN(n13399), .Q(n13413) );
  nnd3s1 U15657 ( .DIN1(n14212), .DIN2(n15302), .DIN3(n15303), .Q(n15183) );
  nnd2s1 U15658 ( .DIN1(n13912), .DIN2(n14165), .Q(n15303) );
  hi1s1 U15659 ( .DIN(n13714), .Q(n14165) );
  nnd2s1 U15660 ( .DIN1(n15261), .DIN2(n15296), .Q(n13714) );
  hi1s1 U15661 ( .DIN(n13931), .Q(n13912) );
  nnd3s1 U15662 ( .DIN1(n1380), .DIN2(n1417), .DIN3(n15289), .Q(n13931) );
  nnd2s1 U15663 ( .DIN1(n13403), .DIN2(n13386), .Q(n15302) );
  hi1s1 U15664 ( .DIN(n14459), .Q(n13386) );
  nnd2s1 U15665 ( .DIN1(n15301), .DIN2(n15262), .Q(n14459) );
  hi1s1 U15666 ( .DIN(n13916), .Q(n13403) );
  nnd2s1 U15667 ( .DIN1(n15304), .DIN2(n15289), .Q(n13916) );
  nnd2s1 U15668 ( .DIN1(n13387), .DIN2(n13901), .Q(n14212) );
  hi1s1 U15669 ( .DIN(n13711), .Q(n13901) );
  nnd2s1 U15670 ( .DIN1(n15262), .DIN2(n15290), .Q(n13711) );
  nor2s1 U15671 ( .DIN1(n1525), .DIN2(n1406), .Q(n15290) );
  nor2s1 U15672 ( .DIN1(sa02[7]), .DIN2(sa02[6]), .Q(n15262) );
  hi1s1 U15673 ( .DIN(n14458), .Q(n13387) );
  nnd3s1 U15674 ( .DIN1(sa02[0]), .DIN2(n1417), .DIN3(n15267), .Q(n14458) );
  nnd4s1 U15675 ( .DIN1(n15305), .DIN2(n15306), .DIN3(n15307), .DIN4(n15308), 
        .Q(n15182) );
  nnd2s1 U15676 ( .DIN1(n14151), .DIN2(n15309), .Q(n15308) );
  nnd2s1 U15677 ( .DIN1(n14146), .DIN2(n14456), .Q(n15309) );
  nnd3s1 U15678 ( .DIN1(n1420), .DIN2(n1377), .DIN3(n15268), .Q(n14456) );
  nor2s1 U15679 ( .DIN1(n1417), .DIN2(n1380), .Q(n15268) );
  nnd3s1 U15680 ( .DIN1(n1420), .DIN2(n1377), .DIN3(n15304), .Q(n14146) );
  hi1s1 U15681 ( .DIN(n13720), .Q(n14151) );
  nnd2s1 U15682 ( .DIN1(n15301), .DIN2(n15282), .Q(n13720) );
  nnd2s1 U15683 ( .DIN1(n13414), .DIN2(n15310), .Q(n15307) );
  nnd2s1 U15684 ( .DIN1(n13910), .DIN2(n13399), .Q(n15310) );
  nnd2s1 U15685 ( .DIN1(n15267), .DIN2(n15304), .Q(n13399) );
  hi1s1 U15686 ( .DIN(n14461), .Q(n13414) );
  nnd2s1 U15687 ( .DIN1(n15301), .DIN2(n15296), .Q(n14461) );
  nor2s1 U15688 ( .DIN1(n1406), .DIN2(sa02[5]), .Q(n15301) );
  nnd2s1 U15689 ( .DIN1(n13397), .DIN2(n15311), .Q(n15306) );
  or2s1 U15690 ( .DIN1(n13723), .DIN2(n13890), .Q(n15311) );
  nnd2s1 U15691 ( .DIN1(n13910), .DIN2(n14153), .Q(n13723) );
  nnd3s1 U15692 ( .DIN1(sa02[1]), .DIN2(n1377), .DIN3(n15304), .Q(n14153) );
  nor2s1 U15693 ( .DIN1(n1417), .DIN2(sa02[0]), .Q(n15304) );
  nnd3s1 U15694 ( .DIN1(n1380), .DIN2(n1417), .DIN3(n15267), .Q(n13910) );
  nor2s1 U15695 ( .DIN1(n1377), .DIN2(sa02[1]), .Q(n15267) );
  hi1s1 U15696 ( .DIN(n14471), .Q(n13397) );
  nnd2s1 U15697 ( .DIN1(n15283), .DIN2(n15296), .Q(n14471) );
  nor2s1 U15698 ( .DIN1(n1407), .DIN2(sa02[7]), .Q(n15296) );
  nor2s1 U15699 ( .DIN1(sa02[5]), .DIN2(sa02[4]), .Q(n15283) );
  nnd2s1 U15700 ( .DIN1(n13381), .DIN2(n15312), .Q(n15305) );
  nnd3s1 U15701 ( .DIN1(n14154), .DIN2(n14201), .DIN3(n13712), .Q(n15312) );
  nor2s1 U15702 ( .DIN1(n13890), .DIN2(n13932), .Q(n13712) );
  hi1s1 U15703 ( .DIN(n14451), .Q(n13932) );
  nnd3s1 U15704 ( .DIN1(sa02[0]), .DIN2(n1420), .DIN3(n15281), .Q(n14451) );
  hi1s1 U15705 ( .DIN(n13911), .Q(n13890) );
  nnd3s1 U15706 ( .DIN1(sa02[0]), .DIN2(sa02[1]), .DIN3(n15281), .Q(n13911) );
  nnd3s1 U15707 ( .DIN1(sa02[1]), .DIN2(n1380), .DIN3(n15281), .Q(n14201) );
  nor2s1 U15708 ( .DIN1(sa02[3]), .DIN2(sa02[2]), .Q(n15281) );
  nnd3s1 U15709 ( .DIN1(n15289), .DIN2(n1417), .DIN3(sa02[0]), .Q(n14154) );
  nor2s1 U15710 ( .DIN1(n1377), .DIN2(n1420), .Q(n15289) );
  hi1s1 U15711 ( .DIN(n13721), .Q(n13381) );
  nnd2s1 U15712 ( .DIN1(n15261), .DIN2(n15282), .Q(n13721) );
  nor2s1 U15713 ( .DIN1(n1524), .DIN2(sa02[6]), .Q(n15282) );
  nor2s1 U15714 ( .DIN1(n1525), .DIN2(sa02[4]), .Q(n15261) );
  hi1s1 U15715 ( .DIN(n14974), .Q(n14977) );
  xnr2s1 U15716 ( .DIN1(n15313), .DIN2(n5039), .Q(n14974) );
  or3s1 U15717 ( .DIN1(n15314), .DIN2(n15315), .DIN3(n15316), .Q(n5039) );
  nnd4s1 U15718 ( .DIN1(n13226), .DIN2(n13176), .DIN3(n13564), .DIN4(n15317), 
        .Q(n15316) );
  and3s1 U15719 ( .DIN1(n15318), .DIN2(n15319), .DIN3(n13238), .Q(n15317) );
  nor2s1 U15720 ( .DIN1(n15320), .DIN2(n15321), .Q(n13238) );
  nnd4s1 U15721 ( .DIN1(n14866), .DIN2(n15322), .DIN3(n15323), .DIN4(n15324), 
        .Q(n15321) );
  nnd2s1 U15722 ( .DIN1(n13248), .DIN2(n15325), .Q(n15324) );
  nnd2s1 U15723 ( .DIN1(n13157), .DIN2(n13255), .Q(n15325) );
  nnd2s1 U15724 ( .DIN1(n13232), .DIN2(n15326), .Q(n15323) );
  nnd3s1 U15725 ( .DIN1(n13594), .DIN2(n13824), .DIN3(n13161), .Q(n15326) );
  nnd2s1 U15726 ( .DIN1(n13170), .DIN2(n13172), .Q(n15322) );
  nnd2s1 U15727 ( .DIN1(n13569), .DIN2(n13231), .Q(n14866) );
  nnd4s1 U15728 ( .DIN1(n15327), .DIN2(n15328), .DIN3(n15329), .DIN4(n15330), 
        .Q(n15320) );
  nnd2s1 U15729 ( .DIN1(n13261), .DIN2(n15331), .Q(n15330) );
  nnd2s1 U15730 ( .DIN1(n14892), .DIN2(n13646), .Q(n15331) );
  nor2s1 U15731 ( .DIN1(n13220), .DIN2(n13182), .Q(n14892) );
  nnd2s1 U15732 ( .DIN1(n13589), .DIN2(n15332), .Q(n15329) );
  nnd2s1 U15733 ( .DIN1(n13585), .DIN2(n14040), .Q(n15332) );
  nnd2s1 U15734 ( .DIN1(n13184), .DIN2(n15333), .Q(n15328) );
  nnd2s1 U15735 ( .DIN1(n13593), .DIN2(n13214), .Q(n15333) );
  nnd2s1 U15736 ( .DIN1(n13159), .DIN2(n14890), .Q(n15327) );
  nnd2s1 U15737 ( .DIN1(n13593), .DIN2(n13644), .Q(n14890) );
  nnd2s1 U15738 ( .DIN1(n13232), .DIN2(n13155), .Q(n15319) );
  nnd2s1 U15739 ( .DIN1(n13578), .DIN2(n13220), .Q(n15318) );
  hi1s1 U15740 ( .DIN(n13593), .Q(n13220) );
  nor3s1 U15741 ( .DIN1(n15334), .DIN2(n15335), .DIN3(n15336), .Q(n13564) );
  nnd4s1 U15742 ( .DIN1(n13175), .DIN2(n13237), .DIN3(n13225), .DIN4(n15337), 
        .Q(n15336) );
  and3s1 U15743 ( .DIN1(n15338), .DIN2(n14946), .DIN3(n15339), .Q(n15337) );
  nnd2s1 U15744 ( .DIN1(n13159), .DIN2(n13243), .Q(n15339) );
  nnd2s1 U15745 ( .DIN1(n13185), .DIN2(n13231), .Q(n14946) );
  nnd2s1 U15746 ( .DIN1(n13628), .DIN2(n13637), .Q(n15338) );
  nor4s1 U15747 ( .DIN1(n15340), .DIN2(n15341), .DIN3(n15342), .DIN4(n15343), 
        .Q(n13225) );
  nnd4s1 U15748 ( .DIN1(n15344), .DIN2(n15345), .DIN3(n15346), .DIN4(n15347), 
        .Q(n15343) );
  nnd2s1 U15749 ( .DIN1(n13181), .DIN2(n15348), .Q(n15347) );
  nnd2s1 U15750 ( .DIN1(n13594), .DIN2(n13588), .Q(n15348) );
  nor2s1 U15751 ( .DIN1(n15349), .DIN2(n15350), .Q(n15346) );
  nor2s1 U15752 ( .DIN1(n15351), .DIN2(n13216), .Q(n15350) );
  and2s1 U15753 ( .DIN1(n13630), .DIN2(n13612), .Q(n15351) );
  nor2s1 U15754 ( .DIN1(n13578), .DIN2(n13184), .Q(n13612) );
  nor2s1 U15755 ( .DIN1(n15352), .DIN2(n13608), .Q(n15349) );
  nor2s1 U15756 ( .DIN1(n13231), .DIN2(n13259), .Q(n15352) );
  hi1s1 U15757 ( .DIN(n13157), .Q(n13259) );
  nnd2s1 U15758 ( .DIN1(n13642), .DIN2(n15353), .Q(n15345) );
  nnd3s1 U15759 ( .DIN1(n13593), .DIN2(n13824), .DIN3(n13218), .Q(n15353) );
  nnd2s1 U15760 ( .DIN1(n13261), .DIN2(n13247), .Q(n15344) );
  nnd3s1 U15761 ( .DIN1(n15354), .DIN2(n14925), .DIN3(n14850), .Q(n15342) );
  nnd2s1 U15762 ( .DIN1(n13579), .DIN2(n13231), .Q(n14850) );
  nnd2s1 U15763 ( .DIN1(n13243), .DIN2(n13221), .Q(n14925) );
  nnd2s1 U15764 ( .DIN1(n13168), .DIN2(n13173), .Q(n15354) );
  nor2s1 U15765 ( .DIN1(n13831), .DIN2(n13256), .Q(n15341) );
  nor2s1 U15766 ( .DIN1(n13258), .DIN2(n13587), .Q(n15340) );
  nor4s1 U15767 ( .DIN1(n15355), .DIN2(n15356), .DIN3(n15357), .DIN4(n15358), 
        .Q(n13237) );
  nnd4s1 U15768 ( .DIN1(n15359), .DIN2(n15360), .DIN3(n15361), .DIN4(n15362), 
        .Q(n15358) );
  and3s1 U15769 ( .DIN1(n15363), .DIN2(n15364), .DIN3(n15365), .Q(n15362) );
  nnd2s1 U15770 ( .DIN1(n13185), .DIN2(n13249), .Q(n15365) );
  nnd2s1 U15771 ( .DIN1(n13183), .DIN2(n15366), .Q(n15364) );
  nnd2s1 U15772 ( .DIN1(n13584), .DIN2(n14042), .Q(n15366) );
  nnd2s1 U15773 ( .DIN1(n13181), .DIN2(n15367), .Q(n15363) );
  nnd2s1 U15774 ( .DIN1(n13593), .DIN2(n13218), .Q(n15367) );
  nnd2s1 U15775 ( .DIN1(n13248), .DIN2(n15368), .Q(n15361) );
  nnd2s1 U15776 ( .DIN1(n13158), .DIN2(n13630), .Q(n15368) );
  nnd2s1 U15777 ( .DIN1(n13223), .DIN2(n15369), .Q(n15360) );
  nnd2s1 U15778 ( .DIN1(n14893), .DIN2(n13647), .Q(n15369) );
  nnd2s1 U15779 ( .DIN1(n13569), .DIN2(n15370), .Q(n15359) );
  nnd2s1 U15780 ( .DIN1(n14370), .DIN2(n13256), .Q(n15370) );
  nnd3s1 U15781 ( .DIN1(n15371), .DIN2(n15372), .DIN3(n15373), .Q(n15357) );
  nnd2s1 U15782 ( .DIN1(n13637), .DIN2(n13182), .Q(n15373) );
  nnd2s1 U15783 ( .DIN1(n13173), .DIN2(n13232), .Q(n15372) );
  hi1s1 U15784 ( .DIN(n13166), .Q(n13232) );
  nnd2s1 U15785 ( .DIN1(n13579), .DIN2(n13171), .Q(n15371) );
  hi1s1 U15786 ( .DIN(n13218), .Q(n13579) );
  nor2s1 U15787 ( .DIN1(n13157), .DIN2(n13161), .Q(n15356) );
  nor2s1 U15788 ( .DIN1(n13609), .DIN2(n13584), .Q(n15355) );
  nor2s1 U15789 ( .DIN1(n15374), .DIN2(n15375), .Q(n13175) );
  nnd4s1 U15790 ( .DIN1(n15376), .DIN2(n15377), .DIN3(n14960), .DIN4(n15378), 
        .Q(n15375) );
  nnd2s1 U15791 ( .DIN1(n13184), .DIN2(n13169), .Q(n15378) );
  nnd2s1 U15792 ( .DIN1(n13587), .DIN2(n13162), .Q(n13169) );
  nnd2s1 U15793 ( .DIN1(n13223), .DIN2(n13159), .Q(n14960) );
  nnd2s1 U15794 ( .DIN1(n13172), .DIN2(n13182), .Q(n15377) );
  nnd2s1 U15795 ( .DIN1(n13642), .DIN2(n13243), .Q(n15376) );
  hi1s1 U15796 ( .DIN(n13255), .Q(n13642) );
  nnd4s1 U15797 ( .DIN1(n15379), .DIN2(n15380), .DIN3(n15381), .DIN4(n15382), 
        .Q(n15374) );
  nnd2s1 U15798 ( .DIN1(n13221), .DIN2(n15383), .Q(n15382) );
  nnd2s1 U15799 ( .DIN1(n13646), .DIN2(n13218), .Q(n15383) );
  hi1s1 U15800 ( .DIN(n13630), .Q(n13221) );
  nnd2s1 U15801 ( .DIN1(n13231), .DIN2(n15384), .Q(n15381) );
  nnd3s1 U15802 ( .DIN1(n13594), .DIN2(n13609), .DIN3(n13161), .Q(n15384) );
  nnd2s1 U15803 ( .DIN1(n13186), .DIN2(n15385), .Q(n15380) );
  nnd4s1 U15804 ( .DIN1(n13593), .DIN2(n14372), .DIN3(n13214), .DIN4(n13646), 
        .Q(n15385) );
  nnd2s1 U15805 ( .DIN1(n13247), .DIN2(n13826), .Q(n15379) );
  nnd3s1 U15806 ( .DIN1(n15386), .DIN2(n15387), .DIN3(n15388), .Q(n15335) );
  nnd2s1 U15807 ( .DIN1(n13172), .DIN2(n13163), .Q(n15388) );
  hi1s1 U15808 ( .DIN(n14042), .Q(n13172) );
  or2s1 U15809 ( .DIN1(n13258), .DIN2(n13834), .Q(n15387) );
  nor2s1 U15810 ( .DIN1(n13248), .DIN2(n13155), .Q(n13834) );
  hi1s1 U15811 ( .DIN(n13646), .Q(n13155) );
  nnd2s1 U15812 ( .DIN1(n13170), .DIN2(n13249), .Q(n15386) );
  nnd4s1 U15813 ( .DIN1(n15389), .DIN2(n15390), .DIN3(n15391), .DIN4(n15392), 
        .Q(n15334) );
  nnd2s1 U15814 ( .DIN1(n13173), .DIN2(n15393), .Q(n15392) );
  nnd2s1 U15815 ( .DIN1(n14373), .DIN2(n13630), .Q(n15393) );
  nor2s1 U15816 ( .DIN1(n13181), .DIN2(n13186), .Q(n14373) );
  hi1s1 U15817 ( .DIN(n13591), .Q(n13186) );
  nnd2s1 U15818 ( .DIN1(n13168), .DIN2(n15394), .Q(n15391) );
  nnd2s1 U15819 ( .DIN1(n13831), .DIN2(n13218), .Q(n15394) );
  nnd3s1 U15820 ( .DIN1(sa20[5]), .DIN2(sa20[4]), .DIN3(n15395), .Q(n13218) );
  nnd2s1 U15821 ( .DIN1(n13184), .DIN2(n15396), .Q(n15390) );
  nnd2s1 U15822 ( .DIN1(n13588), .DIN2(n13608), .Q(n15396) );
  or2s1 U15823 ( .DIN1(n13255), .DIN2(n14956), .Q(n15389) );
  nor2s1 U15824 ( .DIN1(n13569), .DIN2(n13223), .Q(n14956) );
  nor4s1 U15825 ( .DIN1(n15397), .DIN2(n15398), .DIN3(n15399), .DIN4(n15400), 
        .Q(n13176) );
  nnd4s1 U15826 ( .DIN1(n14945), .DIN2(n15401), .DIN3(n14884), .DIN4(n15402), 
        .Q(n15400) );
  nnd2s1 U15827 ( .DIN1(n13569), .DIN2(n13224), .Q(n15402) );
  nnd2s1 U15828 ( .DIN1(n13157), .DIN2(n13258), .Q(n13224) );
  nnd2s1 U15829 ( .DIN1(n13171), .DIN2(n13243), .Q(n14884) );
  nnd2s1 U15830 ( .DIN1(n13159), .DIN2(n13182), .Q(n15401) );
  nnd2s1 U15831 ( .DIN1(n13184), .DIN2(n13248), .Q(n14945) );
  hi1s1 U15832 ( .DIN(n14893), .Q(n13184) );
  nnd3s1 U15833 ( .DIN1(n15403), .DIN2(n15404), .DIN3(n15405), .Q(n15399) );
  nnd2s1 U15834 ( .DIN1(n13231), .DIN2(n15406), .Q(n15405) );
  nnd2s1 U15835 ( .DIN1(n13588), .DIN2(n13162), .Q(n15406) );
  nnd2s1 U15836 ( .DIN1(n13247), .DIN2(n15407), .Q(n15404) );
  nnd2s1 U15837 ( .DIN1(n13167), .DIN2(n13255), .Q(n15407) );
  nor2s1 U15838 ( .DIN1(n13578), .DIN2(n13171), .Q(n13167) );
  hi1s1 U15839 ( .DIN(n13258), .Q(n13171) );
  nnd2s1 U15840 ( .DIN1(n13249), .DIN2(n15408), .Q(n15403) );
  nnd2s1 U15841 ( .DIN1(n13161), .DIN2(n13593), .Q(n15408) );
  nnd3s1 U15842 ( .DIN1(n1371), .DIN2(n1423), .DIN3(n15409), .Q(n13593) );
  nor2s1 U15843 ( .DIN1(n13648), .DIN2(n13630), .Q(n15398) );
  nor2s1 U15844 ( .DIN1(n13182), .DIN2(n13223), .Q(n13648) );
  nor2s1 U15845 ( .DIN1(n15410), .DIN2(n13646), .Q(n15397) );
  nnd3s1 U15846 ( .DIN1(sa20[7]), .DIN2(n1385), .DIN3(n15411), .Q(n13646) );
  nor2s1 U15847 ( .DIN1(n13168), .DIN2(n13181), .Q(n15410) );
  nor4s1 U15848 ( .DIN1(n15412), .DIN2(n15413), .DIN3(n15414), .DIN4(n15415), 
        .Q(n13226) );
  nnd4s1 U15849 ( .DIN1(n15416), .DIN2(n15417), .DIN3(n15418), .DIN4(n15419), 
        .Q(n15415) );
  nor2s1 U15850 ( .DIN1(n15420), .DIN2(n15421), .Q(n15419) );
  nor2s1 U15851 ( .DIN1(n13608), .DIN2(n13591), .Q(n15421) );
  nor2s1 U15852 ( .DIN1(n13831), .DIN2(n13166), .Q(n15420) );
  nnd3s1 U15853 ( .DIN1(n15422), .DIN2(sa20[0]), .DIN3(sa20[3]), .Q(n13166) );
  nnd2s1 U15854 ( .DIN1(n13261), .DIN2(n13243), .Q(n15418) );
  or2s1 U15855 ( .DIN1(n13258), .DIN2(n14388), .Q(n15417) );
  nor2s1 U15856 ( .DIN1(n13182), .DIN2(n13173), .Q(n14388) );
  hi1s1 U15857 ( .DIN(n13644), .Q(n13173) );
  nnd3s1 U15858 ( .DIN1(n1385), .DIN2(n1423), .DIN3(n15411), .Q(n13644) );
  hi1s1 U15859 ( .DIN(n13608), .Q(n13182) );
  nnd2s1 U15860 ( .DIN1(n13569), .DIN2(n13249), .Q(n15416) );
  hi1s1 U15861 ( .DIN(n13647), .Q(n13249) );
  hi1s1 U15862 ( .DIN(n13216), .Q(n13569) );
  nnd3s1 U15863 ( .DIN1(n15423), .DIN2(n15424), .DIN3(n15425), .Q(n15414) );
  nnd2s1 U15864 ( .DIN1(n13628), .DIN2(n15426), .Q(n15425) );
  nnd2s1 U15865 ( .DIN1(n14893), .DIN2(n13258), .Q(n15426) );
  nnd3s1 U15866 ( .DIN1(sa20[0]), .DIN2(n1437), .DIN3(n15422), .Q(n13258) );
  hi1s1 U15867 ( .DIN(n13161), .Q(n13628) );
  nnd2s1 U15868 ( .DIN1(n13247), .DIN2(n15427), .Q(n15424) );
  nnd2s1 U15869 ( .DIN1(n13630), .DIN2(n14042), .Q(n15427) );
  nnd3s1 U15870 ( .DIN1(n15428), .DIN2(n1359), .DIN3(sa20[3]), .Q(n14042) );
  nnd3s1 U15871 ( .DIN1(sa20[0]), .DIN2(n1387), .DIN3(n15429), .Q(n13630) );
  hi1s1 U15872 ( .DIN(n13214), .Q(n13247) );
  nnd3s1 U15873 ( .DIN1(n15430), .DIN2(n1385), .DIN3(sa20[4]), .Q(n13214) );
  nnd2s1 U15874 ( .DIN1(n13589), .DIN2(n13826), .Q(n15423) );
  nnd2s1 U15875 ( .DIN1(n14370), .DIN2(n13647), .Q(n13826) );
  nnd3s1 U15876 ( .DIN1(sa20[0]), .DIN2(n15428), .DIN3(sa20[3]), .Q(n13647) );
  nor2s1 U15877 ( .DIN1(n15431), .DIN2(n13585), .Q(n15413) );
  nor2s1 U15878 ( .DIN1(n13223), .DIN2(n13248), .Q(n15431) );
  hi1s1 U15879 ( .DIN(n14372), .Q(n13223) );
  nnd2s1 U15880 ( .DIN1(n15432), .DIN2(n15430), .Q(n14372) );
  nor2s1 U15881 ( .DIN1(n15433), .DIN2(n13824), .Q(n15412) );
  nor2s1 U15882 ( .DIN1(n13231), .DIN2(n13168), .Q(n15433) );
  hi1s1 U15883 ( .DIN(n13158), .Q(n13231) );
  nnd3s1 U15884 ( .DIN1(sa20[0]), .DIN2(sa20[2]), .DIN3(n15434), .Q(n13158) );
  nnd3s1 U15885 ( .DIN1(n15435), .DIN2(n15436), .DIN3(n15437), .Q(n15315) );
  nnd2s1 U15886 ( .DIN1(n13637), .DIN2(n13589), .Q(n15437) );
  hi1s1 U15887 ( .DIN(n13609), .Q(n13589) );
  nnd3s1 U15888 ( .DIN1(sa20[5]), .DIN2(n1423), .DIN3(n15411), .Q(n13609) );
  hi1s1 U15889 ( .DIN(n13256), .Q(n13637) );
  nnd3s1 U15890 ( .DIN1(n1359), .DIN2(n1387), .DIN3(n15434), .Q(n13256) );
  nnd2s1 U15891 ( .DIN1(n13163), .DIN2(n13636), .Q(n15436) );
  nnd2s1 U15892 ( .DIN1(n14370), .DIN2(n13255), .Q(n13636) );
  nnd3s1 U15893 ( .DIN1(n15428), .DIN2(n1437), .DIN3(sa20[0]), .Q(n13255) );
  hi1s1 U15894 ( .DIN(n13588), .Q(n13163) );
  nnd3s1 U15895 ( .DIN1(sa20[7]), .DIN2(n1371), .DIN3(n15432), .Q(n13588) );
  nnd2s1 U15896 ( .DIN1(n13170), .DIN2(n13261), .Q(n15435) );
  hi1s1 U15897 ( .DIN(n13165), .Q(n13261) );
  nnd3s1 U15898 ( .DIN1(n1359), .DIN2(n1437), .DIN3(n15422), .Q(n13165) );
  hi1s1 U15899 ( .DIN(n13162), .Q(n13170) );
  nnd2s1 U15900 ( .DIN1(n15395), .DIN2(n15409), .Q(n13162) );
  nnd4s1 U15901 ( .DIN1(n15438), .DIN2(n15439), .DIN3(n15440), .DIN4(n15441), 
        .Q(n15314) );
  nnd2s1 U15902 ( .DIN1(n13168), .DIN2(n15442), .Q(n15441) );
  nnd2s1 U15903 ( .DIN1(n13216), .DIN2(n13608), .Q(n15442) );
  nnd3s1 U15904 ( .DIN1(sa20[5]), .DIN2(sa20[7]), .DIN3(n15411), .Q(n13608) );
  and2s1 U15905 ( .DIN1(sa20[4]), .DIN2(n1371), .Q(n15411) );
  nnd3s1 U15906 ( .DIN1(n1371), .DIN2(n1423), .DIN3(n15432), .Q(n13216) );
  hi1s1 U15907 ( .DIN(n14040), .Q(n13168) );
  nnd3s1 U15908 ( .DIN1(n1359), .DIN2(n1387), .DIN3(n15429), .Q(n14040) );
  nnd2s1 U15909 ( .DIN1(n13243), .DIN2(n15443), .Q(n15440) );
  nnd2s1 U15910 ( .DIN1(n13157), .DIN2(n14893), .Q(n15443) );
  nnd3s1 U15911 ( .DIN1(n15422), .DIN2(n1359), .DIN3(sa20[3]), .Q(n14893) );
  nor2s1 U15912 ( .DIN1(n1507), .DIN2(sa20[2]), .Q(n15422) );
  nnd3s1 U15913 ( .DIN1(sa20[2]), .DIN2(n1359), .DIN3(n15434), .Q(n13157) );
  hi1s1 U15914 ( .DIN(n13594), .Q(n13243) );
  nnd2s1 U15915 ( .DIN1(n15409), .DIN2(n15430), .Q(n13594) );
  nnd2s1 U15916 ( .DIN1(n13248), .DIN2(n15444), .Q(n15439) );
  nnd2s1 U15917 ( .DIN1(n13631), .DIN2(n13591), .Q(n15444) );
  nnd3s1 U15918 ( .DIN1(sa20[2]), .DIN2(n1359), .DIN3(n15429), .Q(n13591) );
  nor2s1 U15919 ( .DIN1(n13578), .DIN2(n13159), .Q(n13631) );
  hi1s1 U15920 ( .DIN(n14370), .Q(n13159) );
  nnd3s1 U15921 ( .DIN1(n1359), .DIN2(n1437), .DIN3(n15428), .Q(n14370) );
  nor2s1 U15922 ( .DIN1(n1387), .DIN2(n1507), .Q(n15428) );
  hi1s1 U15923 ( .DIN(n13584), .Q(n13578) );
  nnd3s1 U15924 ( .DIN1(sa20[0]), .DIN2(n1387), .DIN3(n15434), .Q(n13584) );
  nor2s1 U15925 ( .DIN1(sa20[3]), .DIN2(sa20[1]), .Q(n15434) );
  hi1s1 U15926 ( .DIN(n13831), .Q(n13248) );
  nnd3s1 U15927 ( .DIN1(sa20[7]), .DIN2(n1371), .DIN3(n15409), .Q(n13831) );
  nor2s1 U15928 ( .DIN1(sa20[5]), .DIN2(sa20[4]), .Q(n15409) );
  nnd2s1 U15929 ( .DIN1(n13181), .DIN2(n15445), .Q(n15438) );
  nnd2s1 U15930 ( .DIN1(n14390), .DIN2(n13161), .Q(n15445) );
  nnd3s1 U15931 ( .DIN1(sa20[4]), .DIN2(n15430), .DIN3(sa20[5]), .Q(n13161) );
  nor2s1 U15932 ( .DIN1(n1423), .DIN2(n1371), .Q(n15430) );
  nor2s1 U15933 ( .DIN1(n13185), .DIN2(n13183), .Q(n14390) );
  hi1s1 U15934 ( .DIN(n13824), .Q(n13183) );
  nnd2s1 U15935 ( .DIN1(n15432), .DIN2(n15395), .Q(n13824) );
  nor2s1 U15936 ( .DIN1(n1385), .DIN2(sa20[4]), .Q(n15432) );
  hi1s1 U15937 ( .DIN(n13587), .Q(n13185) );
  nnd3s1 U15938 ( .DIN1(sa20[4]), .DIN2(n1385), .DIN3(n15395), .Q(n13587) );
  nor2s1 U15939 ( .DIN1(n1371), .DIN2(sa20[7]), .Q(n15395) );
  hi1s1 U15940 ( .DIN(n13585), .Q(n13181) );
  nnd3s1 U15941 ( .DIN1(sa20[0]), .DIN2(sa20[2]), .DIN3(n15429), .Q(n13585) );
  nor2s1 U15942 ( .DIN1(n1437), .DIN2(sa20[1]), .Q(n15429) );
  xor2s1 U15943 ( .DIN1(n5015), .DIN2(w2[2]), .Q(n15313) );
  or3s1 U15944 ( .DIN1(n15446), .DIN2(n15447), .DIN3(n15448), .Q(n5015) );
  nnd4s1 U15945 ( .DIN1(n15449), .DIN2(n15450), .DIN3(n13451), .DIN4(n15451), 
        .Q(n15448) );
  and3s1 U15946 ( .DIN1(n14478), .DIN2(n14800), .DIN3(n14773), .Q(n15451) );
  nor4s1 U15947 ( .DIN1(n15452), .DIN2(n15453), .DIN3(n15454), .DIN4(n15455), 
        .Q(n14773) );
  nnd4s1 U15948 ( .DIN1(n15456), .DIN2(n15457), .DIN3(n14333), .DIN4(n15458), 
        .Q(n15455) );
  nnd2s1 U15949 ( .DIN1(n13431), .DIN2(n13427), .Q(n15458) );
  nnd2s1 U15950 ( .DIN1(n13793), .DIN2(n13953), .Q(n13427) );
  nnd2s1 U15951 ( .DIN1(n13787), .DIN2(n14311), .Q(n14333) );
  nnd2s1 U15952 ( .DIN1(n13799), .DIN2(n13765), .Q(n15457) );
  nnd2s1 U15953 ( .DIN1(n13766), .DIN2(n13969), .Q(n15456) );
  nnd3s1 U15954 ( .DIN1(n15459), .DIN2(n15460), .DIN3(n15461), .Q(n15454) );
  nnd2s1 U15955 ( .DIN1(n13428), .DIN2(n15462), .Q(n15461) );
  nnd2s1 U15956 ( .DIN1(n14234), .DIN2(n13674), .Q(n15462) );
  nnd2s1 U15957 ( .DIN1(n13950), .DIN2(n15463), .Q(n15460) );
  nnd2s1 U15958 ( .DIN1(n13438), .DIN2(n13681), .Q(n15463) );
  nnd2s1 U15959 ( .DIN1(n13783), .DIN2(n15464), .Q(n15459) );
  nnd2s1 U15960 ( .DIN1(n13665), .DIN2(n14232), .Q(n15464) );
  nor2s1 U15961 ( .DIN1(n14233), .DIN2(n13789), .Q(n15453) );
  nor2s1 U15962 ( .DIN1(n13765), .DIN2(n13426), .Q(n14233) );
  nor2s1 U15963 ( .DIN1(n15465), .DIN2(n13673), .Q(n15452) );
  nor2s1 U15964 ( .DIN1(n13778), .DIN2(n13436), .Q(n15465) );
  nor2s1 U15965 ( .DIN1(n15466), .DIN2(n15467), .Q(n14800) );
  nnd4s1 U15966 ( .DIN1(n14220), .DIN2(n15468), .DIN3(n15469), .DIN4(n15470), 
        .Q(n15467) );
  nnd2s1 U15967 ( .DIN1(n13783), .DIN2(n13666), .Q(n15470) );
  nnd2s1 U15968 ( .DIN1(n13956), .DIN2(n14004), .Q(n13666) );
  nnd2s1 U15969 ( .DIN1(n13446), .DIN2(n13969), .Q(n15469) );
  nnd2s1 U15970 ( .DIN1(n13799), .DIN2(n13678), .Q(n15468) );
  hi1s1 U15971 ( .DIN(n14232), .Q(n13678) );
  nnd2s1 U15972 ( .DIN1(n13766), .DIN2(n14017), .Q(n14220) );
  nnd4s1 U15973 ( .DIN1(n15471), .DIN2(n15472), .DIN3(n15473), .DIN4(n15474), 
        .Q(n15466) );
  nnd2s1 U15974 ( .DIN1(n13431), .DIN2(n15475), .Q(n15474) );
  nnd2s1 U15975 ( .DIN1(n13673), .DIN2(n13444), .Q(n15475) );
  nnd2s1 U15976 ( .DIN1(n13787), .DIN2(n15476), .Q(n15473) );
  nnd2s1 U15977 ( .DIN1(n14234), .DIN2(n14257), .Q(n15476) );
  nnd2s1 U15978 ( .DIN1(n13428), .DIN2(n15477), .Q(n15472) );
  nnd3s1 U15979 ( .DIN1(n13680), .DIN2(n13438), .DIN3(n13664), .Q(n15477) );
  nnd2s1 U15980 ( .DIN1(n13456), .DIN2(n15478), .Q(n15471) );
  nnd4s1 U15981 ( .DIN1(n13439), .DIN2(n13673), .DIN3(n13681), .DIN4(n13953), 
        .Q(n15478) );
  nor2s1 U15982 ( .DIN1(n15479), .DIN2(n15480), .Q(n14478) );
  nnd4s1 U15983 ( .DIN1(n15481), .DIN2(n15482), .DIN3(n15483), .DIN4(n15484), 
        .Q(n15480) );
  nnd2s1 U15984 ( .DIN1(n13776), .DIN2(n13995), .Q(n15484) );
  nnd2s1 U15985 ( .DIN1(n14232), .DIN2(n13791), .Q(n13995) );
  nnd2s1 U15986 ( .DIN1(n13430), .DIN2(n13426), .Q(n15483) );
  nnd2s1 U15987 ( .DIN1(n13968), .DIN2(n13660), .Q(n15482) );
  nnd2s1 U15988 ( .DIN1(n13436), .DIN2(n13424), .Q(n15481) );
  nnd4s1 U15989 ( .DIN1(n15485), .DIN2(n15486), .DIN3(n15487), .DIN4(n15488), 
        .Q(n15479) );
  nnd2s1 U15990 ( .DIN1(n13659), .DIN2(n15489), .Q(n15488) );
  or2s1 U15991 ( .DIN1(n13425), .DIN2(n13787), .Q(n15489) );
  nnd2s1 U15992 ( .DIN1(n13949), .DIN2(n14004), .Q(n13425) );
  nnd2s1 U15993 ( .DIN1(n13799), .DIN2(n13974), .Q(n15487) );
  nnd2s1 U15994 ( .DIN1(n14004), .DIN2(n13443), .Q(n13974) );
  nnd2s1 U15995 ( .DIN1(n13458), .DIN2(n15490), .Q(n15486) );
  nnd2s1 U15996 ( .DIN1(n13793), .DIN2(n13664), .Q(n15490) );
  nnd2s1 U15997 ( .DIN1(n13429), .DIN2(n15491), .Q(n15485) );
  nnd3s1 U15998 ( .DIN1(n13443), .DIN2(n13949), .DIN3(n14815), .Q(n15491) );
  nor2s1 U15999 ( .DIN1(n13807), .DIN2(n13787), .Q(n14815) );
  nor3s1 U16000 ( .DIN1(n15492), .DIN2(n15493), .DIN3(n15494), .Q(n13451) );
  nnd4s1 U16001 ( .DIN1(n14480), .DIN2(n14799), .DIN3(n14777), .DIN4(n15495), 
        .Q(n15494) );
  and3s1 U16002 ( .DIN1(n15496), .DIN2(n14245), .DIN3(n15497), .Q(n15495) );
  nnd2s1 U16003 ( .DIN1(n13766), .DIN2(n13968), .Q(n15497) );
  nnd2s1 U16004 ( .DIN1(n13440), .DIN2(n13431), .Q(n14245) );
  nnd2s1 U16005 ( .DIN1(n13428), .DIN2(n13783), .Q(n15496) );
  hi1s1 U16006 ( .DIN(n13439), .Q(n13783) );
  nor2s1 U16007 ( .DIN1(n15498), .DIN2(n15499), .Q(n14777) );
  nnd4s1 U16008 ( .DIN1(n14247), .DIN2(n15500), .DIN3(n15501), .DIN4(n15502), 
        .Q(n15499) );
  nnd2s1 U16009 ( .DIN1(n13766), .DIN2(n14274), .Q(n15502) );
  nnd2s1 U16010 ( .DIN1(n13681), .DIN2(n14277), .Q(n14274) );
  nnd2s1 U16011 ( .DIN1(n13458), .DIN2(n15503), .Q(n15501) );
  nnd3s1 U16012 ( .DIN1(n13667), .DIN2(n13438), .DIN3(n13680), .Q(n15503) );
  nnd2s1 U16013 ( .DIN1(n13440), .DIN2(n13446), .Q(n15500) );
  nnd2s1 U16014 ( .DIN1(n13428), .DIN2(n13455), .Q(n14247) );
  nnd4s1 U16015 ( .DIN1(n15504), .DIN2(n15505), .DIN3(n15506), .DIN4(n15507), 
        .Q(n15498) );
  nnd2s1 U16016 ( .DIN1(n13776), .DIN2(n15508), .Q(n15507) );
  nnd2s1 U16017 ( .DIN1(n13785), .DIN2(n13805), .Q(n15508) );
  nnd2s1 U16018 ( .DIN1(n14311), .DIN2(n15509), .Q(n15506) );
  nnd2s1 U16019 ( .DIN1(n13949), .DIN2(n14232), .Q(n15509) );
  nnd2s1 U16020 ( .DIN1(n13787), .DIN2(n15510), .Q(n15505) );
  nnd2s1 U16021 ( .DIN1(n13439), .DIN2(n13681), .Q(n15510) );
  nnd2s1 U16022 ( .DIN1(n15511), .DIN2(n15512), .Q(n13439) );
  nnd2s1 U16023 ( .DIN1(n13660), .DIN2(n15513), .Q(n15504) );
  nnd2s1 U16024 ( .DIN1(n14276), .DIN2(n13673), .Q(n15513) );
  nor2s1 U16025 ( .DIN1(n13969), .DIN2(n13430), .Q(n14276) );
  and4s1 U16026 ( .DIN1(n15514), .DIN2(n15515), .DIN3(n15516), .DIN4(n15517), 
        .Q(n14799) );
  nor4s1 U16027 ( .DIN1(n15518), .DIN2(n15519), .DIN3(n15520), .DIN4(n15521), 
        .Q(n15517) );
  nor2s1 U16028 ( .DIN1(n15522), .DIN2(n13953), .Q(n15521) );
  nor2s1 U16029 ( .DIN1(n13950), .DIN2(n13787), .Q(n15522) );
  nor2s1 U16030 ( .DIN1(n15523), .DIN2(n13677), .Q(n15520) );
  nor2s1 U16031 ( .DIN1(n13431), .DIN2(n13428), .Q(n15523) );
  hi1s1 U16032 ( .DIN(n14323), .Q(n13428) );
  nor2s1 U16033 ( .DIN1(n15524), .DIN2(n13789), .Q(n15519) );
  nor2s1 U16034 ( .DIN1(n13773), .DIN2(n13766), .Q(n15524) );
  nnd3s1 U16035 ( .DIN1(n15525), .DIN2(n15526), .DIN3(n15527), .Q(n15518) );
  nnd2s1 U16036 ( .DIN1(n13446), .DIN2(n13968), .Q(n15527) );
  nnd2s1 U16037 ( .DIN1(n13807), .DIN2(n15528), .Q(n15526) );
  nnd2s1 U16038 ( .DIN1(n13778), .DIN2(n15529), .Q(n15525) );
  nnd2s1 U16039 ( .DIN1(n13681), .DIN2(n13444), .Q(n15529) );
  and3s1 U16040 ( .DIN1(n15530), .DIN2(n15531), .DIN3(n15532), .Q(n15516) );
  nnd2s1 U16041 ( .DIN1(n13659), .DIN2(n13765), .Q(n15532) );
  nnd2s1 U16042 ( .DIN1(n13773), .DIN2(n13969), .Q(n15531) );
  hi1s1 U16043 ( .DIN(n13443), .Q(n13773) );
  nnd2s1 U16044 ( .DIN1(n13429), .DIN2(n13458), .Q(n15530) );
  hi1s1 U16045 ( .DIN(n13957), .Q(n13458) );
  nnd2s1 U16046 ( .DIN1(n13950), .DIN2(n13457), .Q(n15515) );
  nnd2s1 U16047 ( .DIN1(n13426), .DIN2(n13777), .Q(n15514) );
  nor4s1 U16048 ( .DIN1(n15533), .DIN2(n15534), .DIN3(n15535), .DIN4(n15536), 
        .Q(n14480) );
  nnd4s1 U16049 ( .DIN1(n15537), .DIN2(n15538), .DIN3(n15539), .DIN4(n15540), 
        .Q(n15536) );
  nnd2s1 U16050 ( .DIN1(n13659), .DIN2(n13807), .Q(n15540) );
  hi1s1 U16051 ( .DIN(n13444), .Q(n13659) );
  nnd2s1 U16052 ( .DIN1(n13950), .DIN2(n13954), .Q(n15539) );
  nnd2s1 U16053 ( .DIN1(n13436), .DIN2(n14017), .Q(n15538) );
  hi1s1 U16054 ( .DIN(n13953), .Q(n14017) );
  nnd2s1 U16055 ( .DIN1(n15541), .DIN2(n15512), .Q(n13953) );
  hi1s1 U16056 ( .DIN(n13785), .Q(n13436) );
  nnd2s1 U16057 ( .DIN1(n13455), .DIN2(n13660), .Q(n15537) );
  hi1s1 U16058 ( .DIN(n13789), .Q(n13455) );
  nnd2s1 U16059 ( .DIN1(n15542), .DIN2(n15541), .Q(n13789) );
  nnd3s1 U16060 ( .DIN1(n15543), .DIN2(n15544), .DIN3(n15545), .Q(n15535) );
  nnd2s1 U16061 ( .DIN1(n13440), .DIN2(n15546), .Q(n15545) );
  nnd3s1 U16062 ( .DIN1(n13805), .DIN2(n13957), .DIN3(n14251), .Q(n15546) );
  nnd2s1 U16063 ( .DIN1(n13431), .DIN2(n15547), .Q(n15544) );
  nnd2s1 U16064 ( .DIN1(n14257), .DIN2(n13674), .Q(n15547) );
  nnd2s1 U16065 ( .DIN1(n13765), .DIN2(n15528), .Q(n15543) );
  nnd2s1 U16066 ( .DIN1(n13667), .DIN2(n13664), .Q(n15528) );
  nor2s1 U16067 ( .DIN1(n13442), .DIN2(n13664), .Q(n15534) );
  and2s1 U16068 ( .DIN1(n13446), .DIN2(n15548), .Q(n15533) );
  nnd4s1 U16069 ( .DIN1(n13680), .DIN2(n13438), .DIN3(n13444), .DIN4(n13681), 
        .Q(n15548) );
  nnd2s1 U16070 ( .DIN1(n15549), .DIN2(n15550), .Q(n13444) );
  nnd3s1 U16071 ( .DIN1(n15551), .DIN2(n15552), .DIN3(n15553), .Q(n15493) );
  nnd2s1 U16072 ( .DIN1(n13799), .DIN2(n13456), .Q(n15553) );
  hi1s1 U16073 ( .DIN(n13442), .Q(n13456) );
  hi1s1 U16074 ( .DIN(n13680), .Q(n13799) );
  nnd2s1 U16075 ( .DIN1(n15554), .DIN2(n15512), .Q(n13680) );
  nnd2s1 U16076 ( .DIN1(n13446), .DIN2(n13954), .Q(n15552) );
  nnd2s1 U16077 ( .DIN1(n14311), .DIN2(n13950), .Q(n15551) );
  hi1s1 U16078 ( .DIN(n14004), .Q(n13950) );
  nnd2s1 U16079 ( .DIN1(n15555), .DIN2(n15556), .Q(n14004) );
  hi1s1 U16080 ( .DIN(n13677), .Q(n14311) );
  nnd4s1 U16081 ( .DIN1(n15557), .DIN2(n15558), .DIN3(n15559), .DIN4(n15560), 
        .Q(n15492) );
  nnd2s1 U16082 ( .DIN1(n13457), .DIN2(n15561), .Q(n15560) );
  nnd2s1 U16083 ( .DIN1(n14232), .DIN2(n13443), .Q(n15561) );
  nnd3s1 U16084 ( .DIN1(n15556), .DIN2(n1378), .DIN3(sa31[1]), .Q(n14232) );
  nnd2s1 U16085 ( .DIN1(n13430), .DIN2(n15562), .Q(n15559) );
  nnd4s1 U16086 ( .DIN1(n13443), .DIN2(n13957), .DIN3(n14323), .DIN4(n13786), 
        .Q(n15562) );
  nnd3s1 U16087 ( .DIN1(n1379), .DIN2(n1421), .DIN3(n15563), .Q(n13443) );
  hi1s1 U16088 ( .DIN(n13681), .Q(n13430) );
  nnd2s1 U16089 ( .DIN1(n15554), .DIN2(n15542), .Q(n13681) );
  nnd2s1 U16090 ( .DIN1(n13426), .DIN2(n14273), .Q(n15558) );
  nnd2s1 U16091 ( .DIN1(n14234), .DIN2(n13667), .Q(n14273) );
  hi1s1 U16092 ( .DIN(n13949), .Q(n13426) );
  nnd2s1 U16093 ( .DIN1(n13660), .DIN2(n13958), .Q(n15557) );
  nnd2s1 U16094 ( .DIN1(n13677), .DIN2(n13664), .Q(n13958) );
  nnd2s1 U16095 ( .DIN1(n15554), .DIN2(n15564), .Q(n13677) );
  hi1s1 U16096 ( .DIN(n14003), .Q(n13660) );
  nnd2s1 U16097 ( .DIN1(n13766), .DIN2(n13777), .Q(n15450) );
  hi1s1 U16098 ( .DIN(n13438), .Q(n13777) );
  nnd2s1 U16099 ( .DIN1(n15550), .DIN2(n15512), .Q(n13438) );
  and2s1 U16100 ( .DIN1(sa31[7]), .DIN2(sa31[6]), .Q(n15512) );
  hi1s1 U16101 ( .DIN(n13956), .Q(n13766) );
  nnd2s1 U16102 ( .DIN1(n13778), .DIN2(n13969), .Q(n15449) );
  hi1s1 U16103 ( .DIN(n13793), .Q(n13969) );
  nnd2s1 U16104 ( .DIN1(n15564), .DIN2(n15550), .Q(n13793) );
  hi1s1 U16105 ( .DIN(n13805), .Q(n13778) );
  nnd2s1 U16106 ( .DIN1(n15565), .DIN2(n15556), .Q(n13805) );
  nnd3s1 U16107 ( .DIN1(n14015), .DIN2(n15566), .DIN3(n15567), .Q(n15447) );
  nnd2s1 U16108 ( .DIN1(n13787), .DIN2(n13968), .Q(n15567) );
  hi1s1 U16109 ( .DIN(n13667), .Q(n13968) );
  nnd2s1 U16110 ( .DIN1(n15549), .DIN2(n15541), .Q(n13667) );
  hi1s1 U16111 ( .DIN(n13806), .Q(n13787) );
  nnd3s1 U16112 ( .DIN1(n1379), .DIN2(n1418), .DIN3(n15555), .Q(n13806) );
  nnd2s1 U16113 ( .DIN1(n13446), .DIN2(n13429), .Q(n15566) );
  hi1s1 U16114 ( .DIN(n14277), .Q(n13429) );
  nnd2s1 U16115 ( .DIN1(n15511), .DIN2(n15542), .Q(n14277) );
  hi1s1 U16116 ( .DIN(n13791), .Q(n13446) );
  nnd2s1 U16117 ( .DIN1(n15568), .DIN2(n15555), .Q(n13791) );
  nnd2s1 U16118 ( .DIN1(n13776), .DIN2(n13431), .Q(n14015) );
  hi1s1 U16119 ( .DIN(n14237), .Q(n13431) );
  nnd3s1 U16120 ( .DIN1(sa31[0]), .DIN2(n1418), .DIN3(n15565), .Q(n14237) );
  hi1s1 U16121 ( .DIN(n13664), .Q(n13776) );
  nnd2s1 U16122 ( .DIN1(n15542), .DIN2(n15550), .Q(n13664) );
  nor2s1 U16123 ( .DIN1(n1511), .DIN2(n1408), .Q(n15550) );
  nor2s1 U16124 ( .DIN1(sa31[7]), .DIN2(sa31[6]), .Q(n15542) );
  nnd4s1 U16125 ( .DIN1(n15569), .DIN2(n15570), .DIN3(n15571), .DIN4(n15572), 
        .Q(n15446) );
  nnd2s1 U16126 ( .DIN1(n13954), .DIN2(n15573), .Q(n15572) );
  nnd2s1 U16127 ( .DIN1(n13949), .DIN2(n14323), .Q(n15573) );
  nnd3s1 U16128 ( .DIN1(n1421), .DIN2(n1378), .DIN3(n15556), .Q(n14323) );
  nor2s1 U16129 ( .DIN1(n1418), .DIN2(n1379), .Q(n15556) );
  nnd3s1 U16130 ( .DIN1(n1421), .DIN2(n1378), .DIN3(n15568), .Q(n13949) );
  hi1s1 U16131 ( .DIN(n13673), .Q(n13954) );
  nnd2s1 U16132 ( .DIN1(n15564), .DIN2(n15511), .Q(n13673) );
  nnd2s1 U16133 ( .DIN1(n13457), .DIN2(n15574), .Q(n15571) );
  nnd2s1 U16134 ( .DIN1(n13785), .DIN2(n13442), .Q(n15574) );
  nnd2s1 U16135 ( .DIN1(n15568), .DIN2(n15565), .Q(n13442) );
  hi1s1 U16136 ( .DIN(n14257), .Q(n13457) );
  nnd2s1 U16137 ( .DIN1(n15549), .DIN2(n15511), .Q(n14257) );
  nor2s1 U16138 ( .DIN1(n1511), .DIN2(sa31[5]), .Q(n15511) );
  nnd2s1 U16139 ( .DIN1(n13440), .DIN2(n15575), .Q(n15570) );
  or2s1 U16140 ( .DIN1(n13676), .DIN2(n13765), .Q(n15575) );
  nnd2s1 U16141 ( .DIN1(n13785), .DIN2(n13956), .Q(n13676) );
  nnd3s1 U16142 ( .DIN1(sa31[1]), .DIN2(n1378), .DIN3(n15568), .Q(n13956) );
  nor2s1 U16143 ( .DIN1(n1418), .DIN2(sa31[0]), .Q(n15568) );
  nnd3s1 U16144 ( .DIN1(n1379), .DIN2(n1418), .DIN3(n15565), .Q(n13785) );
  nor2s1 U16145 ( .DIN1(n1378), .DIN2(sa31[1]), .Q(n15565) );
  hi1s1 U16146 ( .DIN(n14234), .Q(n13440) );
  nnd2s1 U16147 ( .DIN1(n15554), .DIN2(n15549), .Q(n14234) );
  and2s1 U16148 ( .DIN1(sa31[6]), .DIN2(n1539), .Q(n15549) );
  nor2s1 U16149 ( .DIN1(sa31[5]), .DIN2(sa31[4]), .Q(n15554) );
  nnd2s1 U16150 ( .DIN1(n13424), .DIN2(n15576), .Q(n15569) );
  nnd3s1 U16151 ( .DIN1(n14003), .DIN2(n13957), .DIN3(n13665), .Q(n15576) );
  nor2s1 U16152 ( .DIN1(n13765), .DIN2(n13807), .Q(n13665) );
  hi1s1 U16153 ( .DIN(n14251), .Q(n13807) );
  nnd3s1 U16154 ( .DIN1(sa31[0]), .DIN2(n1421), .DIN3(n15563), .Q(n14251) );
  hi1s1 U16155 ( .DIN(n13786), .Q(n13765) );
  nnd3s1 U16156 ( .DIN1(sa31[1]), .DIN2(sa31[0]), .DIN3(n15563), .Q(n13786) );
  nnd3s1 U16157 ( .DIN1(sa31[0]), .DIN2(n1418), .DIN3(n15555), .Q(n13957) );
  nor2s1 U16158 ( .DIN1(n1378), .DIN2(n1421), .Q(n15555) );
  nnd3s1 U16159 ( .DIN1(sa31[1]), .DIN2(n1379), .DIN3(n15563), .Q(n14003) );
  nor2s1 U16160 ( .DIN1(sa31[3]), .DIN2(sa31[2]), .Q(n15563) );
  hi1s1 U16161 ( .DIN(n13674), .Q(n13424) );
  nnd2s1 U16162 ( .DIN1(n15564), .DIN2(n15541), .Q(n13674) );
  nor2s1 U16163 ( .DIN1(n1408), .DIN2(sa31[4]), .Q(n15541) );
  nor2s1 U16164 ( .DIN1(n1539), .DIN2(sa31[6]), .Q(n15564) );
endmodule

