
module dlx ( clk, \DM_read_data[31] , \DM_read_data[30] , 
        \DM_read_data[29] , \DM_read_data[28] , \DM_read_data[27] , 
        \DM_read_data[26] , \DM_read_data[25] , \DM_read_data[24] , 
        \DM_read_data[23] , \DM_read_data[22] , \DM_read_data[21] , 
        \DM_read_data[20] , \DM_read_data[19] , \DM_read_data[18] , 
        \DM_read_data[17] , \DM_read_data[16] , \DM_read_data[15] , 
        \DM_read_data[14] , \DM_read_data[13] , \DM_read_data[12] , 
        \DM_read_data[11] , \DM_read_data[10] , \DM_read_data[9] , 
        \DM_read_data[8] , \DM_read_data[7] , \DM_read_data[6] , 
        \DM_read_data[5] , \DM_read_data[4] , \DM_read_data[3] , 
        \DM_read_data[2] , \DM_read_data[1] , \DM_read_data[0] , 
        \DM_write_data[31] , \DM_write_data[30] , \DM_write_data[29] , 
        \DM_write_data[28] , \DM_write_data[27] , \DM_write_data[26] , 
        \DM_write_data[25] , \DM_write_data[24] , \DM_write_data[23] , 
        \DM_write_data[22] , \DM_write_data[21] , \DM_write_data[20] , 
        \DM_write_data[19] , \DM_write_data[18] , \DM_write_data[17] , 
        \DM_write_data[16] , \DM_write_data[15] , \DM_write_data[14] , 
        \DM_write_data[13] , \DM_write_data[12] , \DM_write_data[11] , 
        \DM_write_data[10] , \DM_write_data[9] , \DM_write_data[8] , 
        \DM_write_data[7] , \DM_write_data[6] , \DM_write_data[5] , 
        \DM_write_data[4] , \DM_write_data[3] , \DM_write_data[2] , 
        \DM_write_data[1] , \DM_write_data[0] , \DM_addr[31] , \DM_addr[30] , 
        \DM_addr[29] , \DM_addr[28] , \DM_addr[27] , \DM_addr[26] , 
        \DM_addr[25] , \DM_addr[24] , \DM_addr[23] , \DM_addr[22] , 
        \DM_addr[21] , \DM_addr[20] , \DM_addr[19] , \DM_addr[18] , 
        \DM_addr[17] , \DM_addr[16] , \DM_addr[15] , \DM_addr[14] , 
        \DM_addr[13] , \DM_addr[12] , \DM_addr[11] , \DM_addr[10] , 
        \DM_addr[9] , \DM_addr[8] , \DM_addr[7] , \DM_addr[6] , \DM_addr[5] , 
        \DM_addr[4] , \DM_addr[3] , \DM_addr[2] , \DM_addr[1] , \DM_addr[0] , 
        DM_write, DM_read, \NPC[31] , \NPC[30] , \NPC[29] , \NPC[28] , 
        \NPC[27] , \NPC[26] , \NPC[25] , \NPC[24] , \NPC[23] , \NPC[22] , 
        \NPC[21] , \NPC[20] , \NPC[19] , \NPC[18] , \NPC[17] , \NPC[16] , 
        \NPC[15] , \NPC[14] , \NPC[13] , \NPC[12] , \NPC[11] , \NPC[10] , 
        \NPC[9] , \NPC[8] , \NPC[7] , \NPC[6] , \NPC[5] , \NPC[4] , \NPC[3] , 
        \NPC[2] , \NPC[1] , \NPC[0] , reset, \IR[31] , \IR[30] , \IR[29] , 
        \IR[28] , \IR[27] , \IR[26] , \IR[25] , \IR[24] , \IR[23] , \IR[22] , 
        \IR[21] , \IR[20] , \IR[19] , \IR[18] , \IR[17] , \IR[16] , \IR[15] , 
        \IR[14] , \IR[13] , \IR[12] , \IR[11] , \IR[10] , \IR[9] , \IR[8] , 
        \IR[7] , \IR[6] , \IR[5] , \IR[4] , \IR[3] , \IR[2] , \IR[1] , \IR[0] , 
        byte, word, INT, CLI, PIPEEMPTY, FREEZE );
  input clk, \DM_read_data[31] , \DM_read_data[30] , \DM_read_data[29] ,
         \DM_read_data[28] , \DM_read_data[27] , \DM_read_data[26] ,
         \DM_read_data[25] , \DM_read_data[24] , \DM_read_data[23] ,
         \DM_read_data[22] , \DM_read_data[21] , \DM_read_data[20] ,
         \DM_read_data[19] , \DM_read_data[18] , \DM_read_data[17] ,
         \DM_read_data[16] , \DM_read_data[15] , \DM_read_data[14] ,
         \DM_read_data[13] , \DM_read_data[12] , \DM_read_data[11] ,
         \DM_read_data[10] , \DM_read_data[9] , \DM_read_data[8] ,
         \DM_read_data[7] , \DM_read_data[6] , \DM_read_data[5] ,
         \DM_read_data[4] , \DM_read_data[3] , \DM_read_data[2] ,
         \DM_read_data[1] , \DM_read_data[0] , reset, \IR[31] , \IR[30] ,
         \IR[29] , \IR[28] , \IR[27] , \IR[26] , \IR[25] , \IR[24] , \IR[23] ,
         \IR[22] , \IR[21] , \IR[20] , \IR[19] , \IR[18] , \IR[17] , \IR[16] ,
         \IR[15] , \IR[14] , \IR[13] , \IR[12] , \IR[11] , \IR[10] , \IR[9] ,
         \IR[8] , \IR[7] , \IR[6] , \IR[5] , \IR[4] , \IR[3] , \IR[2] ,
         \IR[1] , \IR[0] , INT, FREEZE;
  output \DM_write_data[31] , \DM_write_data[30] , \DM_write_data[29] ,
         \DM_write_data[28] , \DM_write_data[27] , \DM_write_data[26] ,
         \DM_write_data[25] , \DM_write_data[24] , \DM_write_data[23] ,
         \DM_write_data[22] , \DM_write_data[21] , \DM_write_data[20] ,
         \DM_write_data[19] , \DM_write_data[18] , \DM_write_data[17] ,
         \DM_write_data[16] , \DM_write_data[15] , \DM_write_data[14] ,
         \DM_write_data[13] , \DM_write_data[12] , \DM_write_data[11] ,
         \DM_write_data[10] , \DM_write_data[9] , \DM_write_data[8] ,
         \DM_write_data[7] , \DM_write_data[6] , \DM_write_data[5] ,
         \DM_write_data[4] , \DM_write_data[3] , \DM_write_data[2] ,
         \DM_write_data[1] , \DM_write_data[0] , \DM_addr[31] , \DM_addr[30] ,
         \DM_addr[29] , \DM_addr[28] , \DM_addr[27] , \DM_addr[26] ,
         \DM_addr[25] , \DM_addr[24] , \DM_addr[23] , \DM_addr[22] ,
         \DM_addr[21] , \DM_addr[20] , \DM_addr[19] , \DM_addr[18] ,
         \DM_addr[17] , \DM_addr[16] , \DM_addr[15] , \DM_addr[14] ,
         \DM_addr[13] , \DM_addr[12] , \DM_addr[11] , \DM_addr[10] ,
         \DM_addr[9] , \DM_addr[8] , \DM_addr[7] , \DM_addr[6] , \DM_addr[5] ,
         \DM_addr[4] , \DM_addr[3] , \DM_addr[2] , \DM_addr[1] , \DM_addr[0] ,
         DM_write, DM_read, \NPC[31] , \NPC[30] , \NPC[29] , \NPC[28] ,
         \NPC[27] , \NPC[26] , \NPC[25] , \NPC[24] , \NPC[23] , \NPC[22] ,
         \NPC[21] , \NPC[20] , \NPC[19] , \NPC[18] , \NPC[17] , \NPC[16] ,
         \NPC[15] , \NPC[14] , \NPC[13] , \NPC[12] , \NPC[11] , \NPC[10] ,
         \NPC[9] , \NPC[8] , \NPC[7] , \NPC[6] , \NPC[5] , \NPC[4] , \NPC[3] ,
         \NPC[2] , \NPC[1] , \NPC[0] , byte, word, CLI, PIPEEMPTY;
  wire   stall, reg_dst, reg_write, reg_write_MEM, reg_write_EX, \IFinst/n848 ,
         \IFinst/n847 , \IFinst/n846 , \IFinst/n845 , \IFinst/n844 ,
         \IFinst/n843 , \IFinst/n842 , \IFinst/n841 , \IFinst/n840 ,
         \IFinst/n839 , \IFinst/n838 , \IFinst/n837 , \IFinst/n836 ,
         \IFinst/n835 , \IFinst/n834 , \IFinst/n833 , \IFinst/n832 ,
         \IFinst/n831 , \IFinst/n830 , \IFinst/n829 , \IFinst/n828 ,
         \IFinst/n827 , \IFinst/n826 , \IFinst/n825 , \IFinst/n824 ,
         \IFinst/n823 , \IFinst/n822 , \IFinst/n821 , \IFinst/n820 ,
         \IFinst/n819 , \IFinst/n818 , \IFinst/n817 , \IFinst/n816 ,
         \IFinst/n749 , \IFinst/n746 , \IFinst/n744 , \IFinst/n741 ,
         \IFinst/n739 , \IFinst/n736 , \IFinst/n734 , \IFinst/n731 ,
         \IFinst/n729 , \IFinst/n726 , \IFinst/n724 , \IFinst/n721 ,
         \IFinst/n719 , \IFinst/n716 , \IFinst/n714 , \IFinst/n711 ,
         \IFinst/n709 , \IFinst/n706 , \IFinst/n704 , \IFinst/n701 ,
         \IFinst/n699 , \IFinst/n696 , \IFinst/n694 , \IFinst/n691 ,
         \IFinst/n689 , \IFinst/n686 , \IFinst/n684 , \IFinst/n681 ,
         \IFinst/n679 , \IFinst/n676 , \IFinst/n674 , \IFinst/n671 ,
         \IFinst/n669 , \IFinst/n666 , \IFinst/n664 , \IFinst/n661 ,
         \IFinst/n659 , \IFinst/n656 , \IFinst/n654 , \IFinst/n651 ,
         \IFinst/n649 , \IFinst/n646 , \IFinst/n644 , \IFinst/n641 ,
         \IFinst/n639 , \IFinst/n636 , \IFinst/n634 , \IFinst/n631 ,
         \IFinst/n629 , \IFinst/n626 , \IFinst/n624 , \IFinst/n621 ,
         \IFinst/n619 , \IFinst/n616 , \IFinst/n614 , \IFinst/n611 ,
         \IFinst/n609 , \IFinst/n606 , \IFinst/n604 , \IFinst/n601 ,
         \IFinst/n599 , \IFinst/n596 , \IFinst/n594 , \IFinst/n591 ,
         \IFinst/N135 , \IFinst/N134 , \IFinst/N133 , \IFinst/N132 ,
         \IFinst/N131 , \IFinst/N130 , \IFinst/N129 , \IFinst/N128 ,
         \IFinst/N127 , \IFinst/N126 , \IFinst/N125 , \IFinst/N124 ,
         \IFinst/N123 , \IFinst/N122 , \IFinst/N121 , \IFinst/N120 ,
         \IFinst/N119 , \IFinst/N118 , \IFinst/N117 , \IFinst/N116 ,
         \IFinst/N115 , \IFinst/N114 , \IFinst/N113 , \IFinst/N112 ,
         \IFinst/N111 , \IFinst/N110 , \IFinst/N109 , \IFinst/N108 ,
         \IFinst/N107 , \IFinst/N106 , \IFinst/N105 , \IFinst/N104 ,
         \IFinst/N103 , \IFinst/N102 , \IFinst/N101 , \IFinst/N100 ,
         \IFinst/N99 , \IFinst/N98 , \IFinst/N97 , \IFinst/N96 , \IFinst/N95 ,
         \IFinst/N94 , \IFinst/N93 , \IFinst/N92 , \IFinst/N91 , \IFinst/N90 ,
         \IFinst/N89 , \IFinst/N88 , \IFinst/N87 , \IFinst/N86 , \IFinst/N85 ,
         \IFinst/N84 , \IFinst/N83 , \IFinst/N82 , \IFinst/N81 , \IFinst/N80 ,
         \IFinst/N79 , \IFinst/N78 , \IFinst/N77 , \IFinst/N76 , \IFinst/N75 ,
         \IFinst/N74 , \IFinst/N73 , \IFinst/N72 , \IFinst/N8 , \IFinst/N7 ,
         \IDinst/n11835 , \IDinst/n11834 , \IDinst/n11833 , \IDinst/n11832 ,
         \IDinst/n11831 , \IDinst/n11830 , \IDinst/n11829 , \IDinst/n11828 ,
         \IDinst/n11827 , \IDinst/n11826 , \IDinst/n11825 , \IDinst/n11824 ,
         \IDinst/n11823 , \IDinst/n11822 , \IDinst/n11821 , \IDinst/n11820 ,
         \IDinst/n11819 , \IDinst/n11818 , \IDinst/n11817 , \IDinst/n11816 ,
         \IDinst/n11815 , \IDinst/n11814 , \IDinst/n11813 , \IDinst/n11812 ,
         \IDinst/n11811 , \IDinst/n11810 , \IDinst/n11809 , \IDinst/n11808 ,
         \IDinst/n11807 , \IDinst/n11806 , \IDinst/n11805 , \IDinst/n11804 ,
         \IDinst/n11803 , \IDinst/n11802 , \IDinst/n11801 , \IDinst/n11800 ,
         \IDinst/n11799 , \IDinst/n11798 , \IDinst/n11797 , \IDinst/n11796 ,
         \IDinst/n11795 , \IDinst/n11794 , \IDinst/n11793 , \IDinst/n11792 ,
         \IDinst/n11791 , \IDinst/n11790 , \IDinst/n11789 , \IDinst/n11788 ,
         \IDinst/n11787 , \IDinst/n11786 , \IDinst/n11785 , \IDinst/n11784 ,
         \IDinst/n11783 , \IDinst/n11782 , \IDinst/n11781 , \IDinst/n11780 ,
         \IDinst/n11779 , \IDinst/n11778 , \IDinst/n11777 , \IDinst/n11776 ,
         \IDinst/n11775 , \IDinst/n11774 , \IDinst/n11773 , \IDinst/n11772 ,
         \IDinst/n11771 , \IDinst/n11770 , \IDinst/n11769 , \IDinst/n11768 ,
         \IDinst/n11767 , \IDinst/n11766 , \IDinst/n11765 , \IDinst/n11764 ,
         \IDinst/n11763 , \IDinst/n11762 , \IDinst/n11761 , \IDinst/n11760 ,
         \IDinst/n11759 , \IDinst/n11758 , \IDinst/n11757 , \IDinst/n11756 ,
         \IDinst/n11755 , \IDinst/n11754 , \IDinst/n11753 , \IDinst/n11752 ,
         \IDinst/n11751 , \IDinst/n11750 , \IDinst/n11749 , \IDinst/n11748 ,
         \IDinst/n11747 , \IDinst/n11746 , \IDinst/n11745 , \IDinst/n11744 ,
         \IDinst/n11743 , \IDinst/n11742 , \IDinst/n11741 , \IDinst/n11740 ,
         \IDinst/n11739 , \IDinst/n11738 , \IDinst/n11737 , \IDinst/n11736 ,
         \IDinst/n11735 , \IDinst/n11734 , \IDinst/n11733 , \IDinst/n11732 ,
         \IDinst/n11731 , \IDinst/n11730 , \IDinst/n11729 , \IDinst/n11728 ,
         \IDinst/n11727 , \IDinst/n11726 , \IDinst/n11725 , \IDinst/n11724 ,
         \IDinst/n11723 , \IDinst/n11722 , \IDinst/n11721 , \IDinst/n11720 ,
         \IDinst/n11719 , \IDinst/n11718 , \IDinst/n11717 , \IDinst/n11716 ,
         \IDinst/n11715 , \IDinst/n11714 , \IDinst/n11713 , \IDinst/n11712 ,
         \IDinst/n11711 , \IDinst/n11710 , \IDinst/n11709 , \IDinst/n11708 ,
         \IDinst/n11707 , \IDinst/n11706 , \IDinst/n11705 , \IDinst/n11704 ,
         \IDinst/n11703 , \IDinst/n11702 , \IDinst/n11701 , \IDinst/n11700 ,
         \IDinst/n11699 , \IDinst/n11698 , \IDinst/n11697 , \IDinst/n11696 ,
         \IDinst/n11695 , \IDinst/n11694 , \IDinst/n11693 , \IDinst/n11692 ,
         \IDinst/n11691 , \IDinst/n11690 , \IDinst/n11689 , \IDinst/n11688 ,
         \IDinst/n11687 , \IDinst/n11686 , \IDinst/n11685 , \IDinst/n11684 ,
         \IDinst/n11683 , \IDinst/n11682 , \IDinst/n11681 , \IDinst/n11680 ,
         \IDinst/n11679 , \IDinst/n11678 , \IDinst/n11677 , \IDinst/n11676 ,
         \IDinst/n11675 , \IDinst/n11674 , \IDinst/n11673 , \IDinst/n11672 ,
         \IDinst/n11671 , \IDinst/n11670 , \IDinst/n11669 , \IDinst/n11668 ,
         \IDinst/n11667 , \IDinst/n11666 , \IDinst/n11665 , \IDinst/n11664 ,
         \IDinst/n11663 , \IDinst/n11662 , \IDinst/n11661 , \IDinst/n11660 ,
         \IDinst/n11659 , \IDinst/n11658 , \IDinst/n11657 , \IDinst/n11656 ,
         \IDinst/n11655 , \IDinst/n11654 , \IDinst/n11653 , \IDinst/n11652 ,
         \IDinst/n11651 , \IDinst/n11650 , \IDinst/n11649 , \IDinst/n11648 ,
         \IDinst/n11647 , \IDinst/n11646 , \IDinst/n11645 , \IDinst/n11644 ,
         \IDinst/n11643 , \IDinst/n11642 , \IDinst/n11641 , \IDinst/n11640 ,
         \IDinst/n11639 , \IDinst/n11638 , \IDinst/n11637 , \IDinst/n11636 ,
         \IDinst/n11635 , \IDinst/n11634 , \IDinst/n11633 , \IDinst/n11632 ,
         \IDinst/n11631 , \IDinst/n11630 , \IDinst/n11629 , \IDinst/n11628 ,
         \IDinst/n11627 , \IDinst/n11626 , \IDinst/n11625 , \IDinst/n11624 ,
         \IDinst/n11623 , \IDinst/n11622 , \IDinst/n11621 , \IDinst/n11620 ,
         \IDinst/n11619 , \IDinst/n11618 , \IDinst/n11617 , \IDinst/n11616 ,
         \IDinst/n11615 , \IDinst/n11614 , \IDinst/n11613 , \IDinst/n11612 ,
         \IDinst/n11611 , \IDinst/n11610 , \IDinst/n11609 , \IDinst/n11608 ,
         \IDinst/n11607 , \IDinst/n11606 , \IDinst/n11605 , \IDinst/n11604 ,
         \IDinst/n11603 , \IDinst/n11602 , \IDinst/n11601 , \IDinst/n11600 ,
         \IDinst/n11599 , \IDinst/n11598 , \IDinst/n11597 , \IDinst/n11596 ,
         \IDinst/n11595 , \IDinst/n11594 , \IDinst/n11593 , \IDinst/n11592 ,
         \IDinst/n11591 , \IDinst/n11590 , \IDinst/n11589 , \IDinst/n11588 ,
         \IDinst/n11587 , \IDinst/n11586 , \IDinst/n11585 , \IDinst/n11584 ,
         \IDinst/n11583 , \IDinst/n11582 , \IDinst/n11581 , \IDinst/n11580 ,
         \IDinst/n11579 , \IDinst/n11578 , \IDinst/n11577 , \IDinst/n11576 ,
         \IDinst/n11575 , \IDinst/n11574 , \IDinst/n11573 , \IDinst/n11572 ,
         \IDinst/n11571 , \IDinst/n11570 , \IDinst/n11569 , \IDinst/n11568 ,
         \IDinst/n11567 , \IDinst/n11566 , \IDinst/n11565 , \IDinst/n11564 ,
         \IDinst/n11563 , \IDinst/n11562 , \IDinst/n11561 , \IDinst/n11560 ,
         \IDinst/n11559 , \IDinst/n11558 , \IDinst/n11557 , \IDinst/n11556 ,
         \IDinst/n11555 , \IDinst/n11554 , \IDinst/n11553 , \IDinst/n11552 ,
         \IDinst/n11551 , \IDinst/n11550 , \IDinst/n11549 , \IDinst/n11548 ,
         \IDinst/n11547 , \IDinst/n11546 , \IDinst/n11545 , \IDinst/n11544 ,
         \IDinst/n11543 , \IDinst/n11542 , \IDinst/n11541 , \IDinst/n11540 ,
         \IDinst/n11539 , \IDinst/n11538 , \IDinst/n11537 , \IDinst/n11536 ,
         \IDinst/n11535 , \IDinst/n11534 , \IDinst/n11533 , \IDinst/n11532 ,
         \IDinst/n11531 , \IDinst/n11530 , \IDinst/n11529 , \IDinst/n11528 ,
         \IDinst/n11527 , \IDinst/n11526 , \IDinst/n11525 , \IDinst/n11524 ,
         \IDinst/n11523 , \IDinst/n11522 , \IDinst/n11521 , \IDinst/n11520 ,
         \IDinst/n11519 , \IDinst/n11518 , \IDinst/n11517 , \IDinst/n11516 ,
         \IDinst/n11515 , \IDinst/n11514 , \IDinst/n11513 , \IDinst/n11512 ,
         \IDinst/n11511 , \IDinst/n11510 , \IDinst/n11509 , \IDinst/n11508 ,
         \IDinst/n11507 , \IDinst/n11506 , \IDinst/n11505 , \IDinst/n11504 ,
         \IDinst/n11503 , \IDinst/n11502 , \IDinst/n11501 , \IDinst/n11500 ,
         \IDinst/n11499 , \IDinst/n11498 , \IDinst/n11497 , \IDinst/n11496 ,
         \IDinst/n11495 , \IDinst/n11494 , \IDinst/n11493 , \IDinst/n11492 ,
         \IDinst/n11491 , \IDinst/n11490 , \IDinst/n11489 , \IDinst/n11488 ,
         \IDinst/n11487 , \IDinst/n11486 , \IDinst/n11485 , \IDinst/n11484 ,
         \IDinst/n11483 , \IDinst/n11482 , \IDinst/n11481 , \IDinst/n11480 ,
         \IDinst/n11479 , \IDinst/n11478 , \IDinst/n11477 , \IDinst/n11476 ,
         \IDinst/n11475 , \IDinst/n11474 , \IDinst/n11473 , \IDinst/n11472 ,
         \IDinst/n11471 , \IDinst/n11470 , \IDinst/n11469 , \IDinst/n11468 ,
         \IDinst/n11467 , \IDinst/n11466 , \IDinst/n11465 , \IDinst/n11464 ,
         \IDinst/n11463 , \IDinst/n11462 , \IDinst/n11461 , \IDinst/n11460 ,
         \IDinst/n11459 , \IDinst/n11458 , \IDinst/n11457 , \IDinst/n11456 ,
         \IDinst/n11455 , \IDinst/n11454 , \IDinst/n11453 , \IDinst/n11452 ,
         \IDinst/n11451 , \IDinst/n11450 , \IDinst/n11449 , \IDinst/n11448 ,
         \IDinst/n11447 , \IDinst/n11446 , \IDinst/n11445 , \IDinst/n11444 ,
         \IDinst/n11443 , \IDinst/n11442 , \IDinst/n11441 , \IDinst/n11440 ,
         \IDinst/n11439 , \IDinst/n11438 , \IDinst/n11437 , \IDinst/n11436 ,
         \IDinst/n11435 , \IDinst/n11434 , \IDinst/n11433 , \IDinst/n11432 ,
         \IDinst/n11431 , \IDinst/n11430 , \IDinst/n11429 , \IDinst/n11428 ,
         \IDinst/n11427 , \IDinst/n11426 , \IDinst/n11425 , \IDinst/n11424 ,
         \IDinst/n11423 , \IDinst/n11422 , \IDinst/n11421 , \IDinst/n11420 ,
         \IDinst/n11419 , \IDinst/n11418 , \IDinst/n11417 , \IDinst/n11416 ,
         \IDinst/n11415 , \IDinst/n11414 , \IDinst/n11413 , \IDinst/n11412 ,
         \IDinst/n11411 , \IDinst/n11410 , \IDinst/n11409 , \IDinst/n11408 ,
         \IDinst/n11407 , \IDinst/n11406 , \IDinst/n11405 , \IDinst/n11404 ,
         \IDinst/n11403 , \IDinst/n11402 , \IDinst/n11401 , \IDinst/n11400 ,
         \IDinst/n11399 , \IDinst/n11398 , \IDinst/n11397 , \IDinst/n11396 ,
         \IDinst/n11395 , \IDinst/n11394 , \IDinst/n11393 , \IDinst/n11392 ,
         \IDinst/n11391 , \IDinst/n11390 , \IDinst/n11389 , \IDinst/n11388 ,
         \IDinst/n11387 , \IDinst/n11386 , \IDinst/n11385 , \IDinst/n11384 ,
         \IDinst/n11383 , \IDinst/n11382 , \IDinst/n11381 , \IDinst/n11380 ,
         \IDinst/n11379 , \IDinst/n11378 , \IDinst/n11377 , \IDinst/n11376 ,
         \IDinst/n11375 , \IDinst/n11374 , \IDinst/n11373 , \IDinst/n11372 ,
         \IDinst/n11371 , \IDinst/n11370 , \IDinst/n11369 , \IDinst/n11368 ,
         \IDinst/n11367 , \IDinst/n11366 , \IDinst/n11365 , \IDinst/n11364 ,
         \IDinst/n11363 , \IDinst/n11362 , \IDinst/n11361 , \IDinst/n11360 ,
         \IDinst/n11359 , \IDinst/n11358 , \IDinst/n11357 , \IDinst/n11356 ,
         \IDinst/n11355 , \IDinst/n11354 , \IDinst/n11353 , \IDinst/n11352 ,
         \IDinst/n11351 , \IDinst/n11350 , \IDinst/n11349 , \IDinst/n11348 ,
         \IDinst/n11347 , \IDinst/n11346 , \IDinst/n11345 , \IDinst/n11344 ,
         \IDinst/n11343 , \IDinst/n11342 , \IDinst/n11341 , \IDinst/n11340 ,
         \IDinst/n11339 , \IDinst/n11338 , \IDinst/n11337 , \IDinst/n11336 ,
         \IDinst/n11335 , \IDinst/n11334 , \IDinst/n11333 , \IDinst/n11332 ,
         \IDinst/n11331 , \IDinst/n11330 , \IDinst/n11329 , \IDinst/n11328 ,
         \IDinst/n11327 , \IDinst/n11326 , \IDinst/n11325 , \IDinst/n11324 ,
         \IDinst/n11323 , \IDinst/n11322 , \IDinst/n11321 , \IDinst/n11320 ,
         \IDinst/n11319 , \IDinst/n11318 , \IDinst/n11317 , \IDinst/n11316 ,
         \IDinst/n11315 , \IDinst/n11314 , \IDinst/n11313 , \IDinst/n11312 ,
         \IDinst/n11311 , \IDinst/n11310 , \IDinst/n11309 , \IDinst/n11308 ,
         \IDinst/n11307 , \IDinst/n11306 , \IDinst/n11305 , \IDinst/n11304 ,
         \IDinst/n11303 , \IDinst/n11302 , \IDinst/n11301 , \IDinst/n11300 ,
         \IDinst/n11299 , \IDinst/n11298 , \IDinst/n11297 , \IDinst/n11296 ,
         \IDinst/n11295 , \IDinst/n11294 , \IDinst/n11293 , \IDinst/n11292 ,
         \IDinst/n11291 , \IDinst/n11290 , \IDinst/n11289 , \IDinst/n11288 ,
         \IDinst/n11287 , \IDinst/n11286 , \IDinst/n11285 , \IDinst/n11284 ,
         \IDinst/n11283 , \IDinst/n11282 , \IDinst/n11281 , \IDinst/n11280 ,
         \IDinst/n11279 , \IDinst/n11278 , \IDinst/n11277 , \IDinst/n11276 ,
         \IDinst/n11275 , \IDinst/n11274 , \IDinst/n11273 , \IDinst/n11272 ,
         \IDinst/n11271 , \IDinst/n11270 , \IDinst/n11269 , \IDinst/n11268 ,
         \IDinst/n11267 , \IDinst/n11266 , \IDinst/n11265 , \IDinst/n11264 ,
         \IDinst/n11263 , \IDinst/n11262 , \IDinst/n11261 , \IDinst/n11260 ,
         \IDinst/n11259 , \IDinst/n11258 , \IDinst/n11257 , \IDinst/n11256 ,
         \IDinst/n11255 , \IDinst/n11254 , \IDinst/n11253 , \IDinst/n11252 ,
         \IDinst/n11251 , \IDinst/n11250 , \IDinst/n11249 , \IDinst/n11248 ,
         \IDinst/n11247 , \IDinst/n11246 , \IDinst/n11245 , \IDinst/n11244 ,
         \IDinst/n11243 , \IDinst/n11242 , \IDinst/n11241 , \IDinst/n11240 ,
         \IDinst/n11239 , \IDinst/n11238 , \IDinst/n11237 , \IDinst/n11236 ,
         \IDinst/n11235 , \IDinst/n11234 , \IDinst/n11233 , \IDinst/n11232 ,
         \IDinst/n11231 , \IDinst/n11230 , \IDinst/n11229 , \IDinst/n11228 ,
         \IDinst/n11227 , \IDinst/n11226 , \IDinst/n11225 , \IDinst/n11224 ,
         \IDinst/n11223 , \IDinst/n11222 , \IDinst/n11221 , \IDinst/n11220 ,
         \IDinst/n11219 , \IDinst/n11218 , \IDinst/n11217 , \IDinst/n11216 ,
         \IDinst/n11215 , \IDinst/n11214 , \IDinst/n11213 , \IDinst/n11212 ,
         \IDinst/n11211 , \IDinst/n11210 , \IDinst/n11209 , \IDinst/n11208 ,
         \IDinst/n11207 , \IDinst/n11206 , \IDinst/n11205 , \IDinst/n11204 ,
         \IDinst/n11203 , \IDinst/n11202 , \IDinst/n11201 , \IDinst/n11200 ,
         \IDinst/n11199 , \IDinst/n11198 , \IDinst/n11197 , \IDinst/n11196 ,
         \IDinst/n11195 , \IDinst/n11194 , \IDinst/n11193 , \IDinst/n11192 ,
         \IDinst/n11191 , \IDinst/n11190 , \IDinst/n11189 , \IDinst/n11188 ,
         \IDinst/n11187 , \IDinst/n11186 , \IDinst/n11185 , \IDinst/n11184 ,
         \IDinst/n11183 , \IDinst/n11182 , \IDinst/n11181 , \IDinst/n11180 ,
         \IDinst/n11179 , \IDinst/n11178 , \IDinst/n11177 , \IDinst/n11176 ,
         \IDinst/n11175 , \IDinst/n11174 , \IDinst/n11173 , \IDinst/n11172 ,
         \IDinst/n11171 , \IDinst/n11170 , \IDinst/n11169 , \IDinst/n11168 ,
         \IDinst/n11167 , \IDinst/n11166 , \IDinst/n11165 , \IDinst/n11164 ,
         \IDinst/n11163 , \IDinst/n11162 , \IDinst/n11161 , \IDinst/n11160 ,
         \IDinst/n11159 , \IDinst/n11158 , \IDinst/n11157 , \IDinst/n11156 ,
         \IDinst/n11155 , \IDinst/n11154 , \IDinst/n11153 , \IDinst/n11152 ,
         \IDinst/n11151 , \IDinst/n11150 , \IDinst/n11149 , \IDinst/n11148 ,
         \IDinst/n11147 , \IDinst/n11146 , \IDinst/n11145 , \IDinst/n11144 ,
         \IDinst/n11143 , \IDinst/n11142 , \IDinst/n11141 , \IDinst/n11140 ,
         \IDinst/n11139 , \IDinst/n11138 , \IDinst/n11137 , \IDinst/n11136 ,
         \IDinst/n11135 , \IDinst/n11134 , \IDinst/n11133 , \IDinst/n11132 ,
         \IDinst/n11131 , \IDinst/n11130 , \IDinst/n11129 , \IDinst/n11128 ,
         \IDinst/n11127 , \IDinst/n11126 , \IDinst/n11125 , \IDinst/n11124 ,
         \IDinst/n11123 , \IDinst/n11122 , \IDinst/n11121 , \IDinst/n11120 ,
         \IDinst/n11119 , \IDinst/n11118 , \IDinst/n11117 , \IDinst/n11116 ,
         \IDinst/n11115 , \IDinst/n11114 , \IDinst/n11113 , \IDinst/n11112 ,
         \IDinst/n11111 , \IDinst/n11110 , \IDinst/n11109 , \IDinst/n11108 ,
         \IDinst/n11107 , \IDinst/n11106 , \IDinst/n11105 , \IDinst/n11104 ,
         \IDinst/n11103 , \IDinst/n11102 , \IDinst/n11101 , \IDinst/n11100 ,
         \IDinst/n11099 , \IDinst/n11098 , \IDinst/n11097 , \IDinst/n11096 ,
         \IDinst/n11095 , \IDinst/n11094 , \IDinst/n11093 , \IDinst/n11092 ,
         \IDinst/n11091 , \IDinst/n11090 , \IDinst/n11089 , \IDinst/n11088 ,
         \IDinst/n11087 , \IDinst/n11086 , \IDinst/n11085 , \IDinst/n11084 ,
         \IDinst/n11083 , \IDinst/n11082 , \IDinst/n11081 , \IDinst/n11080 ,
         \IDinst/n11079 , \IDinst/n11078 , \IDinst/n11077 , \IDinst/n11076 ,
         \IDinst/n11075 , \IDinst/n11074 , \IDinst/n11073 , \IDinst/n11072 ,
         \IDinst/n11071 , \IDinst/n11070 , \IDinst/n11069 , \IDinst/n11068 ,
         \IDinst/n11067 , \IDinst/n11066 , \IDinst/n11065 , \IDinst/n11064 ,
         \IDinst/n11063 , \IDinst/n11062 , \IDinst/n11061 , \IDinst/n11060 ,
         \IDinst/n11059 , \IDinst/n11058 , \IDinst/n11057 , \IDinst/n11056 ,
         \IDinst/n11055 , \IDinst/n11054 , \IDinst/n11053 , \IDinst/n11052 ,
         \IDinst/n11051 , \IDinst/n11050 , \IDinst/n11049 , \IDinst/n11048 ,
         \IDinst/n11047 , \IDinst/n11046 , \IDinst/n11045 , \IDinst/n11044 ,
         \IDinst/n11043 , \IDinst/n11042 , \IDinst/n11041 , \IDinst/n11040 ,
         \IDinst/n11039 , \IDinst/n11038 , \IDinst/n11037 , \IDinst/n11036 ,
         \IDinst/n11035 , \IDinst/n11034 , \IDinst/n11033 , \IDinst/n11032 ,
         \IDinst/n11031 , \IDinst/n11030 , \IDinst/n11029 , \IDinst/n11028 ,
         \IDinst/n11027 , \IDinst/n11026 , \IDinst/n11025 , \IDinst/n11024 ,
         \IDinst/n11023 , \IDinst/n11022 , \IDinst/n11021 , \IDinst/n11020 ,
         \IDinst/n11019 , \IDinst/n11018 , \IDinst/n11017 , \IDinst/n11016 ,
         \IDinst/n11015 , \IDinst/n11014 , \IDinst/n11013 , \IDinst/n11012 ,
         \IDinst/n11011 , \IDinst/n11010 , \IDinst/n11009 , \IDinst/n11008 ,
         \IDinst/n11007 , \IDinst/n11006 , \IDinst/n11005 , \IDinst/n11004 ,
         \IDinst/n11003 , \IDinst/n11002 , \IDinst/n11001 , \IDinst/n11000 ,
         \IDinst/n10999 , \IDinst/n10998 , \IDinst/n10997 , \IDinst/n10996 ,
         \IDinst/n10995 , \IDinst/n10994 , \IDinst/n10993 , \IDinst/n10992 ,
         \IDinst/n10991 , \IDinst/n10990 , \IDinst/n10989 , \IDinst/n10988 ,
         \IDinst/n10987 , \IDinst/n10986 , \IDinst/n10985 , \IDinst/n10984 ,
         \IDinst/n10983 , \IDinst/n10982 , \IDinst/n10981 , \IDinst/n10980 ,
         \IDinst/n10979 , \IDinst/n10978 , \IDinst/n10977 , \IDinst/n10976 ,
         \IDinst/n10975 , \IDinst/n10974 , \IDinst/n10973 , \IDinst/n10972 ,
         \IDinst/n10971 , \IDinst/n10970 , \IDinst/n10969 , \IDinst/n10968 ,
         \IDinst/n10967 , \IDinst/n10966 , \IDinst/n10965 , \IDinst/n10964 ,
         \IDinst/n10963 , \IDinst/n10962 , \IDinst/n10961 , \IDinst/n10960 ,
         \IDinst/n10959 , \IDinst/n10958 , \IDinst/n10957 , \IDinst/n10956 ,
         \IDinst/n10955 , \IDinst/n10954 , \IDinst/n10953 , \IDinst/n10952 ,
         \IDinst/n10951 , \IDinst/n10950 , \IDinst/n10949 , \IDinst/n10948 ,
         \IDinst/n10947 , \IDinst/n10946 , \IDinst/n10945 , \IDinst/n10944 ,
         \IDinst/n10943 , \IDinst/n10942 , \IDinst/n10941 , \IDinst/n10940 ,
         \IDinst/n10939 , \IDinst/n10938 , \IDinst/n10937 , \IDinst/n10936 ,
         \IDinst/n10935 , \IDinst/n10934 , \IDinst/n10933 , \IDinst/n10932 ,
         \IDinst/n10931 , \IDinst/n10930 , \IDinst/n10929 , \IDinst/n10928 ,
         \IDinst/n10927 , \IDinst/n10926 , \IDinst/n10925 , \IDinst/n10924 ,
         \IDinst/n10923 , \IDinst/n10922 , \IDinst/n10921 , \IDinst/n10920 ,
         \IDinst/n10919 , \IDinst/n10918 , \IDinst/n10917 , \IDinst/n10916 ,
         \IDinst/n10915 , \IDinst/n10914 , \IDinst/n10913 , \IDinst/n10912 ,
         \IDinst/n10911 , \IDinst/n10910 , \IDinst/n10909 , \IDinst/n10908 ,
         \IDinst/n10907 , \IDinst/n10906 , \IDinst/n10905 , \IDinst/n10904 ,
         \IDinst/n10903 , \IDinst/n10902 , \IDinst/n10901 , \IDinst/n10900 ,
         \IDinst/n10899 , \IDinst/n10898 , \IDinst/n10897 , \IDinst/n10896 ,
         \IDinst/n10895 , \IDinst/n10894 , \IDinst/n10893 , \IDinst/n10892 ,
         \IDinst/n10891 , \IDinst/n10890 , \IDinst/n10889 , \IDinst/n10888 ,
         \IDinst/n10887 , \IDinst/n10886 , \IDinst/n10885 , \IDinst/n10884 ,
         \IDinst/n10883 , \IDinst/n10882 , \IDinst/n10881 , \IDinst/n10880 ,
         \IDinst/n10879 , \IDinst/n10878 , \IDinst/n10877 , \IDinst/n10876 ,
         \IDinst/n10875 , \IDinst/n10874 , \IDinst/n10873 , \IDinst/n10872 ,
         \IDinst/n10871 , \IDinst/n10870 , \IDinst/n10869 , \IDinst/n10868 ,
         \IDinst/n10867 , \IDinst/n10866 , \IDinst/n10865 , \IDinst/n10864 ,
         \IDinst/n10863 , \IDinst/n10862 , \IDinst/n10861 , \IDinst/n10860 ,
         \IDinst/n10859 , \IDinst/n10858 , \IDinst/n10857 , \IDinst/n10856 ,
         \IDinst/n10855 , \IDinst/n10854 , \IDinst/n10853 , \IDinst/n10852 ,
         \IDinst/n10851 , \IDinst/n10850 , \IDinst/n10849 , \IDinst/n10848 ,
         \IDinst/n10847 , \IDinst/n10846 , \IDinst/n10845 , \IDinst/n10844 ,
         \IDinst/n10843 , \IDinst/n10842 , \IDinst/n10841 , \IDinst/n10840 ,
         \IDinst/n10839 , \IDinst/n10838 , \IDinst/n10837 , \IDinst/n10836 ,
         \IDinst/n10835 , \IDinst/n10834 , \IDinst/n10833 , \IDinst/n10832 ,
         \IDinst/n10831 , \IDinst/n10830 , \IDinst/n10829 , \IDinst/n10828 ,
         \IDinst/n10827 , \IDinst/n10826 , \IDinst/n10825 , \IDinst/n10824 ,
         \IDinst/n10823 , \IDinst/n10822 , \IDinst/n10821 , \IDinst/n10820 ,
         \IDinst/n10819 , \IDinst/n10818 , \IDinst/n10817 , \IDinst/n10816 ,
         \IDinst/n10815 , \IDinst/n10814 , \IDinst/n10813 , \IDinst/n10812 ,
         \IDinst/n10811 , \IDinst/n10810 , \IDinst/n10809 , \IDinst/n10808 ,
         \IDinst/n10807 , \IDinst/n10806 , \IDinst/n10805 , \IDinst/n10804 ,
         \IDinst/n10803 , \IDinst/n10802 , \IDinst/n10801 , \IDinst/n10800 ,
         \IDinst/n10799 , \IDinst/n10798 , \IDinst/n10797 , \IDinst/n10796 ,
         \IDinst/n10795 , \IDinst/n10794 , \IDinst/n10793 , \IDinst/n10792 ,
         \IDinst/n10791 , \IDinst/n10790 , \IDinst/n10789 , \IDinst/n10788 ,
         \IDinst/n10787 , \IDinst/n10786 , \IDinst/n10785 , \IDinst/n10784 ,
         \IDinst/n10783 , \IDinst/n10782 , \IDinst/n10781 , \IDinst/n10780 ,
         \IDinst/n10779 , \IDinst/n10778 , \IDinst/n10777 , \IDinst/n10776 ,
         \IDinst/n10775 , \IDinst/n10774 , \IDinst/n10773 , \IDinst/n10772 ,
         \IDinst/n10771 , \IDinst/n10770 , \IDinst/n10769 , \IDinst/n10768 ,
         \IDinst/n10767 , \IDinst/n10766 , \IDinst/n10765 , \IDinst/n10764 ,
         \IDinst/n10763 , \IDinst/n10762 , \IDinst/n10761 , \IDinst/n10760 ,
         \IDinst/n10759 , \IDinst/n10758 , \IDinst/n10757 , \IDinst/n10756 ,
         \IDinst/n10755 , \IDinst/n10754 , \IDinst/n10753 , \IDinst/n10752 ,
         \IDinst/n10751 , \IDinst/n10750 , \IDinst/n10749 , \IDinst/n10748 ,
         \IDinst/n10747 , \IDinst/n10746 , \IDinst/n10745 , \IDinst/n10744 ,
         \IDinst/n10743 , \IDinst/n10742 , \IDinst/n10741 , \IDinst/n10740 ,
         \IDinst/n10739 , \IDinst/n10738 , \IDinst/n10737 , \IDinst/n10736 ,
         \IDinst/n10735 , \IDinst/n10734 , \IDinst/n10733 , \IDinst/n10732 ,
         \IDinst/n10731 , \IDinst/n10730 , \IDinst/n10729 , \IDinst/n10728 ,
         \IDinst/n10727 , \IDinst/n10726 , \IDinst/n10725 , \IDinst/n10724 ,
         \IDinst/n10723 , \IDinst/n10722 , \IDinst/n10721 , \IDinst/n10720 ,
         \IDinst/n10719 , \IDinst/n10718 , \IDinst/n10717 , \IDinst/n10716 ,
         \IDinst/n10715 , \IDinst/n10714 , \IDinst/n10713 , \IDinst/n10712 ,
         \IDinst/n10711 , \IDinst/n10710 , \IDinst/n10709 , \IDinst/n10708 ,
         \IDinst/n10707 , \IDinst/n10706 , \IDinst/n10705 , \IDinst/n10704 ,
         \IDinst/n10703 , \IDinst/n10702 , \IDinst/n10701 , \IDinst/n10700 ,
         \IDinst/n10699 , \IDinst/n10698 , \IDinst/n10697 , \IDinst/n10696 ,
         \IDinst/n10695 , \IDinst/n10694 , \IDinst/n10693 , \IDinst/n10692 ,
         \IDinst/n10691 , \IDinst/n10690 , \IDinst/n10689 , \IDinst/n10688 ,
         \IDinst/n10687 , \IDinst/n10686 , \IDinst/n10685 , \IDinst/n10684 ,
         \IDinst/n10683 , \IDinst/n10682 , \IDinst/n10681 , \IDinst/n10680 ,
         \IDinst/n10679 , \IDinst/n10678 , \IDinst/n10677 , \IDinst/n10676 ,
         \IDinst/n10675 , \IDinst/n10674 , \IDinst/n10673 , \IDinst/n10672 ,
         \IDinst/n10671 , \IDinst/n10670 , \IDinst/n10669 , \IDinst/n10668 ,
         \IDinst/n10667 , \IDinst/n10666 , \IDinst/n10665 , \IDinst/n10664 ,
         \IDinst/n10663 , \IDinst/n10662 , \IDinst/n10661 , \IDinst/n10660 ,
         \IDinst/n10659 , \IDinst/n10658 , \IDinst/n10657 , \IDinst/n10656 ,
         \IDinst/n10655 , \IDinst/n10654 , \IDinst/n10653 , \IDinst/n10652 ,
         \IDinst/n10651 , \IDinst/n10650 , \IDinst/n10649 , \IDinst/n10648 ,
         \IDinst/n10647 , \IDinst/n10646 , \IDinst/n10645 , \IDinst/n10644 ,
         \IDinst/n10643 , \IDinst/n10642 , \IDinst/n10641 , \IDinst/n10640 ,
         \IDinst/n10639 , \IDinst/n10638 , \IDinst/n10637 , \IDinst/n10636 ,
         \IDinst/n10635 , \IDinst/n10634 , \IDinst/n10633 , \IDinst/n10632 ,
         \IDinst/n10631 , \IDinst/n10630 , \IDinst/n10629 , \IDinst/n10628 ,
         \IDinst/n10627 , \IDinst/n10626 , \IDinst/n10625 , \IDinst/n10624 ,
         \IDinst/n10623 , \IDinst/n10622 , \IDinst/n10621 , \IDinst/n10620 ,
         \IDinst/n10619 , \IDinst/n10618 , \IDinst/n10617 , \IDinst/n10616 ,
         \IDinst/n10615 , \IDinst/n10614 , \IDinst/n10613 , \IDinst/n10612 ,
         \IDinst/n10611 , \IDinst/n10610 , \IDinst/n10609 , \IDinst/n10608 ,
         \IDinst/n10607 , \IDinst/n10606 , \IDinst/n10605 , \IDinst/n10604 ,
         \IDinst/n10603 , \IDinst/n10602 , \IDinst/n10601 , \IDinst/n10600 ,
         \IDinst/n10599 , \IDinst/n10598 , \IDinst/n10597 , \IDinst/n10596 ,
         \IDinst/n10595 , \IDinst/n10594 , \IDinst/n10593 , \IDinst/n10592 ,
         \IDinst/n10591 , \IDinst/n10590 , \IDinst/n10589 , \IDinst/n10588 ,
         \IDinst/n10587 , \IDinst/n10586 , \IDinst/n10585 , \IDinst/n10584 ,
         \IDinst/n10583 , \IDinst/n10582 , \IDinst/n10581 , \IDinst/n10580 ,
         \IDinst/n10579 , \IDinst/n10578 , \IDinst/n10577 , \IDinst/n10576 ,
         \IDinst/n10575 , \IDinst/n10574 , \IDinst/n10573 , \IDinst/n10572 ,
         \IDinst/n10571 , \IDinst/n10570 , \IDinst/n10569 , \IDinst/n10568 ,
         \IDinst/n10567 , \IDinst/n10566 , \IDinst/n10565 , \IDinst/n10564 ,
         \IDinst/n10563 , \IDinst/n10562 , \IDinst/n10561 , \IDinst/n10560 ,
         \IDinst/n10559 , \IDinst/n10558 , \IDinst/n10557 , \IDinst/n10556 ,
         \IDinst/n10555 , \IDinst/n10554 , \IDinst/n10553 , \IDinst/n10552 ,
         \IDinst/n10551 , \IDinst/n10550 , \IDinst/n10549 , \IDinst/n10548 ,
         \IDinst/n10547 , \IDinst/n10546 , \IDinst/n10545 , \IDinst/n10544 ,
         \IDinst/n10543 , \IDinst/n10542 , \IDinst/n10541 , \IDinst/n10540 ,
         \IDinst/n10539 , \IDinst/n10538 , \IDinst/n10537 , \IDinst/n10536 ,
         \IDinst/n10535 , \IDinst/n10534 , \IDinst/n10533 , \IDinst/n10532 ,
         \IDinst/n10531 , \IDinst/n10530 , \IDinst/n10529 , \IDinst/n10528 ,
         \IDinst/n10527 , \IDinst/n10526 , \IDinst/n10525 , \IDinst/n10524 ,
         \IDinst/n10523 , \IDinst/n10522 , \IDinst/n10521 , \IDinst/n10520 ,
         \IDinst/n10519 , \IDinst/n10518 , \IDinst/n10517 , \IDinst/n10516 ,
         \IDinst/n10515 , \IDinst/n10514 , \IDinst/n10513 , \IDinst/n10512 ,
         \IDinst/n10511 , \IDinst/n10510 , \IDinst/n10509 , \IDinst/n10508 ,
         \IDinst/n10507 , \IDinst/n10506 , \IDinst/n10505 , \IDinst/n10504 ,
         \IDinst/n10503 , \IDinst/n10502 , \IDinst/n10501 , \IDinst/n10500 ,
         \IDinst/n10499 , \IDinst/n10498 , \IDinst/n10497 , \IDinst/n10496 ,
         \IDinst/n10495 , \IDinst/n10494 , \IDinst/n10493 , \IDinst/n10492 ,
         \IDinst/n10491 , \IDinst/n10490 , \IDinst/n10489 , \IDinst/n10488 ,
         \IDinst/n10487 , \IDinst/n10486 , \IDinst/n10485 , \IDinst/n10484 ,
         \IDinst/n10483 , \IDinst/n10482 , \IDinst/n10481 , \IDinst/n10480 ,
         \IDinst/n10479 , \IDinst/n10478 , \IDinst/n10477 , \IDinst/n10476 ,
         \IDinst/n10475 , \IDinst/n10474 , \IDinst/n10473 , \IDinst/n10472 ,
         \IDinst/n10471 , \IDinst/n10470 , \IDinst/n10469 , \IDinst/n10468 ,
         \IDinst/n10467 , \IDinst/n10466 , \IDinst/n10465 , \IDinst/n10464 ,
         \IDinst/n10463 , \IDinst/n10462 , \IDinst/n10461 , \IDinst/n10460 ,
         \IDinst/n10459 , \IDinst/n10458 , \IDinst/n10457 , \IDinst/n10456 ,
         \IDinst/n10455 , \IDinst/n10454 , \IDinst/n10453 , \IDinst/n10452 ,
         \IDinst/n10451 , \IDinst/n10450 , \IDinst/n10449 , \IDinst/n10448 ,
         \IDinst/n10447 , \IDinst/n10446 , \IDinst/n10445 , \IDinst/n10444 ,
         \IDinst/n10443 , \IDinst/n10442 , \IDinst/n10441 , \IDinst/n10440 ,
         \IDinst/n10439 , \IDinst/n10438 , \IDinst/n10437 , \IDinst/n10436 ,
         \IDinst/n10435 , \IDinst/n10434 , \IDinst/n10433 , \IDinst/n10432 ,
         \IDinst/n10431 , \IDinst/n10430 , \IDinst/n10429 , \IDinst/n10428 ,
         \IDinst/n10427 , \IDinst/n10426 , \IDinst/n10425 , \IDinst/n10424 ,
         \IDinst/n10423 , \IDinst/n10422 , \IDinst/n10421 , \IDinst/n10420 ,
         \IDinst/n10419 , \IDinst/n10418 , \IDinst/n10417 , \IDinst/n10416 ,
         \IDinst/n10415 , \IDinst/n10414 , \IDinst/n10413 , \IDinst/n10412 ,
         \IDinst/n10411 , \IDinst/n10410 , \IDinst/n10409 , \IDinst/n10408 ,
         \IDinst/n10407 , \IDinst/n10406 , \IDinst/n10405 , \IDinst/n10404 ,
         \IDinst/n10403 , \IDinst/n10402 , \IDinst/n10401 , \IDinst/n10400 ,
         \IDinst/n10399 , \IDinst/n10398 , \IDinst/n10397 , \IDinst/n10396 ,
         \IDinst/n10395 , \IDinst/n10394 , \IDinst/n10393 , \IDinst/n10392 ,
         \IDinst/n10391 , \IDinst/n10390 , \IDinst/n10389 , \IDinst/n10388 ,
         \IDinst/n10387 , \IDinst/n10386 , \IDinst/n10385 , \IDinst/n10384 ,
         \IDinst/n10383 , \IDinst/n10382 , \IDinst/n10381 , \IDinst/n10380 ,
         \IDinst/n10379 , \IDinst/n10378 , \IDinst/n10377 , \IDinst/n10376 ,
         \IDinst/n10375 , \IDinst/n10374 , \IDinst/n10373 , \IDinst/n10372 ,
         \IDinst/n10371 , \IDinst/n10370 , \IDinst/n10369 , \IDinst/n10368 ,
         \IDinst/n10367 , \IDinst/n10366 , \IDinst/n10365 , \IDinst/n10364 ,
         \IDinst/n10363 , \IDinst/n10362 , \IDinst/n10361 , \IDinst/n10360 ,
         \IDinst/n10359 , \IDinst/n10358 , \IDinst/n10357 , \IDinst/n10356 ,
         \IDinst/n10355 , \IDinst/n10354 , \IDinst/n10353 , \IDinst/n10352 ,
         \IDinst/n10351 , \IDinst/n10350 , \IDinst/n10349 , \IDinst/n10348 ,
         \IDinst/n10347 , \IDinst/n10346 , \IDinst/n10345 , \IDinst/n10344 ,
         \IDinst/n10343 , \IDinst/n10342 , \IDinst/n10341 , \IDinst/n10340 ,
         \IDinst/n10339 , \IDinst/n10338 , \IDinst/n10337 , \IDinst/n10336 ,
         \IDinst/n10335 , \IDinst/n10334 , \IDinst/n10333 , \IDinst/n10332 ,
         \IDinst/n10331 , \IDinst/n10330 , \IDinst/n10329 , \IDinst/n10328 ,
         \IDinst/n10327 , \IDinst/n10326 , \IDinst/n10325 , \IDinst/n10324 ,
         \IDinst/n10323 , \IDinst/n10322 , \IDinst/n10321 , \IDinst/n10320 ,
         \IDinst/n10319 , \IDinst/n10318 , \IDinst/n10317 , \IDinst/n10316 ,
         \IDinst/n10315 , \IDinst/n10314 , \IDinst/n10313 , \IDinst/n10312 ,
         \IDinst/n10311 , \IDinst/n10310 , \IDinst/n10309 , \IDinst/n10308 ,
         \IDinst/n10307 , \IDinst/n10306 , \IDinst/n10305 , \IDinst/n10304 ,
         \IDinst/n10303 , \IDinst/n10302 , \IDinst/n10301 , \IDinst/n10300 ,
         \IDinst/n10299 , \IDinst/n10298 , \IDinst/n10297 , \IDinst/n10296 ,
         \IDinst/n10295 , \IDinst/n10294 , \IDinst/n10293 , \IDinst/n10292 ,
         \IDinst/n10291 , \IDinst/n10290 , \IDinst/n10289 , \IDinst/n10288 ,
         \IDinst/n10287 , \IDinst/n10286 , \IDinst/n10285 , \IDinst/n10284 ,
         \IDinst/n10283 , \IDinst/n10282 , \IDinst/n10281 , \IDinst/n10280 ,
         \IDinst/n10279 , \IDinst/n10278 , \IDinst/n10277 , \IDinst/n10276 ,
         \IDinst/n10275 , \IDinst/n10274 , \IDinst/n10273 , \IDinst/n10272 ,
         \IDinst/n10271 , \IDinst/n10270 , \IDinst/n10269 , \IDinst/n10268 ,
         \IDinst/n10267 , \IDinst/n10266 , \IDinst/n10265 , \IDinst/n10264 ,
         \IDinst/n10263 , \IDinst/n10262 , \IDinst/n10261 , \IDinst/n10260 ,
         \IDinst/n10259 , \IDinst/n10258 , \IDinst/n10257 , \IDinst/n10256 ,
         \IDinst/n10255 , \IDinst/n10254 , \IDinst/n10253 , \IDinst/n10252 ,
         \IDinst/n10251 , \IDinst/n10250 , \IDinst/n10249 , \IDinst/n10248 ,
         \IDinst/n10247 , \IDinst/n10246 , \IDinst/n10245 , \IDinst/n10244 ,
         \IDinst/n10243 , \IDinst/n10242 , \IDinst/n10241 , \IDinst/n10240 ,
         \IDinst/n10239 , \IDinst/n10238 , \IDinst/n10237 , \IDinst/n10236 ,
         \IDinst/n10235 , \IDinst/n10234 , \IDinst/n10233 , \IDinst/n10232 ,
         \IDinst/n10231 , \IDinst/n10230 , \IDinst/n10229 , \IDinst/n10228 ,
         \IDinst/n10227 , \IDinst/n10226 , \IDinst/n10225 , \IDinst/n10224 ,
         \IDinst/n10223 , \IDinst/n10222 , \IDinst/n10221 , \IDinst/n10220 ,
         \IDinst/n10219 , \IDinst/n10218 , \IDinst/n10217 , \IDinst/n10216 ,
         \IDinst/n10215 , \IDinst/n10214 , \IDinst/n10213 , \IDinst/n10212 ,
         \IDinst/n10211 , \IDinst/n10210 , \IDinst/n10209 , \IDinst/n10208 ,
         \IDinst/n10207 , \IDinst/n10206 , \IDinst/n10205 , \IDinst/n10204 ,
         \IDinst/n10203 , \IDinst/n10202 , \IDinst/n10201 , \IDinst/n10200 ,
         \IDinst/n10199 , \IDinst/n10198 , \IDinst/n10197 , \IDinst/n10196 ,
         \IDinst/n10195 , \IDinst/n10194 , \IDinst/n10193 , \IDinst/n10192 ,
         \IDinst/n10191 , \IDinst/n10190 , \IDinst/n10189 , \IDinst/n10188 ,
         \IDinst/n10187 , \IDinst/n10186 , \IDinst/n10185 , \IDinst/n10184 ,
         \IDinst/n10183 , \IDinst/n10182 , \IDinst/n10181 , \IDinst/n10180 ,
         \IDinst/n10179 , \IDinst/n10178 , \IDinst/n10177 , \IDinst/n10176 ,
         \IDinst/n10175 , \IDinst/n10174 , \IDinst/n10173 , \IDinst/n10172 ,
         \IDinst/n10171 , \IDinst/n10170 , \IDinst/n10169 , \IDinst/n10168 ,
         \IDinst/n10167 , \IDinst/n10166 , \IDinst/n10165 , \IDinst/n10164 ,
         \IDinst/n10163 , \IDinst/n10162 , \IDinst/n10161 , \IDinst/n10160 ,
         \IDinst/n10159 , \IDinst/n10158 , \IDinst/n10157 , \IDinst/n10156 ,
         \IDinst/n10155 , \IDinst/n10154 , \IDinst/n10153 , \IDinst/n10152 ,
         \IDinst/n10151 , \IDinst/n10150 , \IDinst/n10149 , \IDinst/n10148 ,
         \IDinst/n10147 , \IDinst/n10146 , \IDinst/n10145 , \IDinst/n10144 ,
         \IDinst/n10143 , \IDinst/n10142 , \IDinst/n10141 , \IDinst/n10140 ,
         \IDinst/n10139 , \IDinst/n10138 , \IDinst/n10137 , \IDinst/n10136 ,
         \IDinst/n10135 , \IDinst/n10134 , \IDinst/n10133 , \IDinst/n10132 ,
         \IDinst/n10131 , \IDinst/n10130 , \IDinst/n10129 , \IDinst/n10128 ,
         \IDinst/n10127 , \IDinst/n10126 , \IDinst/n10125 , \IDinst/n10124 ,
         \IDinst/n10123 , \IDinst/n10122 , \IDinst/n10121 , \IDinst/n10120 ,
         \IDinst/n10119 , \IDinst/n10118 , \IDinst/n10117 , \IDinst/n10116 ,
         \IDinst/n10115 , \IDinst/n10114 , \IDinst/n10113 , \IDinst/n10112 ,
         \IDinst/n10111 , \IDinst/n10110 , \IDinst/n10109 , \IDinst/n10108 ,
         \IDinst/n10107 , \IDinst/n10106 , \IDinst/n10105 , \IDinst/n10104 ,
         \IDinst/n10103 , \IDinst/n10102 , \IDinst/n10101 , \IDinst/n10100 ,
         \IDinst/n10099 , \IDinst/n10098 , \IDinst/n10097 , \IDinst/n10096 ,
         \IDinst/n10095 , \IDinst/n10094 , \IDinst/n10093 , \IDinst/n10092 ,
         \IDinst/n10091 , \IDinst/n10090 , \IDinst/n10089 , \IDinst/n10088 ,
         \IDinst/n10087 , \IDinst/n10086 , \IDinst/n10085 , \IDinst/n10084 ,
         \IDinst/n10083 , \IDinst/n10082 , \IDinst/n10081 , \IDinst/n10080 ,
         \IDinst/n10079 , \IDinst/n10078 , \IDinst/n10077 , \IDinst/n10076 ,
         \IDinst/n10075 , \IDinst/n10074 , \IDinst/n10073 , \IDinst/n10072 ,
         \IDinst/n10071 , \IDinst/n10070 , \IDinst/n10069 , \IDinst/n10068 ,
         \IDinst/n10067 , \IDinst/n10066 , \IDinst/n10065 , \IDinst/n10064 ,
         \IDinst/n10063 , \IDinst/n10062 , \IDinst/n10061 , \IDinst/n10060 ,
         \IDinst/n10059 , \IDinst/n10058 , \IDinst/n10057 , \IDinst/n10056 ,
         \IDinst/n10055 , \IDinst/n10054 , \IDinst/n10053 , \IDinst/n10052 ,
         \IDinst/n10051 , \IDinst/n10050 , \IDinst/n10049 , \IDinst/n10048 ,
         \IDinst/n10047 , \IDinst/n10046 , \IDinst/n10045 , \IDinst/n10044 ,
         \IDinst/n10043 , \IDinst/n10042 , \IDinst/n10041 , \IDinst/n10040 ,
         \IDinst/n10039 , \IDinst/n10038 , \IDinst/n10037 , \IDinst/n10036 ,
         \IDinst/n10035 , \IDinst/n10034 , \IDinst/n10033 , \IDinst/n10032 ,
         \IDinst/n10031 , \IDinst/n10030 , \IDinst/n10029 , \IDinst/n10028 ,
         \IDinst/n10027 , \IDinst/n10026 , \IDinst/n10025 , \IDinst/n10024 ,
         \IDinst/n10023 , \IDinst/n10022 , \IDinst/n10021 , \IDinst/n10020 ,
         \IDinst/n10019 , \IDinst/n10018 , \IDinst/n10017 , \IDinst/n10016 ,
         \IDinst/n10015 , \IDinst/n10014 , \IDinst/n10013 , \IDinst/n10012 ,
         \IDinst/n10011 , \IDinst/n10010 , \IDinst/n10009 , \IDinst/n10008 ,
         \IDinst/n10007 , \IDinst/n10006 , \IDinst/n10005 , \IDinst/n10004 ,
         \IDinst/n10003 , \IDinst/n10002 , \IDinst/n10001 , \IDinst/n10000 ,
         \IDinst/n9999 , \IDinst/n9998 , \IDinst/n9997 , \IDinst/n9996 ,
         \IDinst/n9995 , \IDinst/n9994 , \IDinst/n9993 , \IDinst/n9992 ,
         \IDinst/n9991 , \IDinst/n9990 , \IDinst/n9989 , \IDinst/n9988 ,
         \IDinst/n9987 , \IDinst/n9986 , \IDinst/n9985 , \IDinst/n9984 ,
         \IDinst/n9983 , \IDinst/n9982 , \IDinst/n9981 , \IDinst/n9980 ,
         \IDinst/n9979 , \IDinst/n9978 , \IDinst/n9977 , \IDinst/n9976 ,
         \IDinst/n9975 , \IDinst/n9974 , \IDinst/n9973 , \IDinst/n9972 ,
         \IDinst/n9971 , \IDinst/n9970 , \IDinst/n9969 , \IDinst/n9968 ,
         \IDinst/n9967 , \IDinst/n9966 , \IDinst/n9965 , \IDinst/n9964 ,
         \IDinst/n9963 , \IDinst/n9962 , \IDinst/n9961 , \IDinst/n9960 ,
         \IDinst/n9959 , \IDinst/n9958 , \IDinst/n9957 , \IDinst/n9956 ,
         \IDinst/n9955 , \IDinst/n9954 , \IDinst/n9953 , \IDinst/n9952 ,
         \IDinst/n9951 , \IDinst/n9950 , \IDinst/n9949 , \IDinst/n9948 ,
         \IDinst/n9947 , \IDinst/n9946 , \IDinst/n9945 , \IDinst/n9944 ,
         \IDinst/n9943 , \IDinst/n9942 , \IDinst/n9941 , \IDinst/n9940 ,
         \IDinst/n9939 , \IDinst/n9938 , \IDinst/n9937 , \IDinst/n9936 ,
         \IDinst/n9935 , \IDinst/n9934 , \IDinst/n9933 , \IDinst/n9932 ,
         \IDinst/n9931 , \IDinst/n9930 , \IDinst/n9929 , \IDinst/n9928 ,
         \IDinst/n9927 , \IDinst/n9926 , \IDinst/n9925 , \IDinst/n9924 ,
         \IDinst/n9923 , \IDinst/n9922 , \IDinst/n9921 , \IDinst/n9920 ,
         \IDinst/n9919 , \IDinst/n9918 , \IDinst/n9917 , \IDinst/n9916 ,
         \IDinst/n9915 , \IDinst/n9914 , \IDinst/n9913 , \IDinst/n9912 ,
         \IDinst/n9911 , \IDinst/n9910 , \IDinst/n9909 , \IDinst/n9908 ,
         \IDinst/n9907 , \IDinst/n9906 , \IDinst/n9905 , \IDinst/n9904 ,
         \IDinst/n9903 , \IDinst/n9902 , \IDinst/n9901 , \IDinst/n9900 ,
         \IDinst/n9899 , \IDinst/n9898 , \IDinst/n9897 , \IDinst/n9896 ,
         \IDinst/n9895 , \IDinst/n9894 , \IDinst/n9893 , \IDinst/n9892 ,
         \IDinst/n9891 , \IDinst/n9890 , \IDinst/n9889 , \IDinst/n9888 ,
         \IDinst/n9887 , \IDinst/n9886 , \IDinst/n9885 , \IDinst/n9884 ,
         \IDinst/n9883 , \IDinst/n9882 , \IDinst/n9881 , \IDinst/n9880 ,
         \IDinst/n9879 , \IDinst/n9878 , \IDinst/n9877 , \IDinst/n9876 ,
         \IDinst/n9875 , \IDinst/n9874 , \IDinst/n9873 , \IDinst/n9872 ,
         \IDinst/n9871 , \IDinst/n9870 , \IDinst/n9869 , \IDinst/n9868 ,
         \IDinst/n9867 , \IDinst/n9866 , \IDinst/n9865 , \IDinst/n9864 ,
         \IDinst/n9863 , \IDinst/n9862 , \IDinst/n9861 , \IDinst/n9860 ,
         \IDinst/n9859 , \IDinst/n9858 , \IDinst/n9857 , \IDinst/n9856 ,
         \IDinst/n9855 , \IDinst/n9854 , \IDinst/n9853 , \IDinst/n9852 ,
         \IDinst/n9851 , \IDinst/n9850 , \IDinst/n9849 , \IDinst/n9848 ,
         \IDinst/n9847 , \IDinst/n9846 , \IDinst/n9845 , \IDinst/n9844 ,
         \IDinst/n9843 , \IDinst/n9842 , \IDinst/n9841 , \IDinst/n9840 ,
         \IDinst/n9839 , \IDinst/n9838 , \IDinst/n9837 , \IDinst/n9836 ,
         \IDinst/n9835 , \IDinst/n9834 , \IDinst/n9833 , \IDinst/n9832 ,
         \IDinst/n9831 , \IDinst/n9830 , \IDinst/n9829 , \IDinst/n9828 ,
         \IDinst/n9827 , \IDinst/n9826 , \IDinst/n9825 , \IDinst/n9824 ,
         \IDinst/n9823 , \IDinst/n9822 , \IDinst/n9821 , \IDinst/n9820 ,
         \IDinst/n9819 , \IDinst/n9818 , \IDinst/n9817 , \IDinst/n9816 ,
         \IDinst/n9815 , \IDinst/n9814 , \IDinst/n9813 , \IDinst/n9812 ,
         \IDinst/n9811 , \IDinst/n9810 , \IDinst/n9809 , \IDinst/n9808 ,
         \IDinst/n9807 , \IDinst/n9806 , \IDinst/n9805 , \IDinst/n9804 ,
         \IDinst/n9803 , \IDinst/n9802 , \IDinst/n9801 , \IDinst/n9800 ,
         \IDinst/n9799 , \IDinst/n9798 , \IDinst/n9797 , \IDinst/n9796 ,
         \IDinst/n9795 , \IDinst/n9794 , \IDinst/n9793 , \IDinst/n9792 ,
         \IDinst/n9791 , \IDinst/n9790 , \IDinst/n9789 , \IDinst/n9788 ,
         \IDinst/n9787 , \IDinst/n9786 , \IDinst/n9785 , \IDinst/n9784 ,
         \IDinst/n9783 , \IDinst/n9782 , \IDinst/n9781 , \IDinst/n9780 ,
         \IDinst/n9779 , \IDinst/n9778 , \IDinst/n9777 , \IDinst/n9776 ,
         \IDinst/n9775 , \IDinst/n9774 , \IDinst/n9773 , \IDinst/n9772 ,
         \IDinst/n9771 , \IDinst/n9770 , \IDinst/n9769 , \IDinst/n9768 ,
         \IDinst/n9767 , \IDinst/n9766 , \IDinst/n9765 , \IDinst/n9764 ,
         \IDinst/n9763 , \IDinst/n9762 , \IDinst/n9761 , \IDinst/n9760 ,
         \IDinst/n9759 , \IDinst/n9758 , \IDinst/n9757 , \IDinst/n9756 ,
         \IDinst/n9755 , \IDinst/n9754 , \IDinst/n9753 , \IDinst/n9752 ,
         \IDinst/n9751 , \IDinst/n9750 , \IDinst/n9749 , \IDinst/n9748 ,
         \IDinst/n9747 , \IDinst/n9746 , \IDinst/n9745 , \IDinst/n9744 ,
         \IDinst/n9743 , \IDinst/n9742 , \IDinst/n9741 , \IDinst/n9740 ,
         \IDinst/n9739 , \IDinst/n9738 , \IDinst/n9737 , \IDinst/n9736 ,
         \IDinst/n9735 , \IDinst/n9734 , \IDinst/n9733 , \IDinst/n9732 ,
         \IDinst/n9731 , \IDinst/n9730 , \IDinst/n9729 , \IDinst/n9728 ,
         \IDinst/n9727 , \IDinst/n9726 , \IDinst/n9725 , \IDinst/n9724 ,
         \IDinst/n9723 , \IDinst/n9722 , \IDinst/n9721 , \IDinst/n9720 ,
         \IDinst/n9719 , \IDinst/n9718 , \IDinst/n9717 , \IDinst/n9716 ,
         \IDinst/n9715 , \IDinst/n9714 , \IDinst/n9713 , \IDinst/n9712 ,
         \IDinst/n9711 , \IDinst/n9710 , \IDinst/n9709 , \IDinst/n9708 ,
         \IDinst/n9707 , \IDinst/n9706 , \IDinst/n9705 , \IDinst/n9704 ,
         \IDinst/n9703 , \IDinst/n9702 , \IDinst/n9701 , \IDinst/n9700 ,
         \IDinst/n9699 , \IDinst/n9698 , \IDinst/n9697 , \IDinst/n9696 ,
         \IDinst/n9695 , \IDinst/n9694 , \IDinst/n9693 , \IDinst/n9692 ,
         \IDinst/n9691 , \IDinst/n9690 , \IDinst/n9689 , \IDinst/n9688 ,
         \IDinst/n9687 , \IDinst/n9686 , \IDinst/n9685 , \IDinst/n9684 ,
         \IDinst/n9683 , \IDinst/n9682 , \IDinst/n9681 , \IDinst/n9680 ,
         \IDinst/n9679 , \IDinst/n9678 , \IDinst/n9677 , \IDinst/n9676 ,
         \IDinst/n9675 , \IDinst/n9674 , \IDinst/n9673 , \IDinst/n9672 ,
         \IDinst/n9671 , \IDinst/n9670 , \IDinst/n9669 , \IDinst/n9668 ,
         \IDinst/n9667 , \IDinst/n9666 , \IDinst/n9665 , \IDinst/n9664 ,
         \IDinst/n9663 , \IDinst/n9662 , \IDinst/n9661 , \IDinst/n9660 ,
         \IDinst/n9659 , \IDinst/n9658 , \IDinst/n9657 , \IDinst/n9656 ,
         \IDinst/n9655 , \IDinst/n9654 , \IDinst/n9653 , \IDinst/n9652 ,
         \IDinst/n9651 , \IDinst/n9650 , \IDinst/n9649 , \IDinst/n9648 ,
         \IDinst/n9647 , \IDinst/n9646 , \IDinst/n9645 , \IDinst/n9644 ,
         \IDinst/n9643 , \IDinst/n9642 , \IDinst/n9641 , \IDinst/n9640 ,
         \IDinst/n9639 , \IDinst/n9638 , \IDinst/n9637 , \IDinst/n9636 ,
         \IDinst/n9635 , \IDinst/n9634 , \IDinst/n9633 , \IDinst/n9632 ,
         \IDinst/n9631 , \IDinst/n9630 , \IDinst/n9629 , \IDinst/n9628 ,
         \IDinst/n9627 , \IDinst/n9626 , \IDinst/n9625 , \IDinst/n9624 ,
         \IDinst/n9623 , \IDinst/n9622 , \IDinst/n9621 , \IDinst/n9620 ,
         \IDinst/n9619 , \IDinst/n9618 , \IDinst/n9617 , \IDinst/n9616 ,
         \IDinst/n9615 , \IDinst/n9614 , \IDinst/n9613 , \IDinst/n9612 ,
         \IDinst/n9611 , \IDinst/n9610 , \IDinst/n9609 , \IDinst/n9608 ,
         \IDinst/n9607 , \IDinst/n9606 , \IDinst/n9605 , \IDinst/n9604 ,
         \IDinst/n9603 , \IDinst/n9602 , \IDinst/n9601 , \IDinst/n9600 ,
         \IDinst/n9599 , \IDinst/n9598 , \IDinst/n9597 , \IDinst/n9596 ,
         \IDinst/n9595 , \IDinst/n9594 , \IDinst/n9593 , \IDinst/n9592 ,
         \IDinst/n9591 , \IDinst/n9590 , \IDinst/n9589 , \IDinst/n9588 ,
         \IDinst/n9587 , \IDinst/n9586 , \IDinst/n9585 , \IDinst/n9584 ,
         \IDinst/n9583 , \IDinst/n9582 , \IDinst/n9581 , \IDinst/n9580 ,
         \IDinst/n9579 , \IDinst/n9578 , \IDinst/n9577 , \IDinst/n9576 ,
         \IDinst/n9575 , \IDinst/n9574 , \IDinst/n9573 , \IDinst/n9572 ,
         \IDinst/n9571 , \IDinst/n9570 , \IDinst/n9569 , \IDinst/n9568 ,
         \IDinst/n9567 , \IDinst/n9566 , \IDinst/n9565 , \IDinst/n9564 ,
         \IDinst/n9563 , \IDinst/n9562 , \IDinst/n9561 , \IDinst/n9560 ,
         \IDinst/n9559 , \IDinst/n9558 , \IDinst/n9557 , \IDinst/n9556 ,
         \IDinst/n9555 , \IDinst/n9554 , \IDinst/n9553 , \IDinst/n9552 ,
         \IDinst/n9551 , \IDinst/n9550 , \IDinst/n9549 , \IDinst/n9548 ,
         \IDinst/n9547 , \IDinst/n9546 , \IDinst/n9545 , \IDinst/n9544 ,
         \IDinst/n9543 , \IDinst/n9542 , \IDinst/n9541 , \IDinst/n9540 ,
         \IDinst/n9539 , \IDinst/n9538 , \IDinst/n9537 , \IDinst/n9536 ,
         \IDinst/n9535 , \IDinst/n9534 , \IDinst/n9533 , \IDinst/n9532 ,
         \IDinst/n9531 , \IDinst/n9530 , \IDinst/n9529 , \IDinst/n9528 ,
         \IDinst/n9527 , \IDinst/n9526 , \IDinst/n9525 , \IDinst/n9524 ,
         \IDinst/n9523 , \IDinst/n9522 , \IDinst/n9521 , \IDinst/n9520 ,
         \IDinst/n9519 , \IDinst/n9518 , \IDinst/n9517 , \IDinst/n9516 ,
         \IDinst/n9515 , \IDinst/n9514 , \IDinst/n9513 , \IDinst/n9512 ,
         \IDinst/n9511 , \IDinst/n9510 , \IDinst/n9509 , \IDinst/n9508 ,
         \IDinst/n9507 , \IDinst/n9506 , \IDinst/n9505 , \IDinst/n9504 ,
         \IDinst/n9503 , \IDinst/n9502 , \IDinst/n9501 , \IDinst/n9500 ,
         \IDinst/n9499 , \IDinst/n9498 , \IDinst/n9497 , \IDinst/n9496 ,
         \IDinst/n9495 , \IDinst/n9494 , \IDinst/n9493 , \IDinst/n9492 ,
         \IDinst/n9491 , \IDinst/n9490 , \IDinst/n9489 , \IDinst/n9488 ,
         \IDinst/n9487 , \IDinst/n9486 , \IDinst/n9485 , \IDinst/n9484 ,
         \IDinst/n9483 , \IDinst/n9482 , \IDinst/n9481 , \IDinst/n9480 ,
         \IDinst/n9479 , \IDinst/n9478 , \IDinst/n9477 , \IDinst/n9476 ,
         \IDinst/n9475 , \IDinst/n9474 , \IDinst/n9473 , \IDinst/n9472 ,
         \IDinst/n9471 , \IDinst/n9470 , \IDinst/n9469 , \IDinst/n9468 ,
         \IDinst/n9467 , \IDinst/n9466 , \IDinst/n9465 , \IDinst/n9464 ,
         \IDinst/n9463 , \IDinst/n9462 , \IDinst/n9461 , \IDinst/n9460 ,
         \IDinst/n9459 , \IDinst/n9458 , \IDinst/n9457 , \IDinst/n9456 ,
         \IDinst/n9455 , \IDinst/n9454 , \IDinst/n9453 , \IDinst/n9452 ,
         \IDinst/n9451 , \IDinst/n9450 , \IDinst/n9449 , \IDinst/n9448 ,
         \IDinst/n9447 , \IDinst/n9446 , \IDinst/n9445 , \IDinst/n9444 ,
         \IDinst/n9443 , \IDinst/n9442 , \IDinst/n9441 , \IDinst/n9440 ,
         \IDinst/n9439 , \IDinst/n9438 , \IDinst/n9437 , \IDinst/n9436 ,
         \IDinst/n9435 , \IDinst/n9434 , \IDinst/n9433 , \IDinst/n9432 ,
         \IDinst/n9431 , \IDinst/n9430 , \IDinst/n9429 , \IDinst/n9428 ,
         \IDinst/n9427 , \IDinst/n9426 , \IDinst/n9425 , \IDinst/n9424 ,
         \IDinst/n9423 , \IDinst/n9422 , \IDinst/n9421 , \IDinst/n9420 ,
         \IDinst/n9419 , \IDinst/n9418 , \IDinst/n9417 , \IDinst/n9416 ,
         \IDinst/n9415 , \IDinst/n9414 , \IDinst/n9413 , \IDinst/n9412 ,
         \IDinst/n9411 , \IDinst/n9410 , \IDinst/n9409 , \IDinst/n9408 ,
         \IDinst/n9407 , \IDinst/n9406 , \IDinst/n9405 , \IDinst/n9404 ,
         \IDinst/n9403 , \IDinst/n9402 , \IDinst/n9401 , \IDinst/n9400 ,
         \IDinst/n9399 , \IDinst/n9398 , \IDinst/n9397 , \IDinst/n9396 ,
         \IDinst/n9395 , \IDinst/n9394 , \IDinst/n9393 , \IDinst/n9392 ,
         \IDinst/n9391 , \IDinst/n9390 , \IDinst/n9389 , \IDinst/n9388 ,
         \IDinst/n9387 , \IDinst/n9386 , \IDinst/n9385 , \IDinst/n9384 ,
         \IDinst/n9383 , \IDinst/n9382 , \IDinst/n9381 , \IDinst/n9380 ,
         \IDinst/n9379 , \IDinst/n9378 , \IDinst/n9377 , \IDinst/n9376 ,
         \IDinst/n9375 , \IDinst/n9374 , \IDinst/n9373 , \IDinst/n9372 ,
         \IDinst/n9371 , \IDinst/n9370 , \IDinst/n9369 , \IDinst/n9368 ,
         \IDinst/n9367 , \IDinst/n9366 , \IDinst/n9365 , \IDinst/n9364 ,
         \IDinst/n9363 , \IDinst/n9362 , \IDinst/n9361 , \IDinst/n9360 ,
         \IDinst/n9359 , \IDinst/n9358 , \IDinst/n9357 , \IDinst/n9356 ,
         \IDinst/n9355 , \IDinst/n9354 , \IDinst/n9353 , \IDinst/n9352 ,
         \IDinst/n9351 , \IDinst/n9350 , \IDinst/n9349 , \IDinst/n9348 ,
         \IDinst/n9347 , \IDinst/n9346 , \IDinst/n9345 , \IDinst/n9344 ,
         \IDinst/n9343 , \IDinst/n9342 , \IDinst/n9341 , \IDinst/n9340 ,
         \IDinst/n9339 , \IDinst/n9338 , \IDinst/n9337 , \IDinst/n9336 ,
         \IDinst/n9335 , \IDinst/n9334 , \IDinst/n9333 , \IDinst/n9332 ,
         \IDinst/n9331 , \IDinst/n9330 , \IDinst/n9329 , \IDinst/n9328 ,
         \IDinst/n9327 , \IDinst/n9326 , \IDinst/n9325 , \IDinst/n9324 ,
         \IDinst/n9323 , \IDinst/n9322 , \IDinst/n9321 , \IDinst/n9320 ,
         \IDinst/n9319 , \IDinst/n9318 , \IDinst/n9317 , \IDinst/n9316 ,
         \IDinst/n9315 , \IDinst/n9314 , \IDinst/n9313 , \IDinst/n9312 ,
         \IDinst/n9311 , \IDinst/n9310 , \IDinst/n9309 , \IDinst/n9308 ,
         \IDinst/n9307 , \IDinst/n9306 , \IDinst/n9305 , \IDinst/n9304 ,
         \IDinst/n9303 , \IDinst/n9302 , \IDinst/n9301 , \IDinst/n9300 ,
         \IDinst/n9299 , \IDinst/n9298 , \IDinst/n9297 , \IDinst/n9296 ,
         \IDinst/n9295 , \IDinst/n9294 , \IDinst/n9293 , \IDinst/n9292 ,
         \IDinst/n9291 , \IDinst/n9290 , \IDinst/n9289 , \IDinst/n9288 ,
         \IDinst/n9287 , \IDinst/n9286 , \IDinst/n9285 , \IDinst/n9284 ,
         \IDinst/n9283 , \IDinst/n9282 , \IDinst/n9281 , \IDinst/n9280 ,
         \IDinst/n9279 , \IDinst/n9278 , \IDinst/n9277 , \IDinst/n9276 ,
         \IDinst/n9275 , \IDinst/n9274 , \IDinst/n9273 , \IDinst/n9272 ,
         \IDinst/n9271 , \IDinst/n9270 , \IDinst/n9269 , \IDinst/n9268 ,
         \IDinst/n9267 , \IDinst/n9266 , \IDinst/n9265 , \IDinst/n9264 ,
         \IDinst/n9263 , \IDinst/n9262 , \IDinst/n9261 , \IDinst/n9260 ,
         \IDinst/n9259 , \IDinst/n9258 , \IDinst/n9257 , \IDinst/n9256 ,
         \IDinst/n9255 , \IDinst/n9254 , \IDinst/n9253 , \IDinst/n9252 ,
         \IDinst/n9251 , \IDinst/n9250 , \IDinst/n9249 , \IDinst/n9248 ,
         \IDinst/n9247 , \IDinst/n9246 , \IDinst/n9245 , \IDinst/n9244 ,
         \IDinst/n9243 , \IDinst/n9242 , \IDinst/n9241 , \IDinst/n9240 ,
         \IDinst/n9239 , \IDinst/n9238 , \IDinst/n9237 , \IDinst/n9236 ,
         \IDinst/n9235 , \IDinst/n9234 , \IDinst/n9233 , \IDinst/n9232 ,
         \IDinst/n9231 , \IDinst/n9230 , \IDinst/n9229 , \IDinst/n9228 ,
         \IDinst/n9227 , \IDinst/n9226 , \IDinst/n9225 , \IDinst/n9224 ,
         \IDinst/n9223 , \IDinst/n9222 , \IDinst/n9221 , \IDinst/n9220 ,
         \IDinst/n9219 , \IDinst/n9218 , \IDinst/n9217 , \IDinst/n9216 ,
         \IDinst/n9215 , \IDinst/n9214 , \IDinst/n9213 , \IDinst/n9212 ,
         \IDinst/n9211 , \IDinst/n9210 , \IDinst/n9209 , \IDinst/n9208 ,
         \IDinst/n9207 , \IDinst/n9206 , \IDinst/n9205 , \IDinst/n9204 ,
         \IDinst/n9203 , \IDinst/n9202 , \IDinst/n9201 , \IDinst/n9200 ,
         \IDinst/n9199 , \IDinst/n9198 , \IDinst/n9197 , \IDinst/n9196 ,
         \IDinst/n9195 , \IDinst/n9194 , \IDinst/n9193 , \IDinst/n9192 ,
         \IDinst/n9191 , \IDinst/n9190 , \IDinst/n9189 , \IDinst/n9188 ,
         \IDinst/n9187 , \IDinst/n9186 , \IDinst/n9185 , \IDinst/n9184 ,
         \IDinst/n9183 , \IDinst/n9182 , \IDinst/n9181 , \IDinst/n9180 ,
         \IDinst/n9179 , \IDinst/n9178 , \IDinst/n9177 , \IDinst/n9176 ,
         \IDinst/n9175 , \IDinst/n9174 , \IDinst/n9173 , \IDinst/n9172 ,
         \IDinst/n9171 , \IDinst/n9170 , \IDinst/n9169 , \IDinst/n9168 ,
         \IDinst/n9167 , \IDinst/n9166 , \IDinst/n9165 , \IDinst/n9164 ,
         \IDinst/n9163 , \IDinst/n9162 , \IDinst/n9161 , \IDinst/n9160 ,
         \IDinst/n9159 , \IDinst/n9158 , \IDinst/n9157 , \IDinst/n9156 ,
         \IDinst/n9155 , \IDinst/n9154 , \IDinst/n9153 , \IDinst/n9152 ,
         \IDinst/n9151 , \IDinst/n9150 , \IDinst/n9149 , \IDinst/n9148 ,
         \IDinst/n9147 , \IDinst/n9146 , \IDinst/n9145 , \IDinst/n9144 ,
         \IDinst/n9143 , \IDinst/n9142 , \IDinst/n9141 , \IDinst/n9140 ,
         \IDinst/n9139 , \IDinst/n9138 , \IDinst/n9137 , \IDinst/n9136 ,
         \IDinst/n9135 , \IDinst/n9134 , \IDinst/n9133 , \IDinst/n9132 ,
         \IDinst/n9131 , \IDinst/n9130 , \IDinst/n9129 , \IDinst/n9128 ,
         \IDinst/n9127 , \IDinst/n9126 , \IDinst/n9125 , \IDinst/n9124 ,
         \IDinst/n9123 , \IDinst/n9122 , \IDinst/n9121 , \IDinst/n9120 ,
         \IDinst/n9119 , \IDinst/n9118 , \IDinst/n9117 , \IDinst/n9116 ,
         \IDinst/n9115 , \IDinst/n9114 , \IDinst/n9113 , \IDinst/n9112 ,
         \IDinst/n9111 , \IDinst/n9110 , \IDinst/n9109 , \IDinst/n9108 ,
         \IDinst/n9107 , \IDinst/n9106 , \IDinst/n9105 , \IDinst/n9104 ,
         \IDinst/n9103 , \IDinst/n9102 , \IDinst/n9101 , \IDinst/n9100 ,
         \IDinst/n9099 , \IDinst/n9098 , \IDinst/n9097 , \IDinst/n9096 ,
         \IDinst/n9095 , \IDinst/n9094 , \IDinst/n9093 , \IDinst/n9092 ,
         \IDinst/n9091 , \IDinst/n9090 , \IDinst/n9089 , \IDinst/n9088 ,
         \IDinst/n9087 , \IDinst/n9086 , \IDinst/n9085 , \IDinst/n9084 ,
         \IDinst/n9083 , \IDinst/n9082 , \IDinst/n9081 , \IDinst/n9080 ,
         \IDinst/n9079 , \IDinst/n9078 , \IDinst/n9077 , \IDinst/n9076 ,
         \IDinst/n9075 , \IDinst/n9074 , \IDinst/n9073 , \IDinst/n9072 ,
         \IDinst/n9071 , \IDinst/n9070 , \IDinst/n9069 , \IDinst/n9068 ,
         \IDinst/n9067 , \IDinst/n9066 , \IDinst/n9065 , \IDinst/n9064 ,
         \IDinst/n9063 , \IDinst/n9062 , \IDinst/n9061 , \IDinst/n9060 ,
         \IDinst/n9059 , \IDinst/n9058 , \IDinst/n9057 , \IDinst/n9056 ,
         \IDinst/n9055 , \IDinst/n9054 , \IDinst/n9053 , \IDinst/n9052 ,
         \IDinst/n9051 , \IDinst/n9050 , \IDinst/n9049 , \IDinst/n9048 ,
         \IDinst/n9047 , \IDinst/n9046 , \IDinst/n9045 , \IDinst/n9044 ,
         \IDinst/n9043 , \IDinst/n9042 , \IDinst/n9041 , \IDinst/n9040 ,
         \IDinst/n9039 , \IDinst/n9038 , \IDinst/n9037 , \IDinst/n9036 ,
         \IDinst/n9035 , \IDinst/n9034 , \IDinst/n9033 , \IDinst/n9032 ,
         \IDinst/n9031 , \IDinst/n9030 , \IDinst/n9029 , \IDinst/n9028 ,
         \IDinst/n9027 , \IDinst/n9026 , \IDinst/n9025 , \IDinst/n9024 ,
         \IDinst/n9023 , \IDinst/n9022 , \IDinst/n9021 , \IDinst/n9020 ,
         \IDinst/n9019 , \IDinst/n9018 , \IDinst/n9017 , \IDinst/n9016 ,
         \IDinst/n9015 , \IDinst/n9014 , \IDinst/n9013 , \IDinst/n9012 ,
         \IDinst/n9011 , \IDinst/n9010 , \IDinst/n9009 , \IDinst/n9008 ,
         \IDinst/n9007 , \IDinst/n9006 , \IDinst/n9005 , \IDinst/n9004 ,
         \IDinst/n9003 , \IDinst/n9002 , \IDinst/n9001 , \IDinst/n9000 ,
         \IDinst/n8999 , \IDinst/n8998 , \IDinst/n8997 , \IDinst/n8996 ,
         \IDinst/n8995 , \IDinst/n8994 , \IDinst/n8993 , \IDinst/n8992 ,
         \IDinst/n8991 , \IDinst/n8990 , \IDinst/n8989 , \IDinst/n8988 ,
         \IDinst/n8987 , \IDinst/n8986 , \IDinst/n8985 , \IDinst/n8984 ,
         \IDinst/n8983 , \IDinst/n8982 , \IDinst/n8981 , \IDinst/n8980 ,
         \IDinst/n8979 , \IDinst/n8978 , \IDinst/n8977 , \IDinst/n8976 ,
         \IDinst/n8975 , \IDinst/n8974 , \IDinst/n8973 , \IDinst/n8972 ,
         \IDinst/n8971 , \IDinst/n8970 , \IDinst/n8969 , \IDinst/n8968 ,
         \IDinst/n8967 , \IDinst/n8966 , \IDinst/n8965 , \IDinst/n8964 ,
         \IDinst/n8963 , \IDinst/n8962 , \IDinst/n8961 , \IDinst/n8960 ,
         \IDinst/n8959 , \IDinst/n8958 , \IDinst/n8957 , \IDinst/n8956 ,
         \IDinst/n8955 , \IDinst/n8954 , \IDinst/n8953 , \IDinst/n8952 ,
         \IDinst/n8951 , \IDinst/n8950 , \IDinst/n8949 , \IDinst/n8948 ,
         \IDinst/n8947 , \IDinst/n8946 , \IDinst/n8945 , \IDinst/n8944 ,
         \IDinst/n8943 , \IDinst/n8942 , \IDinst/n8941 , \IDinst/n8940 ,
         \IDinst/n8939 , \IDinst/n8938 , \IDinst/n8937 , \IDinst/n8936 ,
         \IDinst/n8935 , \IDinst/n8934 , \IDinst/n8933 , \IDinst/n8932 ,
         \IDinst/n8931 , \IDinst/n8930 , \IDinst/n8929 , \IDinst/n8928 ,
         \IDinst/n8927 , \IDinst/n8926 , \IDinst/n8925 , \IDinst/n8924 ,
         \IDinst/n8923 , \IDinst/n8922 , \IDinst/n8921 , \IDinst/n8920 ,
         \IDinst/n8919 , \IDinst/n8918 , \IDinst/n8917 , \IDinst/n8916 ,
         \IDinst/n8915 , \IDinst/n8914 , \IDinst/n8913 , \IDinst/n8912 ,
         \IDinst/n8911 , \IDinst/n8910 , \IDinst/n8909 , \IDinst/n8908 ,
         \IDinst/n8907 , \IDinst/n8906 , \IDinst/n8905 , \IDinst/n8904 ,
         \IDinst/n8903 , \IDinst/n8902 , \IDinst/n8901 , \IDinst/n8900 ,
         \IDinst/n8899 , \IDinst/n8898 , \IDinst/n8897 , \IDinst/n8896 ,
         \IDinst/n8895 , \IDinst/n8894 , \IDinst/n8893 , \IDinst/n8892 ,
         \IDinst/n8891 , \IDinst/n8890 , \IDinst/n8889 , \IDinst/n8888 ,
         \IDinst/n8887 , \IDinst/n8886 , \IDinst/n8885 , \IDinst/n8884 ,
         \IDinst/n8883 , \IDinst/n8882 , \IDinst/n8881 , \IDinst/n8880 ,
         \IDinst/n8879 , \IDinst/n8878 , \IDinst/n8877 , \IDinst/n8876 ,
         \IDinst/n8875 , \IDinst/n8874 , \IDinst/n8873 , \IDinst/n8872 ,
         \IDinst/n8871 , \IDinst/n8870 , \IDinst/n8869 , \IDinst/n8868 ,
         \IDinst/n8867 , \IDinst/n8866 , \IDinst/n8865 , \IDinst/n8864 ,
         \IDinst/n8863 , \IDinst/n8862 , \IDinst/n8861 , \IDinst/n8860 ,
         \IDinst/n8859 , \IDinst/n8858 , \IDinst/n8857 , \IDinst/n8856 ,
         \IDinst/n8855 , \IDinst/n8854 , \IDinst/n8853 , \IDinst/n8852 ,
         \IDinst/n8851 , \IDinst/n8850 , \IDinst/n8849 , \IDinst/n8848 ,
         \IDinst/n8847 , \IDinst/n8846 , \IDinst/n8845 , \IDinst/n8844 ,
         \IDinst/n8843 , \IDinst/n8842 , \IDinst/n8841 , \IDinst/n8840 ,
         \IDinst/n8839 , \IDinst/n8838 , \IDinst/n8837 , \IDinst/n8836 ,
         \IDinst/n8835 , \IDinst/n8834 , \IDinst/n8833 , \IDinst/n8832 ,
         \IDinst/n8831 , \IDinst/n8830 , \IDinst/n8829 , \IDinst/n8828 ,
         \IDinst/n8827 , \IDinst/n8826 , \IDinst/n8825 , \IDinst/n8824 ,
         \IDinst/n8823 , \IDinst/n8822 , \IDinst/n8821 , \IDinst/n8820 ,
         \IDinst/n8819 , \IDinst/n8818 , \IDinst/n8817 , \IDinst/n8816 ,
         \IDinst/n8815 , \IDinst/n8814 , \IDinst/n8813 , \IDinst/n8812 ,
         \IDinst/n8811 , \IDinst/n8810 , \IDinst/n8809 , \IDinst/n8808 ,
         \IDinst/n8807 , \IDinst/n8806 , \IDinst/n8805 , \IDinst/n8804 ,
         \IDinst/n8803 , \IDinst/n8802 , \IDinst/n8801 , \IDinst/n8800 ,
         \IDinst/n8799 , \IDinst/n8798 , \IDinst/n8797 , \IDinst/n8796 ,
         \IDinst/n8795 , \IDinst/n8794 , \IDinst/n8793 , \IDinst/n8792 ,
         \IDinst/n8791 , \IDinst/n8790 , \IDinst/n8789 , \IDinst/n8788 ,
         \IDinst/n8787 , \IDinst/n8786 , \IDinst/n8785 , \IDinst/n8784 ,
         \IDinst/n8783 , \IDinst/n8782 , \IDinst/n8781 , \IDinst/n8780 ,
         \IDinst/n8779 , \IDinst/n8778 , \IDinst/n8777 , \IDinst/n8776 ,
         \IDinst/n8775 , \IDinst/n8774 , \IDinst/n8773 , \IDinst/n8772 ,
         \IDinst/n8771 , \IDinst/n8770 , \IDinst/n8769 , \IDinst/n8768 ,
         \IDinst/n8767 , \IDinst/n8766 , \IDinst/n8765 , \IDinst/n8764 ,
         \IDinst/n8763 , \IDinst/n8762 , \IDinst/n8761 , \IDinst/n8760 ,
         \IDinst/n8759 , \IDinst/n8758 , \IDinst/n8757 , \IDinst/n8756 ,
         \IDinst/n8755 , \IDinst/n8754 , \IDinst/n8753 , \IDinst/n8752 ,
         \IDinst/n8751 , \IDinst/n8750 , \IDinst/n8749 , \IDinst/n8748 ,
         \IDinst/n8747 , \IDinst/n8746 , \IDinst/n8745 , \IDinst/n8744 ,
         \IDinst/n8743 , \IDinst/n8742 , \IDinst/n8741 , \IDinst/n8740 ,
         \IDinst/n8739 , \IDinst/n8738 , \IDinst/n8737 , \IDinst/n8736 ,
         \IDinst/n8735 , \IDinst/n8734 , \IDinst/n8733 , \IDinst/n8732 ,
         \IDinst/n8731 , \IDinst/n8730 , \IDinst/n8729 , \IDinst/n8728 ,
         \IDinst/n8727 , \IDinst/n8726 , \IDinst/n8725 , \IDinst/n8724 ,
         \IDinst/n8723 , \IDinst/n8722 , \IDinst/n8721 , \IDinst/n8720 ,
         \IDinst/n8719 , \IDinst/n8718 , \IDinst/n8717 , \IDinst/n8716 ,
         \IDinst/n8715 , \IDinst/n8714 , \IDinst/n8713 , \IDinst/n8712 ,
         \IDinst/n8711 , \IDinst/n8710 , \IDinst/n8709 , \IDinst/n8708 ,
         \IDinst/n8707 , \IDinst/n8706 , \IDinst/n8705 , \IDinst/n8704 ,
         \IDinst/n8703 , \IDinst/n8702 , \IDinst/n8701 , \IDinst/n8700 ,
         \IDinst/n8699 , \IDinst/n8698 , \IDinst/n8697 , \IDinst/n8696 ,
         \IDinst/n8695 , \IDinst/n8694 , \IDinst/n8693 , \IDinst/n8692 ,
         \IDinst/n8691 , \IDinst/n8690 , \IDinst/n8689 , \IDinst/n8688 ,
         \IDinst/n8687 , \IDinst/n8686 , \IDinst/n8685 , \IDinst/n8684 ,
         \IDinst/n8683 , \IDinst/n8682 , \IDinst/n8681 , \IDinst/n8680 ,
         \IDinst/n8679 , \IDinst/n8678 , \IDinst/n8677 , \IDinst/n8676 ,
         \IDinst/n8675 , \IDinst/n8674 , \IDinst/n8673 , \IDinst/n8672 ,
         \IDinst/n8671 , \IDinst/n8670 , \IDinst/n8669 , \IDinst/n8668 ,
         \IDinst/n8667 , \IDinst/n8666 , \IDinst/n8665 , \IDinst/n8664 ,
         \IDinst/n8663 , \IDinst/n8662 , \IDinst/n8661 , \IDinst/n8660 ,
         \IDinst/n8659 , \IDinst/n8658 , \IDinst/n8657 , \IDinst/n8656 ,
         \IDinst/n8655 , \IDinst/n8654 , \IDinst/n8653 , \IDinst/n8652 ,
         \IDinst/n8651 , \IDinst/n8650 , \IDinst/n8649 , \IDinst/n8648 ,
         \IDinst/n8647 , \IDinst/n8646 , \IDinst/n8645 , \IDinst/n8644 ,
         \IDinst/n8643 , \IDinst/n8642 , \IDinst/n8641 , \IDinst/n8640 ,
         \IDinst/n8639 , \IDinst/n8638 , \IDinst/n8637 , \IDinst/n8636 ,
         \IDinst/n8635 , \IDinst/n8634 , \IDinst/n8633 , \IDinst/n8632 ,
         \IDinst/n8631 , \IDinst/n8630 , \IDinst/n8629 , \IDinst/n8628 ,
         \IDinst/n8627 , \IDinst/n8626 , \IDinst/n8625 , \IDinst/n8624 ,
         \IDinst/n8623 , \IDinst/n8622 , \IDinst/n8621 , \IDinst/n8620 ,
         \IDinst/n8619 , \IDinst/n8618 , \IDinst/n8617 , \IDinst/n8616 ,
         \IDinst/n8615 , \IDinst/n8614 , \IDinst/n8613 , \IDinst/n8612 ,
         \IDinst/n8611 , \IDinst/n8610 , \IDinst/n8609 , \IDinst/n8608 ,
         \IDinst/n8607 , \IDinst/n8606 , \IDinst/n8605 , \IDinst/n8604 ,
         \IDinst/n8603 , \IDinst/n8602 , \IDinst/n8601 , \IDinst/n8600 ,
         \IDinst/n8599 , \IDinst/n8598 , \IDinst/n8597 , \IDinst/n8596 ,
         \IDinst/n8595 , \IDinst/n8594 , \IDinst/n8593 , \IDinst/n8592 ,
         \IDinst/n8591 , \IDinst/n8590 , \IDinst/n8589 , \IDinst/n8588 ,
         \IDinst/n8587 , \IDinst/n8586 , \IDinst/n8585 , \IDinst/n8584 ,
         \IDinst/n8583 , \IDinst/n8582 , \IDinst/n8581 , \IDinst/n8580 ,
         \IDinst/n8579 , \IDinst/n8578 , \IDinst/n8577 , \IDinst/n8576 ,
         \IDinst/n8575 , \IDinst/n8574 , \IDinst/n8573 , \IDinst/n8572 ,
         \IDinst/n8571 , \IDinst/n8570 , \IDinst/n8569 , \IDinst/n8568 ,
         \IDinst/n8567 , \IDinst/n8566 , \IDinst/n8565 , \IDinst/n8564 ,
         \IDinst/n8563 , \IDinst/n8562 , \IDinst/n8561 , \IDinst/n8560 ,
         \IDinst/n8559 , \IDinst/n8558 , \IDinst/n8557 , \IDinst/n8556 ,
         \IDinst/n8555 , \IDinst/n8554 , \IDinst/n8553 , \IDinst/n8552 ,
         \IDinst/n8551 , \IDinst/n8550 , \IDinst/n8549 , \IDinst/n8548 ,
         \IDinst/n8547 , \IDinst/n8546 , \IDinst/n8545 , \IDinst/n8544 ,
         \IDinst/n8543 , \IDinst/n8542 , \IDinst/n8541 , \IDinst/n8540 ,
         \IDinst/n8539 , \IDinst/n8538 , \IDinst/n8537 , \IDinst/n8536 ,
         \IDinst/n8535 , \IDinst/n8534 , \IDinst/n8533 , \IDinst/n8532 ,
         \IDinst/n8531 , \IDinst/n8530 , \IDinst/n8529 , \IDinst/n8528 ,
         \IDinst/n8527 , \IDinst/n8526 , \IDinst/n8525 , \IDinst/n8524 ,
         \IDinst/n8523 , \IDinst/n8522 , \IDinst/n8521 , \IDinst/n8520 ,
         \IDinst/n8519 , \IDinst/n8518 , \IDinst/n8517 , \IDinst/n8516 ,
         \IDinst/n8515 , \IDinst/n8514 , \IDinst/n8513 , \IDinst/n8512 ,
         \IDinst/n8511 , \IDinst/n8510 , \IDinst/n8509 , \IDinst/n8508 ,
         \IDinst/n8507 , \IDinst/n8506 , \IDinst/n8505 , \IDinst/n8504 ,
         \IDinst/n8503 , \IDinst/n8502 , \IDinst/n8501 , \IDinst/n8500 ,
         \IDinst/n8499 , \IDinst/n8498 , \IDinst/n8497 , \IDinst/n8496 ,
         \IDinst/n8495 , \IDinst/n8494 , \IDinst/n8493 , \IDinst/n8492 ,
         \IDinst/n8491 , \IDinst/n8490 , \IDinst/n8489 , \IDinst/n8488 ,
         \IDinst/n8487 , \IDinst/n8486 , \IDinst/n8485 , \IDinst/n8484 ,
         \IDinst/n8483 , \IDinst/n8482 , \IDinst/n8481 , \IDinst/n8480 ,
         \IDinst/n8479 , \IDinst/n8478 , \IDinst/n8477 , \IDinst/n8476 ,
         \IDinst/n8475 , \IDinst/n8474 , \IDinst/n8473 , \IDinst/n8472 ,
         \IDinst/n8471 , \IDinst/n8470 , \IDinst/n8469 , \IDinst/n8468 ,
         \IDinst/n8467 , \IDinst/n8466 , \IDinst/n8465 , \IDinst/n8464 ,
         \IDinst/n8463 , \IDinst/n8462 , \IDinst/n8461 , \IDinst/n8460 ,
         \IDinst/n8459 , \IDinst/n8458 , \IDinst/n8457 , \IDinst/n8456 ,
         \IDinst/n8455 , \IDinst/n8454 , \IDinst/n8453 , \IDinst/n8452 ,
         \IDinst/n8451 , \IDinst/n8450 , \IDinst/n8449 , \IDinst/n8448 ,
         \IDinst/n8447 , \IDinst/n8446 , \IDinst/n8445 , \IDinst/n8444 ,
         \IDinst/n8443 , \IDinst/n8442 , \IDinst/n8441 , \IDinst/n8440 ,
         \IDinst/n8439 , \IDinst/n8438 , \IDinst/n8437 , \IDinst/n8436 ,
         \IDinst/n8435 , \IDinst/n8434 , \IDinst/n8433 , \IDinst/n8432 ,
         \IDinst/n8431 , \IDinst/n8430 , \IDinst/n8429 , \IDinst/n8428 ,
         \IDinst/n8427 , \IDinst/n8426 , \IDinst/n8425 , \IDinst/n8424 ,
         \IDinst/n8423 , \IDinst/n8422 , \IDinst/n8421 , \IDinst/n8420 ,
         \IDinst/n8419 , \IDinst/n8418 , \IDinst/n8417 , \IDinst/n8416 ,
         \IDinst/n8415 , \IDinst/n8414 , \IDinst/n8413 , \IDinst/n8412 ,
         \IDinst/n8411 , \IDinst/n8410 , \IDinst/n8409 , \IDinst/n8408 ,
         \IDinst/n8407 , \IDinst/n8406 , \IDinst/n8405 , \IDinst/n8404 ,
         \IDinst/n8403 , \IDinst/n8402 , \IDinst/n8401 , \IDinst/n8400 ,
         \IDinst/n8399 , \IDinst/n8398 , \IDinst/n8397 , \IDinst/n8396 ,
         \IDinst/n8395 , \IDinst/n8394 , \IDinst/n8393 , \IDinst/n8392 ,
         \IDinst/n8391 , \IDinst/n8390 , \IDinst/n8389 , \IDinst/n8388 ,
         \IDinst/n8387 , \IDinst/n8386 , \IDinst/n8385 , \IDinst/n8384 ,
         \IDinst/n8383 , \IDinst/n8382 , \IDinst/n8381 , \IDinst/n8380 ,
         \IDinst/n8379 , \IDinst/n8378 , \IDinst/n8377 , \IDinst/n8376 ,
         \IDinst/n8375 , \IDinst/n8374 , \IDinst/n8373 , \IDinst/n8372 ,
         \IDinst/n8371 , \IDinst/n8370 , \IDinst/n8369 , \IDinst/n8368 ,
         \IDinst/n8367 , \IDinst/n8366 , \IDinst/n8365 , \IDinst/n8364 ,
         \IDinst/n8363 , \IDinst/n8362 , \IDinst/n8361 , \IDinst/n8360 ,
         \IDinst/n8359 , \IDinst/n8358 , \IDinst/n8357 , \IDinst/n8356 ,
         \IDinst/n8355 , \IDinst/n8354 , \IDinst/n8353 , \IDinst/n8352 ,
         \IDinst/n8351 , \IDinst/n8350 , \IDinst/n8349 , \IDinst/n8348 ,
         \IDinst/n8347 , \IDinst/n8346 , \IDinst/n8345 , \IDinst/n8344 ,
         \IDinst/n8343 , \IDinst/n8342 , \IDinst/n8341 , \IDinst/n8340 ,
         \IDinst/n8339 , \IDinst/n8338 , \IDinst/n8337 , \IDinst/n8336 ,
         \IDinst/n8335 , \IDinst/n8334 , \IDinst/n8333 , \IDinst/n8332 ,
         \IDinst/n8331 , \IDinst/n8330 , \IDinst/n8329 , \IDinst/n8328 ,
         \IDinst/n8327 , \IDinst/n8326 , \IDinst/n8325 , \IDinst/n8324 ,
         \IDinst/n8323 , \IDinst/n8322 , \IDinst/n8321 , \IDinst/n8320 ,
         \IDinst/n8319 , \IDinst/n8318 , \IDinst/n8317 , \IDinst/n8316 ,
         \IDinst/n8315 , \IDinst/n8314 , \IDinst/n8313 , \IDinst/n8312 ,
         \IDinst/n8311 , \IDinst/n8310 , \IDinst/n8309 , \IDinst/n8308 ,
         \IDinst/n8307 , \IDinst/n8306 , \IDinst/n8305 , \IDinst/n8304 ,
         \IDinst/n8303 , \IDinst/n8302 , \IDinst/n8301 , \IDinst/n8300 ,
         \IDinst/n8299 , \IDinst/n8298 , \IDinst/n8297 , \IDinst/n8296 ,
         \IDinst/n8295 , \IDinst/n8294 , \IDinst/n8293 , \IDinst/n8292 ,
         \IDinst/n8291 , \IDinst/n8290 , \IDinst/n8289 , \IDinst/n8288 ,
         \IDinst/n8287 , \IDinst/n8286 , \IDinst/n8285 , \IDinst/n8284 ,
         \IDinst/n8283 , \IDinst/n8282 , \IDinst/n8281 , \IDinst/n8280 ,
         \IDinst/n8279 , \IDinst/n8278 , \IDinst/n8277 , \IDinst/n8276 ,
         \IDinst/n8275 , \IDinst/n8274 , \IDinst/n8273 , \IDinst/n8272 ,
         \IDinst/n8271 , \IDinst/n8270 , \IDinst/n8269 , \IDinst/n8268 ,
         \IDinst/n8267 , \IDinst/n8266 , \IDinst/n8265 , \IDinst/n8264 ,
         \IDinst/n8263 , \IDinst/n8262 , \IDinst/n8261 , \IDinst/n8260 ,
         \IDinst/n8259 , \IDinst/n8258 , \IDinst/n8257 , \IDinst/n8256 ,
         \IDinst/n8255 , \IDinst/n8254 , \IDinst/n8253 , \IDinst/n8252 ,
         \IDinst/n8251 , \IDinst/n8250 , \IDinst/n8249 , \IDinst/n8248 ,
         \IDinst/n8247 , \IDinst/n8246 , \IDinst/n8245 , \IDinst/n8244 ,
         \IDinst/n8243 , \IDinst/n8242 , \IDinst/n8241 , \IDinst/n8240 ,
         \IDinst/n8239 , \IDinst/n8238 , \IDinst/n8237 , \IDinst/n8236 ,
         \IDinst/n8235 , \IDinst/n8234 , \IDinst/n8233 , \IDinst/n8232 ,
         \IDinst/n8231 , \IDinst/n8230 , \IDinst/n8229 , \IDinst/n8228 ,
         \IDinst/n8227 , \IDinst/n8226 , \IDinst/n8225 , \IDinst/n8224 ,
         \IDinst/n8223 , \IDinst/n8222 , \IDinst/n8221 , \IDinst/n8220 ,
         \IDinst/n8219 , \IDinst/n8218 , \IDinst/n8217 , \IDinst/n8216 ,
         \IDinst/n8215 , \IDinst/n8214 , \IDinst/n8213 , \IDinst/n8212 ,
         \IDinst/n8211 , \IDinst/n8210 , \IDinst/n8209 , \IDinst/n8208 ,
         \IDinst/n8207 , \IDinst/n8206 , \IDinst/n8205 , \IDinst/n8204 ,
         \IDinst/n8203 , \IDinst/n8202 , \IDinst/n8201 , \IDinst/n8200 ,
         \IDinst/n8199 , \IDinst/n8198 , \IDinst/n8197 , \IDinst/n8196 ,
         \IDinst/n8195 , \IDinst/n8194 , \IDinst/n8193 , \IDinst/n8192 ,
         \IDinst/n8191 , \IDinst/n8190 , \IDinst/n8189 , \IDinst/n8188 ,
         \IDinst/n8187 , \IDinst/n8186 , \IDinst/n8185 , \IDinst/n8184 ,
         \IDinst/n8183 , \IDinst/n8182 , \IDinst/n8181 , \IDinst/n8180 ,
         \IDinst/n8179 , \IDinst/n8178 , \IDinst/n8177 , \IDinst/n8176 ,
         \IDinst/n8175 , \IDinst/n8174 , \IDinst/n8173 , \IDinst/n8172 ,
         \IDinst/n8171 , \IDinst/n8170 , \IDinst/n8169 , \IDinst/n8168 ,
         \IDinst/n8167 , \IDinst/n8166 , \IDinst/n8165 , \IDinst/n8164 ,
         \IDinst/n8163 , \IDinst/n8162 , \IDinst/n8161 , \IDinst/n8160 ,
         \IDinst/n8159 , \IDinst/n8158 , \IDinst/n8157 , \IDinst/n8156 ,
         \IDinst/n8155 , \IDinst/n8154 , \IDinst/n8153 , \IDinst/n8152 ,
         \IDinst/n8151 , \IDinst/n8150 , \IDinst/n8149 , \IDinst/n8148 ,
         \IDinst/n8147 , \IDinst/n8146 , \IDinst/n8145 , \IDinst/n8144 ,
         \IDinst/n8143 , \IDinst/n8142 , \IDinst/n8141 , \IDinst/n8140 ,
         \IDinst/n8139 , \IDinst/n8138 , \IDinst/n8137 , \IDinst/n8136 ,
         \IDinst/n8135 , \IDinst/n8134 , \IDinst/n8133 , \IDinst/n8132 ,
         \IDinst/n8131 , \IDinst/n8130 , \IDinst/n8129 , \IDinst/n8128 ,
         \IDinst/n8127 , \IDinst/n8126 , \IDinst/n8125 , \IDinst/n8124 ,
         \IDinst/n8123 , \IDinst/n8122 , \IDinst/n8121 , \IDinst/n8120 ,
         \IDinst/n8119 , \IDinst/n8118 , \IDinst/n8117 , \IDinst/n8116 ,
         \IDinst/n8115 , \IDinst/n8114 , \IDinst/n8113 , \IDinst/n8112 ,
         \IDinst/n8111 , \IDinst/n8110 , \IDinst/n8109 , \IDinst/n8108 ,
         \IDinst/n8107 , \IDinst/n8106 , \IDinst/n8105 , \IDinst/n8104 ,
         \IDinst/n8103 , \IDinst/n8102 , \IDinst/n8101 , \IDinst/n8100 ,
         \IDinst/n8099 , \IDinst/n8098 , \IDinst/n8097 , \IDinst/n8096 ,
         \IDinst/n8095 , \IDinst/n8094 , \IDinst/n8093 , \IDinst/n8092 ,
         \IDinst/n8091 , \IDinst/n8090 , \IDinst/n8089 , \IDinst/n8088 ,
         \IDinst/n8087 , \IDinst/n8086 , \IDinst/n8085 , \IDinst/n8084 ,
         \IDinst/n8083 , \IDinst/n8082 , \IDinst/n8081 , \IDinst/n8080 ,
         \IDinst/n8079 , \IDinst/n8078 , \IDinst/n8077 , \IDinst/n8076 ,
         \IDinst/n8075 , \IDinst/n8074 , \IDinst/n8073 , \IDinst/n8072 ,
         \IDinst/n8071 , \IDinst/n8070 , \IDinst/n8069 , \IDinst/n8068 ,
         \IDinst/n8067 , \IDinst/n8066 , \IDinst/n8065 , \IDinst/n8064 ,
         \IDinst/n8063 , \IDinst/n8062 , \IDinst/n8061 , \IDinst/n8060 ,
         \IDinst/n8059 , \IDinst/n8058 , \IDinst/n8057 , \IDinst/n8056 ,
         \IDinst/n8055 , \IDinst/n8054 , \IDinst/n8053 , \IDinst/n8052 ,
         \IDinst/n8051 , \IDinst/n8050 , \IDinst/n8049 , \IDinst/n8048 ,
         \IDinst/n8047 , \IDinst/n8046 , \IDinst/n8045 , \IDinst/n8044 ,
         \IDinst/n8043 , \IDinst/n8042 , \IDinst/n8041 , \IDinst/n8040 ,
         \IDinst/n8039 , \IDinst/n8038 , \IDinst/n8037 , \IDinst/n8036 ,
         \IDinst/n8035 , \IDinst/n8034 , \IDinst/n8033 , \IDinst/n8032 ,
         \IDinst/n8031 , \IDinst/n8030 , \IDinst/n8029 , \IDinst/n8028 ,
         \IDinst/n8027 , \IDinst/n8026 , \IDinst/n8025 , \IDinst/n8024 ,
         \IDinst/n8023 , \IDinst/n8022 , \IDinst/n8021 , \IDinst/n8020 ,
         \IDinst/n8019 , \IDinst/n8018 , \IDinst/n8017 , \IDinst/n8016 ,
         \IDinst/n8015 , \IDinst/n8014 , \IDinst/n8013 , \IDinst/n8012 ,
         \IDinst/n8011 , \IDinst/n8010 , \IDinst/n8009 , \IDinst/n8008 ,
         \IDinst/n8007 , \IDinst/n8006 , \IDinst/n8005 , \IDinst/n8004 ,
         \IDinst/n8003 , \IDinst/n8002 , \IDinst/n8001 , \IDinst/n8000 ,
         \IDinst/n7999 , \IDinst/n7998 , \IDinst/n7997 , \IDinst/n7996 ,
         \IDinst/n7995 , \IDinst/n7994 , \IDinst/n7993 , \IDinst/n7992 ,
         \IDinst/n7991 , \IDinst/n7990 , \IDinst/n7989 , \IDinst/n7988 ,
         \IDinst/n7987 , \IDinst/n7986 , \IDinst/n7985 , \IDinst/n7984 ,
         \IDinst/n7983 , \IDinst/n7982 , \IDinst/n7981 , \IDinst/n7980 ,
         \IDinst/n7979 , \IDinst/n7978 , \IDinst/n7977 , \IDinst/n7976 ,
         \IDinst/n7975 , \IDinst/n7974 , \IDinst/n7973 , \IDinst/n7972 ,
         \IDinst/n7971 , \IDinst/n7970 , \IDinst/n7969 , \IDinst/n7968 ,
         \IDinst/n7967 , \IDinst/n7966 , \IDinst/n7965 , \IDinst/n7964 ,
         \IDinst/n7963 , \IDinst/n7962 , \IDinst/n7961 , \IDinst/n7960 ,
         \IDinst/n7959 , \IDinst/n7958 , \IDinst/n7957 , \IDinst/n7956 ,
         \IDinst/n7955 , \IDinst/n7954 , \IDinst/n7953 , \IDinst/n7952 ,
         \IDinst/n7951 , \IDinst/n7950 , \IDinst/n7949 , \IDinst/n7948 ,
         \IDinst/n7947 , \IDinst/n7946 , \IDinst/n7945 , \IDinst/n7944 ,
         \IDinst/n7943 , \IDinst/n7942 , \IDinst/n7941 , \IDinst/n7940 ,
         \IDinst/n7939 , \IDinst/n7938 , \IDinst/n7937 , \IDinst/n7936 ,
         \IDinst/n7935 , \IDinst/n7934 , \IDinst/n7933 , \IDinst/n7932 ,
         \IDinst/n7931 , \IDinst/n7930 , \IDinst/n7929 , \IDinst/n7928 ,
         \IDinst/n7927 , \IDinst/n7926 , \IDinst/n7925 , \IDinst/n7924 ,
         \IDinst/n7923 , \IDinst/n7922 , \IDinst/n7921 , \IDinst/n7920 ,
         \IDinst/n7919 , \IDinst/n7918 , \IDinst/n7917 , \IDinst/n7916 ,
         \IDinst/n7915 , \IDinst/n7914 , \IDinst/n7913 , \IDinst/n7912 ,
         \IDinst/n7911 , \IDinst/n7910 , \IDinst/n7909 , \IDinst/n7908 ,
         \IDinst/n7907 , \IDinst/n7906 , \IDinst/n7905 , \IDinst/n7904 ,
         \IDinst/n7903 , \IDinst/n7902 , \IDinst/n7901 , \IDinst/n7900 ,
         \IDinst/n7899 , \IDinst/n7898 , \IDinst/n7897 , \IDinst/n7896 ,
         \IDinst/n7895 , \IDinst/n7894 , \IDinst/n7893 , \IDinst/n7892 ,
         \IDinst/n7891 , \IDinst/n7890 , \IDinst/n7889 , \IDinst/n7888 ,
         \IDinst/n7887 , \IDinst/n7886 , \IDinst/n7885 , \IDinst/n7884 ,
         \IDinst/n7883 , \IDinst/n7882 , \IDinst/n7881 , \IDinst/n7880 ,
         \IDinst/n7879 , \IDinst/n7878 , \IDinst/n7877 , \IDinst/n7876 ,
         \IDinst/n7875 , \IDinst/n7874 , \IDinst/n7873 , \IDinst/n7872 ,
         \IDinst/n7871 , \IDinst/n7870 , \IDinst/n7869 , \IDinst/n7868 ,
         \IDinst/n7867 , \IDinst/n7866 , \IDinst/n7865 , \IDinst/n7864 ,
         \IDinst/n7863 , \IDinst/n7862 , \IDinst/n7861 , \IDinst/n7860 ,
         \IDinst/n7859 , \IDinst/n7858 , \IDinst/n7857 , \IDinst/n7856 ,
         \IDinst/n7855 , \IDinst/n7854 , \IDinst/n7853 , \IDinst/n7852 ,
         \IDinst/n7851 , \IDinst/n7850 , \IDinst/n7849 , \IDinst/n7848 ,
         \IDinst/n7847 , \IDinst/n7846 , \IDinst/n7845 , \IDinst/n7844 ,
         \IDinst/n7843 , \IDinst/n7842 , \IDinst/n7841 , \IDinst/n7840 ,
         \IDinst/n7839 , \IDinst/n7838 , \IDinst/n7837 , \IDinst/n7836 ,
         \IDinst/n7835 , \IDinst/n7834 , \IDinst/n7833 , \IDinst/n7832 ,
         \IDinst/n7831 , \IDinst/n7830 , \IDinst/n7829 , \IDinst/n7828 ,
         \IDinst/n7827 , \IDinst/n7826 , \IDinst/n7825 , \IDinst/n7824 ,
         \IDinst/n7823 , \IDinst/n7822 , \IDinst/n7821 , \IDinst/n7820 ,
         \IDinst/n7819 , \IDinst/n7818 , \IDinst/n7817 , \IDinst/n7816 ,
         \IDinst/n7815 , \IDinst/n7814 , \IDinst/n7813 , \IDinst/n7812 ,
         \IDinst/n7811 , \IDinst/n7810 , \IDinst/n7809 , \IDinst/n7808 ,
         \IDinst/n7807 , \IDinst/n7806 , \IDinst/n7805 , \IDinst/n7804 ,
         \IDinst/n7803 , \IDinst/n7802 , \IDinst/n7801 , \IDinst/n7800 ,
         \IDinst/n7799 , \IDinst/n7798 , \IDinst/n7797 , \IDinst/n7796 ,
         \IDinst/n7795 , \IDinst/n7794 , \IDinst/n7793 , \IDinst/n7792 ,
         \IDinst/n7791 , \IDinst/n7790 , \IDinst/n7789 , \IDinst/n7788 ,
         \IDinst/n7787 , \IDinst/n7786 , \IDinst/n7785 , \IDinst/n7784 ,
         \IDinst/n7783 , \IDinst/n7782 , \IDinst/n7781 , \IDinst/n7780 ,
         \IDinst/n7779 , \IDinst/n7778 , \IDinst/n7777 , \IDinst/n7776 ,
         \IDinst/n7775 , \IDinst/n7774 , \IDinst/n7773 , \IDinst/n7772 ,
         \IDinst/n7771 , \IDinst/n7770 , \IDinst/n7769 , \IDinst/n7768 ,
         \IDinst/n7767 , \IDinst/n7766 , \IDinst/n7765 , \IDinst/n7764 ,
         \IDinst/n7763 , \IDinst/n7762 , \IDinst/n7761 , \IDinst/n7760 ,
         \IDinst/n7759 , \IDinst/n7758 , \IDinst/n7757 , \IDinst/n7756 ,
         \IDinst/n7755 , \IDinst/n7754 , \IDinst/n7753 , \IDinst/n7752 ,
         \IDinst/n7751 , \IDinst/n7750 , \IDinst/n7749 , \IDinst/n7748 ,
         \IDinst/n7747 , \IDinst/n7746 , \IDinst/n7745 , \IDinst/n7744 ,
         \IDinst/n7743 , \IDinst/n7742 , \IDinst/n7741 , \IDinst/n7740 ,
         \IDinst/n7739 , \IDinst/n7738 , \IDinst/n7737 , \IDinst/n7736 ,
         \IDinst/n7735 , \IDinst/n7734 , \IDinst/n7733 , \IDinst/n7732 ,
         \IDinst/n7731 , \IDinst/n7730 , \IDinst/n7729 , \IDinst/n7728 ,
         \IDinst/n7727 , \IDinst/n7726 , \IDinst/n7725 , \IDinst/n7724 ,
         \IDinst/n7723 , \IDinst/n7722 , \IDinst/n7721 , \IDinst/n7720 ,
         \IDinst/n7719 , \IDinst/n7718 , \IDinst/n7717 , \IDinst/n7716 ,
         \IDinst/n7715 , \IDinst/n7714 , \IDinst/n7713 , \IDinst/n7712 ,
         \IDinst/n7711 , \IDinst/n7710 , \IDinst/n7709 , \IDinst/n7708 ,
         \IDinst/n7707 , \IDinst/n7706 , \IDinst/n7705 , \IDinst/n7704 ,
         \IDinst/n7703 , \IDinst/n7702 , \IDinst/n7701 , \IDinst/n7700 ,
         \IDinst/n7699 , \IDinst/n7698 , \IDinst/n7697 , \IDinst/n7696 ,
         \IDinst/n7695 , \IDinst/n7694 , \IDinst/n7693 , \IDinst/n7692 ,
         \IDinst/n7691 , \IDinst/n7690 , \IDinst/n7689 , \IDinst/n7688 ,
         \IDinst/n7687 , \IDinst/n7686 , \IDinst/n7685 , \IDinst/n7684 ,
         \IDinst/n7683 , \IDinst/n7682 , \IDinst/n7681 , \IDinst/n7680 ,
         \IDinst/n7679 , \IDinst/n7678 , \IDinst/n7677 , \IDinst/n7676 ,
         \IDinst/n7675 , \IDinst/n7674 , \IDinst/n7673 , \IDinst/n7672 ,
         \IDinst/n7671 , \IDinst/n7670 , \IDinst/n7669 , \IDinst/n7668 ,
         \IDinst/n7667 , \IDinst/n7666 , \IDinst/n7665 , \IDinst/n7664 ,
         \IDinst/n7663 , \IDinst/n7662 , \IDinst/n7661 , \IDinst/n7660 ,
         \IDinst/n7659 , \IDinst/n7658 , \IDinst/n7657 , \IDinst/n7656 ,
         \IDinst/n7655 , \IDinst/n7654 , \IDinst/n7653 , \IDinst/n7652 ,
         \IDinst/n7651 , \IDinst/n7650 , \IDinst/n7649 , \IDinst/n7648 ,
         \IDinst/n7647 , \IDinst/n7646 , \IDinst/n7645 , \IDinst/n7644 ,
         \IDinst/n7643 , \IDinst/n7642 , \IDinst/n7641 , \IDinst/n7640 ,
         \IDinst/n7639 , \IDinst/n7638 , \IDinst/n7637 , \IDinst/n7636 ,
         \IDinst/n7635 , \IDinst/n7634 , \IDinst/n7633 , \IDinst/n7632 ,
         \IDinst/n7631 , \IDinst/n7630 , \IDinst/n7629 , \IDinst/n7628 ,
         \IDinst/n7627 , \IDinst/n7626 , \IDinst/n7625 , \IDinst/n7624 ,
         \IDinst/n7623 , \IDinst/n7622 , \IDinst/n7621 , \IDinst/n7620 ,
         \IDinst/n7619 , \IDinst/n7618 , \IDinst/n7617 , \IDinst/n7616 ,
         \IDinst/n7615 , \IDinst/n7614 , \IDinst/n7613 , \IDinst/n7612 ,
         \IDinst/n7611 , \IDinst/n7610 , \IDinst/n7609 , \IDinst/n7608 ,
         \IDinst/n7607 , \IDinst/n7606 , \IDinst/n7605 , \IDinst/n7604 ,
         \IDinst/n7603 , \IDinst/n7602 , \IDinst/n7601 , \IDinst/n7600 ,
         \IDinst/n7599 , \IDinst/n7598 , \IDinst/n7597 , \IDinst/n7596 ,
         \IDinst/n7595 , \IDinst/n7594 , \IDinst/n7593 , \IDinst/n7592 ,
         \IDinst/n7591 , \IDinst/n7590 , \IDinst/n7589 , \IDinst/n7588 ,
         \IDinst/n7587 , \IDinst/n7586 , \IDinst/n7585 , \IDinst/n7584 ,
         \IDinst/n7583 , \IDinst/n7582 , \IDinst/n7581 , \IDinst/n7580 ,
         \IDinst/n7579 , \IDinst/n7578 , \IDinst/n7577 , \IDinst/n7576 ,
         \IDinst/n7575 , \IDinst/n7574 , \IDinst/n7573 , \IDinst/n7572 ,
         \IDinst/n7571 , \IDinst/n7570 , \IDinst/n7569 , \IDinst/n7568 ,
         \IDinst/n7567 , \IDinst/n7566 , \IDinst/n7565 , \IDinst/n7564 ,
         \IDinst/n7563 , \IDinst/n7562 , \IDinst/n7561 , \IDinst/n7560 ,
         \IDinst/n7559 , \IDinst/n7558 , \IDinst/n7557 , \IDinst/n7556 ,
         \IDinst/n7555 , \IDinst/n7554 , \IDinst/n7553 , \IDinst/n7552 ,
         \IDinst/n7551 , \IDinst/n7550 , \IDinst/n7549 , \IDinst/n7548 ,
         \IDinst/n7547 , \IDinst/n7546 , \IDinst/n7545 , \IDinst/n7544 ,
         \IDinst/n7543 , \IDinst/n7542 , \IDinst/n7541 , \IDinst/n7540 ,
         \IDinst/n7539 , \IDinst/n7538 , \IDinst/n7537 , \IDinst/n7536 ,
         \IDinst/n7535 , \IDinst/n7534 , \IDinst/n7533 , \IDinst/n7532 ,
         \IDinst/n7531 , \IDinst/n7530 , \IDinst/n7529 , \IDinst/n7528 ,
         \IDinst/n7527 , \IDinst/n7526 , \IDinst/n7525 , \IDinst/n7524 ,
         \IDinst/n7523 , \IDinst/n7522 , \IDinst/n7521 , \IDinst/n7520 ,
         \IDinst/n7519 , \IDinst/n7518 , \IDinst/n7517 , \IDinst/n7516 ,
         \IDinst/n7515 , \IDinst/n7514 , \IDinst/n7513 , \IDinst/n7512 ,
         \IDinst/n7511 , \IDinst/n7510 , \IDinst/n7509 , \IDinst/n7508 ,
         \IDinst/n7507 , \IDinst/n7506 , \IDinst/n7505 , \IDinst/n7504 ,
         \IDinst/n7503 , \IDinst/n7502 , \IDinst/n7501 , \IDinst/n7500 ,
         \IDinst/n7499 , \IDinst/n7498 , \IDinst/n7497 , \IDinst/n7496 ,
         \IDinst/n7495 , \IDinst/n7494 , \IDinst/n7493 , \IDinst/n7492 ,
         \IDinst/n7491 , \IDinst/n7490 , \IDinst/n7489 , \IDinst/n7488 ,
         \IDinst/n7487 , \IDinst/n7486 , \IDinst/n7485 , \IDinst/n7484 ,
         \IDinst/n7483 , \IDinst/n7482 , \IDinst/n7481 , \IDinst/n7480 ,
         \IDinst/n7479 , \IDinst/n7478 , \IDinst/n7477 , \IDinst/n7476 ,
         \IDinst/n7475 , \IDinst/n7474 , \IDinst/n7473 , \IDinst/n7472 ,
         \IDinst/n7471 , \IDinst/n7470 , \IDinst/n7469 , \IDinst/n7468 ,
         \IDinst/n7467 , \IDinst/n7466 , \IDinst/n7465 , \IDinst/n7464 ,
         \IDinst/n7463 , \IDinst/n7462 , \IDinst/n7461 , \IDinst/n7460 ,
         \IDinst/n7459 , \IDinst/n7458 , \IDinst/n7457 , \IDinst/n7456 ,
         \IDinst/n7455 , \IDinst/n7454 , \IDinst/n7453 , \IDinst/n7452 ,
         \IDinst/n7451 , \IDinst/n7450 , \IDinst/n7449 , \IDinst/n7448 ,
         \IDinst/n7447 , \IDinst/n7446 , \IDinst/n7445 , \IDinst/n7444 ,
         \IDinst/n7443 , \IDinst/n7442 , \IDinst/n7441 , \IDinst/n7440 ,
         \IDinst/n7439 , \IDinst/n7438 , \IDinst/n7437 , \IDinst/n7436 ,
         \IDinst/n7435 , \IDinst/n7434 , \IDinst/n7433 , \IDinst/n7432 ,
         \IDinst/n7431 , \IDinst/n7430 , \IDinst/n7429 , \IDinst/n7428 ,
         \IDinst/n7427 , \IDinst/n7426 , \IDinst/n7425 , \IDinst/n7424 ,
         \IDinst/n7423 , \IDinst/n7422 , \IDinst/n7421 , \IDinst/n7420 ,
         \IDinst/n7419 , \IDinst/n7418 , \IDinst/n7417 , \IDinst/n7416 ,
         \IDinst/n7415 , \IDinst/n7414 , \IDinst/n7413 , \IDinst/n7412 ,
         \IDinst/n7411 , \IDinst/n7410 , \IDinst/n7409 , \IDinst/n7408 ,
         \IDinst/n7407 , \IDinst/n7406 , \IDinst/n7405 , \IDinst/n7404 ,
         \IDinst/n7403 , \IDinst/n7402 , \IDinst/n7401 , \IDinst/n7400 ,
         \IDinst/n7399 , \IDinst/n7398 , \IDinst/n7397 , \IDinst/n7396 ,
         \IDinst/n7395 , \IDinst/n7394 , \IDinst/n7393 , \IDinst/n7392 ,
         \IDinst/n7391 , \IDinst/n7390 , \IDinst/n7389 , \IDinst/n7388 ,
         \IDinst/n7387 , \IDinst/n7386 , \IDinst/n7385 , \IDinst/n7384 ,
         \IDinst/n7383 , \IDinst/n7382 , \IDinst/n7381 , \IDinst/n7380 ,
         \IDinst/n7379 , \IDinst/n7378 , \IDinst/n7377 , \IDinst/n7376 ,
         \IDinst/n7375 , \IDinst/n7374 , \IDinst/n7373 , \IDinst/n7372 ,
         \IDinst/n7371 , \IDinst/n7370 , \IDinst/n7369 , \IDinst/n7368 ,
         \IDinst/n7367 , \IDinst/n7366 , \IDinst/n7365 , \IDinst/n7364 ,
         \IDinst/n7363 , \IDinst/n7362 , \IDinst/n7361 , \IDinst/n7360 ,
         \IDinst/n7359 , \IDinst/n7358 , \IDinst/n7357 , \IDinst/n7356 ,
         \IDinst/n7355 , \IDinst/n7354 , \IDinst/n7353 , \IDinst/n7352 ,
         \IDinst/n7351 , \IDinst/n7350 , \IDinst/n7349 , \IDinst/n7348 ,
         \IDinst/n7347 , \IDinst/n7346 , \IDinst/n7345 , \IDinst/n7344 ,
         \IDinst/n7343 , \IDinst/n7342 , \IDinst/n7341 , \IDinst/n7340 ,
         \IDinst/n7339 , \IDinst/n7338 , \IDinst/n7337 , \IDinst/n7336 ,
         \IDinst/n7335 , \IDinst/n7334 , \IDinst/n7333 , \IDinst/n7332 ,
         \IDinst/n7331 , \IDinst/n7330 , \IDinst/n7329 , \IDinst/n7328 ,
         \IDinst/n7327 , \IDinst/n7326 , \IDinst/n7325 , \IDinst/n7324 ,
         \IDinst/n7323 , \IDinst/n7322 , \IDinst/n7321 , \IDinst/n7320 ,
         \IDinst/n7319 , \IDinst/n7318 , \IDinst/n7317 , \IDinst/n7316 ,
         \IDinst/n7315 , \IDinst/n7314 , \IDinst/n7313 , \IDinst/n7312 ,
         \IDinst/n7311 , \IDinst/n7310 , \IDinst/n7309 , \IDinst/n7308 ,
         \IDinst/n7307 , \IDinst/n7306 , \IDinst/n7305 , \IDinst/n7304 ,
         \IDinst/n7303 , \IDinst/n7302 , \IDinst/n7301 , \IDinst/n7300 ,
         \IDinst/n7299 , \IDinst/n7298 , \IDinst/n7297 , \IDinst/n7296 ,
         \IDinst/n7295 , \IDinst/n7294 , \IDinst/n7293 , \IDinst/n7292 ,
         \IDinst/n7291 , \IDinst/n7290 , \IDinst/n7289 , \IDinst/n7288 ,
         \IDinst/n7287 , \IDinst/n7286 , \IDinst/n7285 , \IDinst/n7284 ,
         \IDinst/n7283 , \IDinst/n7282 , \IDinst/n7281 , \IDinst/n7280 ,
         \IDinst/n7279 , \IDinst/n7278 , \IDinst/n7277 , \IDinst/n7276 ,
         \IDinst/n7275 , \IDinst/n7274 , \IDinst/n7273 , \IDinst/n7272 ,
         \IDinst/n7271 , \IDinst/n7270 , \IDinst/n7269 , \IDinst/n7268 ,
         \IDinst/n7267 , \IDinst/n7266 , \IDinst/n7265 , \IDinst/n7264 ,
         \IDinst/n7263 , \IDinst/n7262 , \IDinst/n7261 , \IDinst/n7260 ,
         \IDinst/n7259 , \IDinst/n7258 , \IDinst/n7257 , \IDinst/n7256 ,
         \IDinst/n7255 , \IDinst/n7254 , \IDinst/n7253 , \IDinst/n7252 ,
         \IDinst/n7251 , \IDinst/n7250 , \IDinst/n7249 , \IDinst/n7248 ,
         \IDinst/n7247 , \IDinst/n7246 , \IDinst/n7245 , \IDinst/n7244 ,
         \IDinst/n7243 , \IDinst/n7242 , \IDinst/n7241 , \IDinst/n7240 ,
         \IDinst/n7239 , \IDinst/n7238 , \IDinst/n7237 , \IDinst/n7236 ,
         \IDinst/n7235 , \IDinst/n7234 , \IDinst/n7233 , \IDinst/n7232 ,
         \IDinst/n7231 , \IDinst/n7230 , \IDinst/n7229 , \IDinst/n7228 ,
         \IDinst/n7227 , \IDinst/n7226 , \IDinst/n7225 , \IDinst/n7224 ,
         \IDinst/n7223 , \IDinst/n7222 , \IDinst/n7221 , \IDinst/n7220 ,
         \IDinst/n7219 , \IDinst/n7218 , \IDinst/n7217 , \IDinst/n7216 ,
         \IDinst/n7215 , \IDinst/n7214 , \IDinst/n7213 , \IDinst/n7212 ,
         \IDinst/n7211 , \IDinst/n7210 , \IDinst/n7209 , \IDinst/n7208 ,
         \IDinst/n7207 , \IDinst/n7206 , \IDinst/n7205 , \IDinst/n7204 ,
         \IDinst/n7203 , \IDinst/n7202 , \IDinst/n7201 , \IDinst/n7200 ,
         \IDinst/n7199 , \IDinst/n7198 , \IDinst/n7197 , \IDinst/n7196 ,
         \IDinst/n7195 , \IDinst/n7194 , \IDinst/n7193 , \IDinst/n7192 ,
         \IDinst/n7191 , \IDinst/n7190 , \IDinst/n7189 , \IDinst/n7188 ,
         \IDinst/n7187 , \IDinst/n7186 , \IDinst/n7185 , \IDinst/n7184 ,
         \IDinst/n7183 , \IDinst/n7182 , \IDinst/n7181 , \IDinst/n7180 ,
         \IDinst/n7179 , \IDinst/n7178 , \IDinst/n7177 , \IDinst/n7176 ,
         \IDinst/n7175 , \IDinst/n7174 , \IDinst/n7173 , \IDinst/n7172 ,
         \IDinst/n7171 , \IDinst/n7170 , \IDinst/n7169 , \IDinst/n7168 ,
         \IDinst/n7167 , \IDinst/n7166 , \IDinst/n7165 , \IDinst/n7164 ,
         \IDinst/n7163 , \IDinst/n7162 , \IDinst/n7161 , \IDinst/n7160 ,
         \IDinst/n7159 , \IDinst/n7158 , \IDinst/n7157 , \IDinst/n7156 ,
         \IDinst/n7155 , \IDinst/n7154 , \IDinst/n7153 , \IDinst/n7152 ,
         \IDinst/n7151 , \IDinst/n7150 , \IDinst/n7149 , \IDinst/n7148 ,
         \IDinst/n7147 , \IDinst/n7146 , \IDinst/n7145 , \IDinst/n7144 ,
         \IDinst/n7143 , \IDinst/n7142 , \IDinst/n7141 , \IDinst/n7140 ,
         \IDinst/n7139 , \IDinst/n7138 , \IDinst/n7137 , \IDinst/n7136 ,
         \IDinst/n7135 , \IDinst/n7134 , \IDinst/n7133 , \IDinst/n7132 ,
         \IDinst/n7131 , \IDinst/n7130 , \IDinst/n7129 , \IDinst/n7128 ,
         \IDinst/n7127 , \IDinst/n7126 , \IDinst/n7125 , \IDinst/n7124 ,
         \IDinst/n7123 , \IDinst/n7122 , \IDinst/n7121 , \IDinst/n7120 ,
         \IDinst/n7119 , \IDinst/n7118 , \IDinst/n7117 , \IDinst/n7116 ,
         \IDinst/n7115 , \IDinst/n7114 , \IDinst/n7113 , \IDinst/n7112 ,
         \IDinst/n7111 , \IDinst/n7110 , \IDinst/n7109 , \IDinst/n7108 ,
         \IDinst/n7107 , \IDinst/n7106 , \IDinst/n7105 , \IDinst/n7104 ,
         \IDinst/n7103 , \IDinst/n7102 , \IDinst/n7101 , \IDinst/n7100 ,
         \IDinst/n7099 , \IDinst/n7098 , \IDinst/n7097 , \IDinst/n7096 ,
         \IDinst/n7095 , \IDinst/n7094 , \IDinst/n7093 , \IDinst/n7092 ,
         \IDinst/n7091 , \IDinst/n7090 , \IDinst/n7089 , \IDinst/n7088 ,
         \IDinst/n7087 , \IDinst/n7086 , \IDinst/n7085 , \IDinst/n7084 ,
         \IDinst/n7083 , \IDinst/n7082 , \IDinst/n7081 , \IDinst/n7080 ,
         \IDinst/n7079 , \IDinst/n7078 , \IDinst/n7077 , \IDinst/n7076 ,
         \IDinst/n7075 , \IDinst/n7074 , \IDinst/n7073 , \IDinst/n7072 ,
         \IDinst/n7071 , \IDinst/n7070 , \IDinst/n7069 , \IDinst/n7068 ,
         \IDinst/n7067 , \IDinst/n7066 , \IDinst/n7065 , \IDinst/n7064 ,
         \IDinst/n7063 , \IDinst/n7062 , \IDinst/n7061 , \IDinst/n7060 ,
         \IDinst/n7059 , \IDinst/n7058 , \IDinst/n7057 , \IDinst/n7056 ,
         \IDinst/n7055 , \IDinst/n7054 , \IDinst/n7053 , \IDinst/n7052 ,
         \IDinst/n7051 , \IDinst/n7050 , \IDinst/n7049 , \IDinst/n7048 ,
         \IDinst/n7047 , \IDinst/n7046 , \IDinst/n7045 , \IDinst/n7044 ,
         \IDinst/n7043 , \IDinst/n7042 , \IDinst/n7041 , \IDinst/n7040 ,
         \IDinst/n7039 , \IDinst/n7038 , \IDinst/n7037 , \IDinst/n7036 ,
         \IDinst/n7035 , \IDinst/n7034 , \IDinst/n7033 , \IDinst/n7032 ,
         \IDinst/n7031 , \IDinst/n7030 , \IDinst/n7029 , \IDinst/n7028 ,
         \IDinst/n7027 , \IDinst/n7026 , \IDinst/n7025 , \IDinst/n7024 ,
         \IDinst/n7023 , \IDinst/n7022 , \IDinst/n7021 , \IDinst/n7020 ,
         \IDinst/n7019 , \IDinst/n7018 , \IDinst/n7017 , \IDinst/n7016 ,
         \IDinst/n7015 , \IDinst/n7014 , \IDinst/n7013 , \IDinst/n7012 ,
         \IDinst/n7011 , \IDinst/n7010 , \IDinst/n7009 , \IDinst/n7008 ,
         \IDinst/n7007 , \IDinst/n7006 , \IDinst/n7005 , \IDinst/n7004 ,
         \IDinst/n7003 , \IDinst/n7002 , \IDinst/n7001 , \IDinst/n7000 ,
         \IDinst/n6999 , \IDinst/n6998 , \IDinst/n6997 , \IDinst/n6996 ,
         \IDinst/n6995 , \IDinst/n6994 , \IDinst/n6993 , \IDinst/n6992 ,
         \IDinst/n6991 , \IDinst/n6990 , \IDinst/n6989 , \IDinst/n6988 ,
         \IDinst/n6987 , \IDinst/n6986 , \IDinst/n6985 , \IDinst/n6984 ,
         \IDinst/n6983 , \IDinst/n6982 , \IDinst/n6981 , \IDinst/n6980 ,
         \IDinst/n6979 , \IDinst/n6978 , \IDinst/n6977 , \IDinst/n6976 ,
         \IDinst/n6975 , \IDinst/n6974 , \IDinst/n6973 , \IDinst/n6972 ,
         \IDinst/n6971 , \IDinst/n6970 , \IDinst/n6969 , \IDinst/n6968 ,
         \IDinst/n6967 , \IDinst/n6966 , \IDinst/n6965 , \IDinst/n6964 ,
         \IDinst/n6963 , \IDinst/n6962 , \IDinst/n6961 , \IDinst/n6960 ,
         \IDinst/n6959 , \IDinst/n6958 , \IDinst/n6957 , \IDinst/n6956 ,
         \IDinst/n6955 , \IDinst/n6954 , \IDinst/n6953 , \IDinst/n6952 ,
         \IDinst/n6951 , \IDinst/n6950 , \IDinst/n6949 , \IDinst/n6948 ,
         \IDinst/n6947 , \IDinst/n6946 , \IDinst/n6945 , \IDinst/n6944 ,
         \IDinst/n6943 , \IDinst/n6942 , \IDinst/n6941 , \IDinst/n6940 ,
         \IDinst/n6939 , \IDinst/n6938 , \IDinst/n6937 , \IDinst/n6936 ,
         \IDinst/n6935 , \IDinst/n6934 , \IDinst/n6933 , \IDinst/n6932 ,
         \IDinst/n6931 , \IDinst/n6930 , \IDinst/n6929 , \IDinst/n6928 ,
         \IDinst/n6927 , \IDinst/n6926 , \IDinst/n6925 , \IDinst/n6924 ,
         \IDinst/n6923 , \IDinst/n6922 , \IDinst/n6921 , \IDinst/n6920 ,
         \IDinst/n6919 , \IDinst/n6918 , \IDinst/n6917 , \IDinst/n6916 ,
         \IDinst/n6915 , \IDinst/n6914 , \IDinst/n6913 , \IDinst/n6912 ,
         \IDinst/n6911 , \IDinst/n6910 , \IDinst/n6909 , \IDinst/n6908 ,
         \IDinst/n6907 , \IDinst/n6906 , \IDinst/n6905 , \IDinst/n6904 ,
         \IDinst/n6903 , \IDinst/n6902 , \IDinst/n6901 , \IDinst/n6900 ,
         \IDinst/n6899 , \IDinst/n6898 , \IDinst/n6897 , \IDinst/n6896 ,
         \IDinst/n6895 , \IDinst/n6894 , \IDinst/n6893 , \IDinst/n6892 ,
         \IDinst/n6891 , \IDinst/n6890 , \IDinst/n6889 , \IDinst/n6888 ,
         \IDinst/n6887 , \IDinst/n6886 , \IDinst/n6885 , \IDinst/n6884 ,
         \IDinst/n6883 , \IDinst/n6882 , \IDinst/n6881 , \IDinst/n6880 ,
         \IDinst/n6879 , \IDinst/n6878 , \IDinst/n6877 , \IDinst/n6876 ,
         \IDinst/n6875 , \IDinst/n6874 , \IDinst/n6873 , \IDinst/n6872 ,
         \IDinst/n6871 , \IDinst/n6870 , \IDinst/n6869 , \IDinst/n6868 ,
         \IDinst/n6867 , \IDinst/n6866 , \IDinst/n6865 , \IDinst/n6864 ,
         \IDinst/n6863 , \IDinst/n6862 , \IDinst/n6861 , \IDinst/n6860 ,
         \IDinst/n6859 , \IDinst/n6858 , \IDinst/n6857 , \IDinst/n6856 ,
         \IDinst/n6855 , \IDinst/n6854 , \IDinst/n6853 , \IDinst/n6852 ,
         \IDinst/n6851 , \IDinst/n6850 , \IDinst/n6849 , \IDinst/n6848 ,
         \IDinst/n6847 , \IDinst/n6846 , \IDinst/n6845 , \IDinst/n6844 ,
         \IDinst/n6843 , \IDinst/n6842 , \IDinst/n6841 , \IDinst/n6840 ,
         \IDinst/n6839 , \IDinst/n6838 , \IDinst/n6837 , \IDinst/n6836 ,
         \IDinst/n6835 , \IDinst/n6834 , \IDinst/n6833 , \IDinst/n6832 ,
         \IDinst/n6831 , \IDinst/n6830 , \IDinst/n6829 , \IDinst/n6828 ,
         \IDinst/n6827 , \IDinst/n6826 , \IDinst/n6825 , \IDinst/n6824 ,
         \IDinst/n6823 , \IDinst/n6822 , \IDinst/n6821 , \IDinst/n6820 ,
         \IDinst/n6819 , \IDinst/n6818 , \IDinst/n6817 , \IDinst/n6816 ,
         \IDinst/n6815 , \IDinst/n6814 , \IDinst/n6813 , \IDinst/n6812 ,
         \IDinst/n6811 , \IDinst/n6810 , \IDinst/n6809 , \IDinst/n6808 ,
         \IDinst/n6807 , \IDinst/n6806 , \IDinst/n6805 , \IDinst/n6804 ,
         \IDinst/n6803 , \IDinst/n6802 , \IDinst/n6801 , \IDinst/n6800 ,
         \IDinst/n6799 , \IDinst/n6798 , \IDinst/n6797 , \IDinst/n6796 ,
         \IDinst/n6795 , \IDinst/n6794 , \IDinst/n6793 , \IDinst/n6792 ,
         \IDinst/n6791 , \IDinst/n6790 , \IDinst/n6789 , \IDinst/n6788 ,
         \IDinst/n6787 , \IDinst/n6786 , \IDinst/n6785 , \IDinst/n6784 ,
         \IDinst/n6783 , \IDinst/n6782 , \IDinst/n6781 , \IDinst/n6780 ,
         \IDinst/n6779 , \IDinst/n6778 , \IDinst/n6777 , \IDinst/n6776 ,
         \IDinst/n6775 , \IDinst/n6774 , \IDinst/n6773 , \IDinst/n6772 ,
         \IDinst/n6771 , \IDinst/n6770 , \IDinst/n6769 , \IDinst/n6768 ,
         \IDinst/n6767 , \IDinst/n6766 , \IDinst/n6765 , \IDinst/n6764 ,
         \IDinst/n6763 , \IDinst/n6762 , \IDinst/n6761 , \IDinst/n6760 ,
         \IDinst/n6759 , \IDinst/n6758 , \IDinst/n6757 , \IDinst/n6756 ,
         \IDinst/n6755 , \IDinst/n6754 , \IDinst/n6753 , \IDinst/n6752 ,
         \IDinst/n6751 , \IDinst/n6750 , \IDinst/n6749 , \IDinst/n6748 ,
         \IDinst/n6747 , \IDinst/n6746 , \IDinst/n6745 , \IDinst/n6744 ,
         \IDinst/n6743 , \IDinst/n6742 , \IDinst/n6741 , \IDinst/n6740 ,
         \IDinst/n6739 , \IDinst/n6738 , \IDinst/n6737 , \IDinst/n6736 ,
         \IDinst/n6735 , \IDinst/n6734 , \IDinst/n6733 , \IDinst/n6732 ,
         \IDinst/n6731 , \IDinst/n6730 , \IDinst/n6729 , \IDinst/n6728 ,
         \IDinst/n6727 , \IDinst/n6726 , \IDinst/n6725 , \IDinst/n6724 ,
         \IDinst/n6723 , \IDinst/n6722 , \IDinst/n6721 , \IDinst/n6720 ,
         \IDinst/n6719 , \IDinst/n6718 , \IDinst/n6717 , \IDinst/n6716 ,
         \IDinst/n6715 , \IDinst/n6714 , \IDinst/n6713 , \IDinst/n6712 ,
         \IDinst/n6711 , \IDinst/n6710 , \IDinst/n6709 , \IDinst/n6708 ,
         \IDinst/n6707 , \IDinst/n6706 , \IDinst/n6705 , \IDinst/n6704 ,
         \IDinst/n6703 , \IDinst/n6702 , \IDinst/n6701 , \IDinst/n6700 ,
         \IDinst/n6699 , \IDinst/n6698 , \IDinst/n6697 , \IDinst/n6696 ,
         \IDinst/n6695 , \IDinst/n6694 , \IDinst/n6693 , \IDinst/n6692 ,
         \IDinst/n6691 , \IDinst/n6690 , \IDinst/n6689 , \IDinst/n6688 ,
         \IDinst/n6687 , \IDinst/n6686 , \IDinst/n6685 , \IDinst/n6684 ,
         \IDinst/n6683 , \IDinst/n6682 , \IDinst/n6681 , \IDinst/n6680 ,
         \IDinst/n6679 , \IDinst/n6678 , \IDinst/n6677 , \IDinst/n6676 ,
         \IDinst/n6675 , \IDinst/n6674 , \IDinst/n6673 , \IDinst/n6672 ,
         \IDinst/n6671 , \IDinst/n6670 , \IDinst/n6669 , \IDinst/n6668 ,
         \IDinst/n6667 , \IDinst/n6666 , \IDinst/n6665 , \IDinst/n6664 ,
         \IDinst/n6663 , \IDinst/n6662 , \IDinst/n6661 , \IDinst/n6660 ,
         \IDinst/n6659 , \IDinst/n6658 , \IDinst/n6657 , \IDinst/n6656 ,
         \IDinst/n6655 , \IDinst/n6654 , \IDinst/n6653 , \IDinst/n6652 ,
         \IDinst/n6651 , \IDinst/n6650 , \IDinst/n6649 , \IDinst/n6648 ,
         \IDinst/n6647 , \IDinst/n6646 , \IDinst/n6645 , \IDinst/n6644 ,
         \IDinst/n6643 , \IDinst/n6642 , \IDinst/n6641 , \IDinst/n6640 ,
         \IDinst/n6639 , \IDinst/n6638 , \IDinst/n6637 , \IDinst/n6636 ,
         \IDinst/n6635 , \IDinst/n6634 , \IDinst/n6633 , \IDinst/n6632 ,
         \IDinst/n6631 , \IDinst/n6630 , \IDinst/n6629 , \IDinst/n6628 ,
         \IDinst/n6627 , \IDinst/n6626 , \IDinst/n6625 , \IDinst/n6624 ,
         \IDinst/n6623 , \IDinst/n6622 , \IDinst/n6621 , \IDinst/n6620 ,
         \IDinst/n6619 , \IDinst/n6618 , \IDinst/n6617 , \IDinst/n6616 ,
         \IDinst/n6615 , \IDinst/n6614 , \IDinst/n6613 , \IDinst/n6612 ,
         \IDinst/n6611 , \IDinst/n6610 , \IDinst/n6609 , \IDinst/n6608 ,
         \IDinst/n6607 , \IDinst/n6606 , \IDinst/n6605 , \IDinst/n6604 ,
         \IDinst/n6603 , \IDinst/n6602 , \IDinst/n6601 , \IDinst/n6600 ,
         \IDinst/n6599 , \IDinst/n6598 , \IDinst/n6597 , \IDinst/n6596 ,
         \IDinst/n6595 , \IDinst/n6594 , \IDinst/n6593 , \IDinst/n6592 ,
         \IDinst/n6591 , \IDinst/n6590 , \IDinst/n6589 , \IDinst/n6588 ,
         \IDinst/n6587 , \IDinst/n6586 , \IDinst/n6585 , \IDinst/n6584 ,
         \IDinst/n6583 , \IDinst/n6582 , \IDinst/n6581 , \IDinst/n6580 ,
         \IDinst/n6579 , \IDinst/n6578 , \IDinst/n6577 , \IDinst/n6576 ,
         \IDinst/n6575 , \IDinst/n6574 , \IDinst/n6573 , \IDinst/n6572 ,
         \IDinst/n6571 , \IDinst/n6570 , \IDinst/n6569 , \IDinst/n6568 ,
         \IDinst/n6567 , \IDinst/n6566 , \IDinst/n6565 , \IDinst/n6564 ,
         \IDinst/n6563 , \IDinst/n6562 , \IDinst/n6561 , \IDinst/n6560 ,
         \IDinst/n6559 , \IDinst/n6558 , \IDinst/n6557 , \IDinst/n6556 ,
         \IDinst/n6555 , \IDinst/n6554 , \IDinst/n6553 , \IDinst/n6552 ,
         \IDinst/n6551 , \IDinst/n6550 , \IDinst/n6549 , \IDinst/n6548 ,
         \IDinst/n6547 , \IDinst/n6546 , \IDinst/n6545 , \IDinst/n6544 ,
         \IDinst/n6543 , \IDinst/n6542 , \IDinst/n6541 , \IDinst/n6540 ,
         \IDinst/n6539 , \IDinst/n6538 , \IDinst/n6537 , \IDinst/n6536 ,
         \IDinst/n6535 , \IDinst/n6534 , \IDinst/n6533 , \IDinst/n6532 ,
         \IDinst/n6531 , \IDinst/n6530 , \IDinst/n6529 , \IDinst/n6528 ,
         \IDinst/n6527 , \IDinst/n6526 , \IDinst/n6525 , \IDinst/n6524 ,
         \IDinst/n6523 , \IDinst/n6522 , \IDinst/n6521 , \IDinst/n6520 ,
         \IDinst/n6519 , \IDinst/n6518 , \IDinst/n6517 , \IDinst/n6516 ,
         \IDinst/n6515 , \IDinst/n6514 , \IDinst/n6513 , \IDinst/n6512 ,
         \IDinst/n6511 , \IDinst/n6510 , \IDinst/n6509 , \IDinst/n6508 ,
         \IDinst/n6507 , \IDinst/n6506 , \IDinst/n6505 , \IDinst/n6504 ,
         \IDinst/n6503 , \IDinst/n6502 , \IDinst/n6501 , \IDinst/n6500 ,
         \IDinst/n6499 , \IDinst/n6498 , \IDinst/n6497 , \IDinst/n6496 ,
         \IDinst/n6495 , \IDinst/n6494 , \IDinst/n6493 , \IDinst/n6492 ,
         \IDinst/n6491 , \IDinst/n6490 , \IDinst/n6489 , \IDinst/n6488 ,
         \IDinst/n6487 , \IDinst/n6486 , \IDinst/n6485 , \IDinst/n6484 ,
         \IDinst/n6483 , \IDinst/n6482 , \IDinst/n6481 , \IDinst/n6480 ,
         \IDinst/n6479 , \IDinst/n6478 , \IDinst/n6477 , \IDinst/n6476 ,
         \IDinst/n6475 , \IDinst/n6474 , \IDinst/n6473 , \IDinst/n6472 ,
         \IDinst/n6471 , \IDinst/n6470 , \IDinst/n6469 , \IDinst/n6468 ,
         \IDinst/n6467 , \IDinst/n6466 , \IDinst/n6465 , \IDinst/n6464 ,
         \IDinst/n6463 , \IDinst/n6462 , \IDinst/n6461 , \IDinst/n6460 ,
         \IDinst/n6459 , \IDinst/n6458 , \IDinst/n6457 , \IDinst/n6456 ,
         \IDinst/n6455 , \IDinst/n6454 , \IDinst/n6453 , \IDinst/n6452 ,
         \IDinst/n6451 , \IDinst/n6450 , \IDinst/n6449 , \IDinst/n6448 ,
         \IDinst/n6447 , \IDinst/n6446 , \IDinst/n6445 , \IDinst/n6444 ,
         \IDinst/n6443 , \IDinst/n6442 , \IDinst/n6441 , \IDinst/n6440 ,
         \IDinst/n6439 , \IDinst/n6438 , \IDinst/n6437 , \IDinst/n6436 ,
         \IDinst/n6435 , \IDinst/n6434 , \IDinst/n6433 , \IDinst/n6432 ,
         \IDinst/n6431 , \IDinst/n6430 , \IDinst/n6429 , \IDinst/n6428 ,
         \IDinst/n6427 , \IDinst/n6426 , \IDinst/n6425 , \IDinst/n6424 ,
         \IDinst/n6423 , \IDinst/n6422 , \IDinst/n6421 , \IDinst/n6420 ,
         \IDinst/n6419 , \IDinst/n6418 , \IDinst/n6417 , \IDinst/n6416 ,
         \IDinst/n6415 , \IDinst/n6414 , \IDinst/n6413 , \IDinst/n6412 ,
         \IDinst/n6411 , \IDinst/n6410 , \IDinst/n6409 , \IDinst/n6408 ,
         \IDinst/n6407 , \IDinst/n6406 , \IDinst/n6405 , \IDinst/n6404 ,
         \IDinst/n6403 , \IDinst/n6402 , \IDinst/n6401 , \IDinst/n6400 ,
         \IDinst/n6399 , \IDinst/n6398 , \IDinst/n6397 , \IDinst/n6396 ,
         \IDinst/n6395 , \IDinst/n6394 , \IDinst/n6393 , \IDinst/n6392 ,
         \IDinst/n6391 , \IDinst/n6390 , \IDinst/n6389 , \IDinst/n6388 ,
         \IDinst/n6387 , \IDinst/n6386 , \IDinst/n6385 , \IDinst/n6384 ,
         \IDinst/n6383 , \IDinst/n6382 , \IDinst/n6381 , \IDinst/n6380 ,
         \IDinst/n6379 , \IDinst/n6378 , \IDinst/n6377 , \IDinst/n6376 ,
         \IDinst/n6375 , \IDinst/n6374 , \IDinst/n6373 , \IDinst/n6372 ,
         \IDinst/n6371 , \IDinst/n6370 , \IDinst/n6369 , \IDinst/n6368 ,
         \IDinst/n6367 , \IDinst/n6366 , \IDinst/n6365 , \IDinst/n6364 ,
         \IDinst/n6363 , \IDinst/n6362 , \IDinst/n6361 , \IDinst/n6360 ,
         \IDinst/n6359 , \IDinst/n6358 , \IDinst/n6357 , \IDinst/n6356 ,
         \IDinst/n6355 , \IDinst/n6354 , \IDinst/n6353 , \IDinst/n6352 ,
         \IDinst/n6351 , \IDinst/n6350 , \IDinst/n6349 , \IDinst/n6348 ,
         \IDinst/n6347 , \IDinst/n6346 , \IDinst/n6345 , \IDinst/n6344 ,
         \IDinst/n6343 , \IDinst/n6342 , \IDinst/n6341 , \IDinst/n6340 ,
         \IDinst/n6339 , \IDinst/n6338 , \IDinst/n6337 , \IDinst/n6336 ,
         \IDinst/n6335 , \IDinst/n6334 , \IDinst/n6333 , \IDinst/n6332 ,
         \IDinst/n6331 , \IDinst/n6330 , \IDinst/n6329 , \IDinst/n6328 ,
         \IDinst/n6327 , \IDinst/n6326 , \IDinst/n6325 , \IDinst/n6324 ,
         \IDinst/n6323 , \IDinst/n6322 , \IDinst/n6321 , \IDinst/n6320 ,
         \IDinst/n6319 , \IDinst/n6318 , \IDinst/n6317 , \IDinst/n6316 ,
         \IDinst/n6315 , \IDinst/n6314 , \IDinst/n6313 , \IDinst/n6312 ,
         \IDinst/n6311 , \IDinst/n6310 , \IDinst/n6309 , \IDinst/n6308 ,
         \IDinst/n6307 , \IDinst/n6306 , \IDinst/n6305 , \IDinst/n6304 ,
         \IDinst/n6303 , \IDinst/n6302 , \IDinst/n6301 , \IDinst/n6300 ,
         \IDinst/n6299 , \IDinst/n6298 , \IDinst/n6297 , \IDinst/n6296 ,
         \IDinst/n6295 , \IDinst/n6294 , \IDinst/n6293 , \IDinst/n6292 ,
         \IDinst/n6291 , \IDinst/n6290 , \IDinst/n6289 , \IDinst/n6288 ,
         \IDinst/n6287 , \IDinst/n6286 , \IDinst/n6285 , \IDinst/n6284 ,
         \IDinst/n6283 , \IDinst/n6282 , \IDinst/n6281 , \IDinst/n6280 ,
         \IDinst/n6279 , \IDinst/n6278 , \IDinst/n6277 , \IDinst/n6276 ,
         \IDinst/n6275 , \IDinst/n6274 , \IDinst/n6273 , \IDinst/n6272 ,
         \IDinst/n6271 , \IDinst/n6270 , \IDinst/n6269 , \IDinst/n6268 ,
         \IDinst/n6267 , \IDinst/n6266 , \IDinst/n6265 , \IDinst/n6264 ,
         \IDinst/n6263 , \IDinst/n6262 , \IDinst/n6261 , \IDinst/n6260 ,
         \IDinst/n6259 , \IDinst/n6258 , \IDinst/n6257 , \IDinst/n6256 ,
         \IDinst/n6255 , \IDinst/n6254 , \IDinst/n6253 , \IDinst/n6252 ,
         \IDinst/n6251 , \IDinst/n6250 , \IDinst/n6249 , \IDinst/n6248 ,
         \IDinst/n6247 , \IDinst/n6246 , \IDinst/n6245 , \IDinst/n6244 ,
         \IDinst/n6243 , \IDinst/n6242 , \IDinst/n6241 , \IDinst/n6240 ,
         \IDinst/n6239 , \IDinst/n6238 , \IDinst/n6237 , \IDinst/n6236 ,
         \IDinst/n6235 , \IDinst/n6234 , \IDinst/n6233 , \IDinst/n6232 ,
         \IDinst/n6231 , \IDinst/n6230 , \IDinst/n6229 , \IDinst/n6228 ,
         \IDinst/n6227 , \IDinst/n6226 , \IDinst/n6225 , \IDinst/n6224 ,
         \IDinst/n6223 , \IDinst/n6222 , \IDinst/n6221 , \IDinst/n6220 ,
         \IDinst/n6219 , \IDinst/n6218 , \IDinst/n6217 , \IDinst/n6216 ,
         \IDinst/n6215 , \IDinst/n6214 , \IDinst/n6213 , \IDinst/n6212 ,
         \IDinst/n6211 , \IDinst/n6210 , \IDinst/n6209 , \IDinst/n6208 ,
         \IDinst/n6207 , \IDinst/n6206 , \IDinst/n6205 , \IDinst/n6204 ,
         \IDinst/n6203 , \IDinst/n6202 , \IDinst/n6201 , \IDinst/n6200 ,
         \IDinst/n6199 , \IDinst/n6198 , \IDinst/n6197 , \IDinst/n6196 ,
         \IDinst/n6195 , \IDinst/n6194 , \IDinst/n6193 , \IDinst/n6192 ,
         \IDinst/n6191 , \IDinst/n6190 , \IDinst/n6189 , \IDinst/n6188 ,
         \IDinst/n6187 , \IDinst/n6186 , \IDinst/n6185 , \IDinst/n6184 ,
         \IDinst/n6183 , \IDinst/n6182 , \IDinst/n6181 , \IDinst/n6180 ,
         \IDinst/n6179 , \IDinst/n6178 , \IDinst/n6177 , \IDinst/n6176 ,
         \IDinst/n6175 , \IDinst/n6174 , \IDinst/n6173 , \IDinst/n6172 ,
         \IDinst/n6171 , \IDinst/n6170 , \IDinst/n6169 , \IDinst/n6168 ,
         \IDinst/n6167 , \IDinst/n6166 , \IDinst/n6165 , \IDinst/n6164 ,
         \IDinst/n6163 , \IDinst/n6162 , \IDinst/n6161 , \IDinst/n6160 ,
         \IDinst/n6159 , \IDinst/n6158 , \IDinst/n6157 , \IDinst/n6156 ,
         \IDinst/n6155 , \IDinst/n6154 , \IDinst/n6153 , \IDinst/n6152 ,
         \IDinst/n6151 , \IDinst/n6150 , \IDinst/n6149 , \IDinst/n6148 ,
         \IDinst/n6147 , \IDinst/n6146 , \IDinst/n6145 , \IDinst/n6144 ,
         \IDinst/n6143 , \IDinst/n6142 , \IDinst/n6141 , \IDinst/n6140 ,
         \IDinst/n6139 , \IDinst/n6138 , \IDinst/n6137 , \IDinst/n6136 ,
         \IDinst/n6135 , \IDinst/n6134 , \IDinst/n6133 , \IDinst/n6132 ,
         \IDinst/n6131 , \IDinst/n6130 , \IDinst/n6129 , \IDinst/n6128 ,
         \IDinst/n6127 , \IDinst/n6126 , \IDinst/n6125 , \IDinst/n6124 ,
         \IDinst/n6123 , \IDinst/n6122 , \IDinst/n6121 , \IDinst/n6120 ,
         \IDinst/n6119 , \IDinst/n6118 , \IDinst/n6117 , \IDinst/n6116 ,
         \IDinst/n6115 , \IDinst/n6114 , \IDinst/n6113 , \IDinst/n6112 ,
         \IDinst/n6111 , \IDinst/n6110 , \IDinst/n6109 , \IDinst/n6108 ,
         \IDinst/n6107 , \IDinst/n6106 , \IDinst/n6105 , \IDinst/n6104 ,
         \IDinst/n6103 , \IDinst/n6102 , \IDinst/n6101 , \IDinst/n6100 ,
         \IDinst/n6099 , \IDinst/n6098 , \IDinst/n6097 , \IDinst/n6096 ,
         \IDinst/n6095 , \IDinst/n6094 , \IDinst/n6093 , \IDinst/n6092 ,
         \IDinst/n6091 , \IDinst/n6090 , \IDinst/n6089 , \IDinst/n6088 ,
         \IDinst/n6087 , \IDinst/n6086 , \IDinst/n6085 , \IDinst/n6084 ,
         \IDinst/n6083 , \IDinst/n6082 , \IDinst/n6081 , \IDinst/n6080 ,
         \IDinst/n6079 , \IDinst/n6078 , \IDinst/n6077 , \IDinst/n6076 ,
         \IDinst/n6075 , \IDinst/n6074 , \IDinst/n6073 , \IDinst/n6072 ,
         \IDinst/n6071 , \IDinst/n6070 , \IDinst/n6069 , \IDinst/n6068 ,
         \IDinst/n6067 , \IDinst/n6066 , \IDinst/n6065 , \IDinst/n6064 ,
         \IDinst/n6063 , \IDinst/n6062 , \IDinst/n6061 , \IDinst/n6060 ,
         \IDinst/n6059 , \IDinst/n6058 , \IDinst/n6057 , \IDinst/n6056 ,
         \IDinst/n6055 , \IDinst/n6054 , \IDinst/n6053 , \IDinst/n6052 ,
         \IDinst/n6051 , \IDinst/n6050 , \IDinst/n6049 , \IDinst/n6048 ,
         \IDinst/n6047 , \IDinst/n6046 , \IDinst/n6045 , \IDinst/n6044 ,
         \IDinst/n6043 , \IDinst/n6042 , \IDinst/n6041 , \IDinst/n6040 ,
         \IDinst/n6039 , \IDinst/n6038 , \IDinst/n6037 , \IDinst/n6036 ,
         \IDinst/n6035 , \IDinst/n6034 , \IDinst/n6033 , \IDinst/n6032 ,
         \IDinst/n6031 , \IDinst/n6030 , \IDinst/n6029 , \IDinst/n6028 ,
         \IDinst/n6027 , \IDinst/n6026 , \IDinst/n6025 , \IDinst/n6024 ,
         \IDinst/n6023 , \IDinst/n6022 , \IDinst/n6021 , \IDinst/n6020 ,
         \IDinst/n6019 , \IDinst/n6018 , \IDinst/n6017 , \IDinst/n6016 ,
         \IDinst/n6015 , \IDinst/n6014 , \IDinst/n6013 , \IDinst/n6012 ,
         \IDinst/n6011 , \IDinst/n6010 , \IDinst/n6009 , \IDinst/n6008 ,
         \IDinst/n6007 , \IDinst/n6006 , \IDinst/n6005 , \IDinst/n6004 ,
         \IDinst/n6003 , \IDinst/n6002 , \IDinst/n6001 , \IDinst/n6000 ,
         \IDinst/n5999 , \IDinst/n5998 , \IDinst/n5997 , \IDinst/n5996 ,
         \IDinst/n5995 , \IDinst/n5994 , \IDinst/n5993 , \IDinst/n5992 ,
         \IDinst/n5991 , \IDinst/n5990 , \IDinst/n5989 , \IDinst/n5988 ,
         \IDinst/n5987 , \IDinst/n5986 , \IDinst/n5985 , \IDinst/n5984 ,
         \IDinst/n5983 , \IDinst/n5982 , \IDinst/n5981 , \IDinst/n5980 ,
         \IDinst/n5979 , \IDinst/n5978 , \IDinst/n5977 , \IDinst/n5976 ,
         \IDinst/n5975 , \IDinst/n5974 , \IDinst/n5973 , \IDinst/n5972 ,
         \IDinst/n5971 , \IDinst/n5970 , \IDinst/n5969 , \IDinst/n5968 ,
         \IDinst/n5967 , \IDinst/n5966 , \IDinst/n5965 , \IDinst/n5964 ,
         \IDinst/n5963 , \IDinst/n5962 , \IDinst/n5961 , \IDinst/n5960 ,
         \IDinst/n5959 , \IDinst/n5958 , \IDinst/n5957 , \IDinst/n5956 ,
         \IDinst/n5955 , \IDinst/n5954 , \IDinst/n5953 , \IDinst/n5952 ,
         \IDinst/n5951 , \IDinst/n5950 , \IDinst/n5949 , \IDinst/n5948 ,
         \IDinst/n5947 , \IDinst/n5946 , \IDinst/n5945 , \IDinst/n5944 ,
         \IDinst/n5943 , \IDinst/n5926 , \IDinst/n5925 , \IDinst/n5924 ,
         \IDinst/n5923 , \IDinst/n5922 , \IDinst/n5921 , \IDinst/n5920 ,
         \IDinst/n5919 , \IDinst/n5918 , \IDinst/n5917 , \IDinst/n5916 ,
         \IDinst/n5915 , \IDinst/n5914 , \IDinst/n5913 , \IDinst/n5912 ,
         \IDinst/n5911 , \IDinst/n5910 , \IDinst/n5909 , \IDinst/n5908 ,
         \IDinst/n5907 , \IDinst/n5906 , \IDinst/n5905 , \IDinst/n5904 ,
         \IDinst/n5903 , \IDinst/n5902 , \IDinst/n5901 , \IDinst/n5900 ,
         \IDinst/n5899 , \IDinst/n5898 , \IDinst/n5897 , \IDinst/n5896 ,
         \IDinst/n5895 , \IDinst/n5894 , \IDinst/n5893 , \IDinst/n5892 ,
         \IDinst/n5891 , \IDinst/n5890 , \IDinst/n5889 , \IDinst/n5888 ,
         \IDinst/n5887 , \IDinst/n5886 , \IDinst/n5885 , \IDinst/n5884 ,
         \IDinst/n5883 , \IDinst/n5882 , \IDinst/n5881 , \IDinst/n5880 ,
         \IDinst/n5879 , \IDinst/n5878 , \IDinst/n5877 , \IDinst/n5876 ,
         \IDinst/n5875 , \IDinst/n5874 , \IDinst/n5873 , \IDinst/n5872 ,
         \IDinst/n5871 , \IDinst/n5870 , \IDinst/n5869 , \IDinst/n5868 ,
         \IDinst/n5867 , \IDinst/n5866 , \IDinst/n5865 , \IDinst/n5864 ,
         \IDinst/n5863 , \IDinst/n5862 , \IDinst/n5861 , \IDinst/n5860 ,
         \IDinst/n5859 , \IDinst/n5858 , \IDinst/n5857 , \IDinst/n5856 ,
         \IDinst/n5855 , \IDinst/n5854 , \IDinst/n5853 , \IDinst/n5852 ,
         \IDinst/n5851 , \IDinst/n5850 , \IDinst/n5849 , \IDinst/n5848 ,
         \IDinst/n5847 , \IDinst/n5846 , \IDinst/n5845 , \IDinst/n5844 ,
         \IDinst/n5843 , \IDinst/n5842 , \IDinst/n5841 , \IDinst/n5840 ,
         \IDinst/n5839 , \IDinst/n5838 , \IDinst/n5837 , \IDinst/n5836 ,
         \IDinst/n5835 , \IDinst/n5834 , \IDinst/n5833 , \IDinst/n5832 ,
         \IDinst/n5831 , \IDinst/n5830 , \IDinst/n5829 , \IDinst/n5828 ,
         \IDinst/n5827 , \IDinst/n5826 , \IDinst/n5825 , \IDinst/n5824 ,
         \IDinst/n5823 , \IDinst/n5822 , \IDinst/n5821 , \IDinst/n5820 ,
         \IDinst/n5819 , \IDinst/n5818 , \IDinst/n5817 , \IDinst/n5816 ,
         \IDinst/n5815 , \IDinst/n5814 , \IDinst/n5813 , \IDinst/n5812 ,
         \IDinst/n5811 , \IDinst/n5810 , \IDinst/n5809 , \IDinst/n5808 ,
         \IDinst/n5807 , \IDinst/n5806 , \IDinst/n5805 , \IDinst/n5804 ,
         \IDinst/n5803 , \IDinst/n5802 , \IDinst/n5801 , \IDinst/n5800 ,
         \IDinst/n5799 , \IDinst/n5798 , \IDinst/n5797 , \IDinst/n5796 ,
         \IDinst/n5795 , \IDinst/n5794 , \IDinst/n5793 , \IDinst/n5792 ,
         \IDinst/n5791 , \IDinst/n5790 , \IDinst/n5789 , \IDinst/n5788 ,
         \IDinst/n5787 , \IDinst/n5786 , \IDinst/n5785 , \IDinst/n5784 ,
         \IDinst/n5783 , \IDinst/n5782 , \IDinst/n5781 , \IDinst/n5780 ,
         \IDinst/n5779 , \IDinst/n5778 , \IDinst/n5777 , \IDinst/n5776 ,
         \IDinst/n5775 , \IDinst/n5774 , \IDinst/n5773 , \IDinst/n5772 ,
         \IDinst/n5771 , \IDinst/n5770 , \IDinst/n5769 , \IDinst/n5768 ,
         \IDinst/n5767 , \IDinst/n5766 , \IDinst/n5765 , \IDinst/n5764 ,
         \IDinst/n5763 , \IDinst/n5762 , \IDinst/n5761 , \IDinst/n5760 ,
         \IDinst/n5759 , \IDinst/n5758 , \IDinst/n5757 , \IDinst/n5756 ,
         \IDinst/n5755 , \IDinst/n5754 , \IDinst/n5753 , \IDinst/n5752 ,
         \IDinst/n5751 , \IDinst/n5750 , \IDinst/n5749 , \IDinst/n5748 ,
         \IDinst/n5747 , \IDinst/n5746 , \IDinst/n5745 , \IDinst/n5744 ,
         \IDinst/n5743 , \IDinst/n5742 , \IDinst/n5741 , \IDinst/n5740 ,
         \IDinst/n5739 , \IDinst/n5738 , \IDinst/n5737 , \IDinst/n5736 ,
         \IDinst/n5735 , \IDinst/n5734 , \IDinst/n5733 , \IDinst/n5732 ,
         \IDinst/n5731 , \IDinst/n5730 , \IDinst/n5729 , \IDinst/n5728 ,
         \IDinst/n5727 , \IDinst/n5726 , \IDinst/n5725 , \IDinst/n5724 ,
         \IDinst/n5723 , \IDinst/n5722 , \IDinst/n5721 , \IDinst/n5720 ,
         \IDinst/n5719 , \IDinst/n5718 , \IDinst/n5717 , \IDinst/n5716 ,
         \IDinst/n5715 , \IDinst/n5714 , \IDinst/n5713 , \IDinst/n5712 ,
         \IDinst/n5711 , \IDinst/n5710 , \IDinst/n5709 , \IDinst/n5708 ,
         \IDinst/n5707 , \IDinst/n5706 , \IDinst/n5705 , \IDinst/n5704 ,
         \IDinst/n5703 , \IDinst/n5702 , \IDinst/n5701 , \IDinst/n5700 ,
         \IDinst/n5699 , \IDinst/n5698 , \IDinst/n5697 , \IDinst/n5696 ,
         \IDinst/n5695 , \IDinst/n5694 , \IDinst/n5693 , \IDinst/n5692 ,
         \IDinst/n5691 , \IDinst/n5690 , \IDinst/n5689 , \IDinst/n5688 ,
         \IDinst/n5687 , \IDinst/n5686 , \IDinst/n5685 , \IDinst/n5684 ,
         \IDinst/n5683 , \IDinst/n5682 , \IDinst/n5681 , \IDinst/n5680 ,
         \IDinst/n5679 , \IDinst/n5678 , \IDinst/n5677 , \IDinst/n5676 ,
         \IDinst/n5675 , \IDinst/n5674 , \IDinst/n5673 , \IDinst/n5672 ,
         \IDinst/n5671 , \IDinst/n5670 , \IDinst/n5669 , \IDinst/n5668 ,
         \IDinst/n5667 , \IDinst/n5666 , \IDinst/n5665 , \IDinst/n5664 ,
         \IDinst/n5663 , \IDinst/n5662 , \IDinst/n5661 , \IDinst/n5660 ,
         \IDinst/n5659 , \IDinst/n5658 , \IDinst/n5657 , \IDinst/n5656 ,
         \IDinst/n5655 , \IDinst/n5654 , \IDinst/n5653 , \IDinst/n5652 ,
         \IDinst/n5651 , \IDinst/n5650 , \IDinst/n5649 , \IDinst/n5648 ,
         \IDinst/n5647 , \IDinst/n5646 , \IDinst/n5645 , \IDinst/n5644 ,
         \IDinst/n5643 , \IDinst/n5642 , \IDinst/n5641 , \IDinst/n5640 ,
         \IDinst/n5639 , \IDinst/n5638 , \IDinst/n5637 , \IDinst/n5636 ,
         \IDinst/n5635 , \IDinst/n5634 , \IDinst/n5633 , \IDinst/n5632 ,
         \IDinst/n5631 , \IDinst/n5630 , \IDinst/n5629 , \IDinst/n5628 ,
         \IDinst/n5627 , \IDinst/n5626 , \IDinst/n5625 , \IDinst/n5624 ,
         \IDinst/n5623 , \IDinst/n5622 , \IDinst/n5621 , \IDinst/n5620 ,
         \IDinst/n5619 , \IDinst/n5618 , \IDinst/n5617 , \IDinst/n5616 ,
         \IDinst/n5615 , \IDinst/n5614 , \IDinst/n5613 , \IDinst/n5612 ,
         \IDinst/n5611 , \IDinst/n5610 , \IDinst/n5609 , \IDinst/n5608 ,
         \IDinst/n5607 , \IDinst/n5606 , \IDinst/n5605 , \IDinst/n5604 ,
         \IDinst/n5603 , \IDinst/n5602 , \IDinst/n5601 , \IDinst/n5600 ,
         \IDinst/n5599 , \IDinst/n5598 , \IDinst/n5597 , \IDinst/n5596 ,
         \IDinst/n5595 , \IDinst/n5594 , \IDinst/n5593 , \IDinst/n5592 ,
         \IDinst/n5591 , \IDinst/n5590 , \IDinst/n5589 , \IDinst/n5588 ,
         \IDinst/n5587 , \IDinst/n5586 , \IDinst/n5585 , \IDinst/n5584 ,
         \IDinst/n5583 , \IDinst/n5582 , \IDinst/n5581 , \IDinst/n5580 ,
         \IDinst/n5579 , \IDinst/n5578 , \IDinst/n5577 , \IDinst/n5576 ,
         \IDinst/n5575 , \IDinst/n5574 , \IDinst/n5573 , \IDinst/n5572 ,
         \IDinst/n5571 , \IDinst/n5570 , \IDinst/n5569 , \IDinst/n5568 ,
         \IDinst/n5567 , \IDinst/n5566 , \IDinst/n5565 , \IDinst/n5564 ,
         \IDinst/n5563 , \IDinst/n5562 , \IDinst/n5561 , \IDinst/n5560 ,
         \IDinst/n5559 , \IDinst/n5558 , \IDinst/n5557 , \IDinst/n5556 ,
         \IDinst/n5555 , \IDinst/n5554 , \IDinst/n5553 , \IDinst/n5552 ,
         \IDinst/n5551 , \IDinst/n5550 , \IDinst/n5549 , \IDinst/n5548 ,
         \IDinst/n5547 , \IDinst/n5546 , \IDinst/n5545 , \IDinst/n5544 ,
         \IDinst/n5543 , \IDinst/n5542 , \IDinst/n5541 , \IDinst/n5540 ,
         \IDinst/n5539 , \IDinst/n5538 , \IDinst/n5537 , \IDinst/n5536 ,
         \IDinst/n5535 , \IDinst/n5534 , \IDinst/n5533 , \IDinst/n5532 ,
         \IDinst/n5531 , \IDinst/n5530 , \IDinst/n5529 , \IDinst/n5528 ,
         \IDinst/n5527 , \IDinst/n5526 , \IDinst/n5525 , \IDinst/n5524 ,
         \IDinst/n5523 , \IDinst/n5522 , \IDinst/n5521 , \IDinst/n5520 ,
         \IDinst/n5519 , \IDinst/n5518 , \IDinst/n5517 , \IDinst/n5516 ,
         \IDinst/n5515 , \IDinst/n5514 , \IDinst/n5513 , \IDinst/n5512 ,
         \IDinst/n5511 , \IDinst/n5510 , \IDinst/n5509 , \IDinst/n5508 ,
         \IDinst/n5507 , \IDinst/n5506 , \IDinst/n5505 , \IDinst/n5504 ,
         \IDinst/n5503 , \IDinst/n5502 , \IDinst/n5501 , \IDinst/n5500 ,
         \IDinst/n5499 , \IDinst/n5498 , \IDinst/n5497 , \IDinst/n5496 ,
         \IDinst/n5495 , \IDinst/n5494 , \IDinst/n5493 , \IDinst/n5492 ,
         \IDinst/n5491 , \IDinst/n5490 , \IDinst/n5489 , \IDinst/n5488 ,
         \IDinst/n5487 , \IDinst/n5486 , \IDinst/n5485 , \IDinst/n5484 ,
         \IDinst/n5483 , \IDinst/n5482 , \IDinst/n5481 , \IDinst/n5480 ,
         \IDinst/n5479 , \IDinst/n5478 , \IDinst/n5477 , \IDinst/n5476 ,
         \IDinst/n5475 , \IDinst/n5474 , \IDinst/n5473 , \IDinst/n5472 ,
         \IDinst/n5471 , \IDinst/n5470 , \IDinst/n5469 , \IDinst/n5468 ,
         \IDinst/n5467 , \IDinst/n5466 , \IDinst/n5465 , \IDinst/n5464 ,
         \IDinst/n5463 , \IDinst/n5462 , \IDinst/n5461 , \IDinst/n5460 ,
         \IDinst/n5459 , \IDinst/n5458 , \IDinst/n5457 , \IDinst/n5456 ,
         \IDinst/n5455 , \IDinst/n5454 , \IDinst/n5453 , \IDinst/n5452 ,
         \IDinst/n5451 , \IDinst/n5450 , \IDinst/n5449 , \IDinst/n5448 ,
         \IDinst/n5447 , \IDinst/n5446 , \IDinst/n5445 , \IDinst/n5444 ,
         \IDinst/n5443 , \IDinst/n5442 , \IDinst/n5441 , \IDinst/n5440 ,
         \IDinst/n5439 , \IDinst/n5438 , \IDinst/n5437 , \IDinst/n5436 ,
         \IDinst/n5435 , \IDinst/n5434 , \IDinst/n5433 , \IDinst/n5432 ,
         \IDinst/n5431 , \IDinst/n5430 , \IDinst/n5429 , \IDinst/n5428 ,
         \IDinst/n5427 , \IDinst/n5426 , \IDinst/n5425 , \IDinst/n5424 ,
         \IDinst/n5423 , \IDinst/n5422 , \IDinst/n5421 , \IDinst/n5420 ,
         \IDinst/n5419 , \IDinst/n5418 , \IDinst/n5417 , \IDinst/n5416 ,
         \IDinst/n5415 , \IDinst/n5414 , \IDinst/n5413 , \IDinst/n5412 ,
         \IDinst/n5411 , \IDinst/n5410 , \IDinst/n5409 , \IDinst/n5408 ,
         \IDinst/n5407 , \IDinst/n5406 , \IDinst/n5405 , \IDinst/n5404 ,
         \IDinst/n5403 , \IDinst/n5402 , \IDinst/n5401 , \IDinst/n5400 ,
         \IDinst/n5399 , \IDinst/n5398 , \IDinst/n5397 , \IDinst/n5396 ,
         \IDinst/n5395 , \IDinst/n5394 , \IDinst/n5393 , \IDinst/n5392 ,
         \IDinst/n5391 , \IDinst/n5390 , \IDinst/n5389 , \IDinst/n5388 ,
         \IDinst/n5387 , \IDinst/n5386 , \IDinst/n5385 , \IDinst/n5384 ,
         \IDinst/n5383 , \IDinst/n5382 , \IDinst/n5381 , \IDinst/n5380 ,
         \IDinst/n5379 , \IDinst/n5378 , \IDinst/n5377 , \IDinst/n5376 ,
         \IDinst/n5375 , \IDinst/n5374 , \IDinst/n5373 , \IDinst/n5372 ,
         \IDinst/n5371 , \IDinst/n5370 , \IDinst/n5369 , \IDinst/n5368 ,
         \IDinst/n5367 , \IDinst/n5366 , \IDinst/n5365 , \IDinst/n5364 ,
         \IDinst/n5363 , \IDinst/n5362 , \IDinst/n5361 , \IDinst/n5360 ,
         \IDinst/n5359 , \IDinst/n5358 , \IDinst/n5357 , \IDinst/n5356 ,
         \IDinst/n5355 , \IDinst/n5354 , \IDinst/n5353 , \IDinst/n5352 ,
         \IDinst/n5351 , \IDinst/n5350 , \IDinst/n5349 , \IDinst/n5348 ,
         \IDinst/n5347 , \IDinst/n5346 , \IDinst/n5345 , \IDinst/n5344 ,
         \IDinst/n5343 , \IDinst/n5342 , \IDinst/n5341 , \IDinst/n5340 ,
         \IDinst/n5339 , \IDinst/n5338 , \IDinst/n5337 , \IDinst/n5336 ,
         \IDinst/n5335 , \IDinst/n5334 , \IDinst/n5333 , \IDinst/n5332 ,
         \IDinst/n5331 , \IDinst/n5330 , \IDinst/n5329 , \IDinst/n5328 ,
         \IDinst/n5327 , \IDinst/n5326 , \IDinst/n5325 , \IDinst/n5324 ,
         \IDinst/n5323 , \IDinst/n5322 , \IDinst/n5321 , \IDinst/n5320 ,
         \IDinst/n5319 , \IDinst/n5318 , \IDinst/n5317 , \IDinst/n5316 ,
         \IDinst/n5315 , \IDinst/n5314 , \IDinst/n5313 , \IDinst/n5312 ,
         \IDinst/n5311 , \IDinst/n5310 , \IDinst/n5309 , \IDinst/n5308 ,
         \IDinst/n5307 , \IDinst/n5306 , \IDinst/n5305 , \IDinst/n5304 ,
         \IDinst/n5303 , \IDinst/n5302 , \IDinst/n5301 , \IDinst/n5300 ,
         \IDinst/n5299 , \IDinst/n5298 , \IDinst/n5297 , \IDinst/n5296 ,
         \IDinst/n5295 , \IDinst/n5294 , \IDinst/n5293 , \IDinst/n5292 ,
         \IDinst/n5291 , \IDinst/n5290 , \IDinst/n5289 , \IDinst/n5288 ,
         \IDinst/n5287 , \IDinst/n5286 , \IDinst/n5285 , \IDinst/n5284 ,
         \IDinst/n5283 , \IDinst/n5282 , \IDinst/n5281 , \IDinst/n5280 ,
         \IDinst/n5279 , \IDinst/n5278 , \IDinst/n5277 , \IDinst/n5276 ,
         \IDinst/n5275 , \IDinst/n5274 , \IDinst/n5273 , \IDinst/n5272 ,
         \IDinst/n5271 , \IDinst/n5270 , \IDinst/n5269 , \IDinst/n5268 ,
         \IDinst/n5267 , \IDinst/n5266 , \IDinst/n5265 , \IDinst/n5264 ,
         \IDinst/n5263 , \IDinst/n5262 , \IDinst/n5261 , \IDinst/n5260 ,
         \IDinst/n5259 , \IDinst/n5258 , \IDinst/n5257 , \IDinst/n5256 ,
         \IDinst/n5255 , \IDinst/n5254 , \IDinst/n5253 , \IDinst/n5252 ,
         \IDinst/n5251 , \IDinst/n5250 , \IDinst/n5249 , \IDinst/n5248 ,
         \IDinst/n5247 , \IDinst/n5246 , \IDinst/n5245 , \IDinst/n5244 ,
         \IDinst/n5243 , \IDinst/n5242 , \IDinst/n5241 , \IDinst/n5240 ,
         \IDinst/n5239 , \IDinst/n5238 , \IDinst/n5237 , \IDinst/n5236 ,
         \IDinst/n5235 , \IDinst/n5234 , \IDinst/n5233 , \IDinst/n5232 ,
         \IDinst/n5231 , \IDinst/n5230 , \IDinst/n5229 , \IDinst/n5228 ,
         \IDinst/n5227 , \IDinst/n5226 , \IDinst/n5225 , \IDinst/n5224 ,
         \IDinst/n5223 , \IDinst/n5222 , \IDinst/n5221 , \IDinst/n5220 ,
         \IDinst/n5219 , \IDinst/n5218 , \IDinst/n5217 , \IDinst/n5216 ,
         \IDinst/n5215 , \IDinst/n5214 , \IDinst/n5213 , \IDinst/n5212 ,
         \IDinst/n5211 , \IDinst/n5210 , \IDinst/n5209 , \IDinst/n5208 ,
         \IDinst/n5207 , \IDinst/n5206 , \IDinst/n5205 , \IDinst/n5204 ,
         \IDinst/n5203 , \IDinst/n5202 , \IDinst/n5201 , \IDinst/n5200 ,
         \IDinst/n5199 , \IDinst/n5198 , \IDinst/n5197 , \IDinst/n5196 ,
         \IDinst/n5195 , \IDinst/n5194 , \IDinst/n5193 , \IDinst/n5192 ,
         \IDinst/n5191 , \IDinst/n5190 , \IDinst/n5189 , \IDinst/n5188 ,
         \IDinst/n5187 , \IDinst/n5186 , \IDinst/n5185 , \IDinst/n5184 ,
         \IDinst/n5183 , \IDinst/n5182 , \IDinst/n5181 , \IDinst/n5180 ,
         \IDinst/n5179 , \IDinst/n5178 , \IDinst/n5177 , \IDinst/n5176 ,
         \IDinst/n5175 , \IDinst/n5174 , \IDinst/n5173 , \IDinst/n5172 ,
         \IDinst/n5171 , \IDinst/n5170 , \IDinst/n5169 , \IDinst/n5168 ,
         \IDinst/n5167 , \IDinst/n5166 , \IDinst/n5165 , \IDinst/n5164 ,
         \IDinst/n5163 , \IDinst/n5162 , \IDinst/n5161 , \IDinst/n5160 ,
         \IDinst/n5159 , \IDinst/n5158 , \IDinst/n5157 , \IDinst/n5156 ,
         \IDinst/n5155 , \IDinst/n5154 , \IDinst/n5153 , \IDinst/n5152 ,
         \IDinst/n5151 , \IDinst/n5150 , \IDinst/n5149 , \IDinst/n5148 ,
         \IDinst/n5147 , \IDinst/n5146 , \IDinst/n5145 , \IDinst/n5144 ,
         \IDinst/n5143 , \IDinst/n5142 , \IDinst/n5141 , \IDinst/n5140 ,
         \IDinst/n5139 , \IDinst/n5138 , \IDinst/n5137 , \IDinst/n5136 ,
         \IDinst/n5135 , \IDinst/n5134 , \IDinst/n5133 , \IDinst/n5132 ,
         \IDinst/n5131 , \IDinst/n5130 , \IDinst/n5129 , \IDinst/n5128 ,
         \IDinst/n5127 , \IDinst/n5126 , \IDinst/n5125 , \IDinst/n5124 ,
         \IDinst/n5123 , \IDinst/n5122 , \IDinst/n5121 , \IDinst/n5120 ,
         \IDinst/n5119 , \IDinst/n5118 , \IDinst/n5117 , \IDinst/n5116 ,
         \IDinst/n5115 , \IDinst/n5114 , \IDinst/n5113 , \IDinst/n5112 ,
         \IDinst/n5111 , \IDinst/n5110 , \IDinst/n5109 , \IDinst/n5108 ,
         \IDinst/n5107 , \IDinst/n5106 , \IDinst/n5105 , \IDinst/n5104 ,
         \IDinst/n5103 , \IDinst/n5102 , \IDinst/n5101 , \IDinst/n5100 ,
         \IDinst/n5099 , \IDinst/n5098 , \IDinst/n5097 , \IDinst/n5096 ,
         \IDinst/n5095 , \IDinst/n5094 , \IDinst/n5093 , \IDinst/n5092 ,
         \IDinst/n5091 , \IDinst/n5090 , \IDinst/n5089 , \IDinst/n5088 ,
         \IDinst/n5087 , \IDinst/n5086 , \IDinst/n5085 , \IDinst/n5084 ,
         \IDinst/n5083 , \IDinst/n5082 , \IDinst/n5081 , \IDinst/n5080 ,
         \IDinst/n5079 , \IDinst/n5078 , \IDinst/n5077 , \IDinst/n5076 ,
         \IDinst/n5075 , \IDinst/n5074 , \IDinst/n5073 , \IDinst/n5072 ,
         \IDinst/n5071 , \IDinst/n5070 , \IDinst/n5069 , \IDinst/n5068 ,
         \IDinst/n5067 , \IDinst/n5066 , \IDinst/n5065 , \IDinst/n5064 ,
         \IDinst/n5063 , \IDinst/n5062 , \IDinst/n5061 , \IDinst/n5060 ,
         \IDinst/n5059 , \IDinst/n5058 , \IDinst/n5057 , \IDinst/n5056 ,
         \IDinst/n5055 , \IDinst/n5054 , \IDinst/n5053 , \IDinst/n5052 ,
         \IDinst/n5051 , \IDinst/n5050 , \IDinst/n5049 , \IDinst/n5048 ,
         \IDinst/n5047 , \IDinst/n5046 , \IDinst/n5045 , \IDinst/n5044 ,
         \IDinst/n5043 , \IDinst/n5042 , \IDinst/n5041 , \IDinst/n5040 ,
         \IDinst/n5039 , \IDinst/n5038 , \IDinst/n5037 , \IDinst/n5036 ,
         \IDinst/n5035 , \IDinst/n5034 , \IDinst/n5033 , \IDinst/n5032 ,
         \IDinst/n5031 , \IDinst/n5030 , \IDinst/n5029 , \IDinst/n5028 ,
         \IDinst/n5027 , \IDinst/n5026 , \IDinst/n5025 , \IDinst/n5024 ,
         \IDinst/n5023 , \IDinst/n5022 , \IDinst/n5021 , \IDinst/n5020 ,
         \IDinst/n5019 , \IDinst/n5018 , \IDinst/n5017 , \IDinst/n5016 ,
         \IDinst/n5015 , \IDinst/n5014 , \IDinst/n5013 , \IDinst/n5012 ,
         \IDinst/n5011 , \IDinst/n5010 , \IDinst/n5009 , \IDinst/n5008 ,
         \IDinst/n5007 , \IDinst/n5006 , \IDinst/n5005 , \IDinst/n5004 ,
         \IDinst/n5003 , \IDinst/n5002 , \IDinst/n5001 , \IDinst/n5000 ,
         \IDinst/n4999 , \IDinst/n4998 , \IDinst/n4997 , \IDinst/n4996 ,
         \IDinst/n4995 , \IDinst/n4994 , \IDinst/n4993 , \IDinst/n4992 ,
         \IDinst/n4991 , \IDinst/n4990 , \IDinst/n4989 , \IDinst/n4988 ,
         \IDinst/n4987 , \IDinst/n4986 , \IDinst/n4985 , \IDinst/n4984 ,
         \IDinst/n4983 , \IDinst/n4982 , \IDinst/n4981 , \IDinst/n4980 ,
         \IDinst/n4979 , \IDinst/n4978 , \IDinst/n4977 , \IDinst/n4976 ,
         \IDinst/n4975 , \IDinst/n4974 , \IDinst/n4973 , \IDinst/n4972 ,
         \IDinst/n4971 , \IDinst/n4970 , \IDinst/n4969 , \IDinst/n4968 ,
         \IDinst/n4967 , \IDinst/n4966 , \IDinst/n4965 , \IDinst/n4964 ,
         \IDinst/n4963 , \IDinst/n4962 , \IDinst/n4961 , \IDinst/n4960 ,
         \IDinst/n4959 , \IDinst/n4958 , \IDinst/n4957 , \IDinst/n4956 ,
         \IDinst/n4955 , \IDinst/n4954 , \IDinst/n4953 , \IDinst/n4952 ,
         \IDinst/n4951 , \IDinst/n4950 , \IDinst/n4949 , \IDinst/n4948 ,
         \IDinst/n4947 , \IDinst/n4946 , \IDinst/n4945 , \IDinst/n4944 ,
         \IDinst/n4943 , \IDinst/n4942 , \IDinst/n4941 , \IDinst/n4940 ,
         \IDinst/n4939 , \IDinst/n4938 , \IDinst/n4937 , \IDinst/n4936 ,
         \IDinst/n4935 , \IDinst/n4934 , \IDinst/n4933 , \IDinst/n4932 ,
         \IDinst/n4931 , \IDinst/n4930 , \IDinst/n4929 , \IDinst/n4928 ,
         \IDinst/n4927 , \IDinst/n4926 , \IDinst/n4925 , \IDinst/n4924 ,
         \IDinst/n4923 , \IDinst/n4922 , \IDinst/n4921 , \IDinst/n4920 ,
         \IDinst/n4919 , \IDinst/n4918 , \IDinst/n4917 , \IDinst/n4916 ,
         \IDinst/n4915 , \IDinst/n4914 , \IDinst/n4913 , \IDinst/n4912 ,
         \IDinst/n4911 , \IDinst/n4910 , \IDinst/n4909 , \IDinst/n4908 ,
         \IDinst/n4907 , \IDinst/n4906 , \IDinst/n4905 , \IDinst/n4904 ,
         \IDinst/n4903 , \IDinst/n4902 , \IDinst/n4901 , \IDinst/n4900 ,
         \IDinst/n4899 , \IDinst/n4898 , \IDinst/n4897 , \IDinst/n4896 ,
         \IDinst/n4895 , \IDinst/n4894 , \IDinst/n4893 , \IDinst/n4892 ,
         \IDinst/n4891 , \IDinst/n4890 , \IDinst/n4889 , \IDinst/n4888 ,
         \IDinst/n4887 , \IDinst/n4886 , \IDinst/n4885 , \IDinst/n4884 ,
         \IDinst/n4883 , \IDinst/n4882 , \IDinst/n4881 , \IDinst/n4880 ,
         \IDinst/n4879 , \IDinst/n4878 , \IDinst/n4877 , \IDinst/n4876 ,
         \IDinst/n4875 , \IDinst/n4874 , \IDinst/n4873 , \IDinst/n4872 ,
         \IDinst/n4871 , \IDinst/n4870 , \IDinst/n4869 , \IDinst/n4868 ,
         \IDinst/n4867 , \IDinst/n4866 , \IDinst/n4865 , \IDinst/n4864 ,
         \IDinst/n4863 , \IDinst/n4862 , \IDinst/n4861 , \IDinst/n4860 ,
         \IDinst/n4859 , \IDinst/n4858 , \IDinst/n4857 , \IDinst/n4856 ,
         \IDinst/n4855 , \IDinst/n4854 , \IDinst/n4853 , \IDinst/n4852 ,
         \IDinst/n4851 , \IDinst/n4850 , \IDinst/n4849 , \IDinst/n4848 ,
         \IDinst/n4847 , \IDinst/n4846 , \IDinst/n4845 , \IDinst/n4844 ,
         \IDinst/n4843 , \IDinst/n4842 , \IDinst/n4841 , \IDinst/n4840 ,
         \IDinst/n4839 , \IDinst/n4838 , \IDinst/n4837 , \IDinst/n4836 ,
         \IDinst/n4835 , \IDinst/n4834 , \IDinst/n4833 , \IDinst/n4832 ,
         \IDinst/n4831 , \IDinst/n4830 , \IDinst/n4829 , \IDinst/n4828 ,
         \IDinst/n4827 , \IDinst/n4826 , \IDinst/n4825 , \IDinst/n4824 ,
         \IDinst/n4823 , \IDinst/n4822 , \IDinst/n4821 , \IDinst/n4820 ,
         \IDinst/n4819 , \IDinst/n4818 , \IDinst/n4817 , \IDinst/n4816 ,
         \IDinst/n4815 , \IDinst/n4814 , \IDinst/n4813 , \IDinst/n4812 ,
         \IDinst/n4811 , \IDinst/n4810 , \IDinst/n4809 , \IDinst/n4808 ,
         \IDinst/n4807 , \IDinst/n4806 , \IDinst/n4805 , \IDinst/n4804 ,
         \IDinst/n4803 , \IDinst/n4802 , \IDinst/n4801 , \IDinst/n4800 ,
         \IDinst/n4799 , \IDinst/n4798 , \IDinst/n4797 , \IDinst/n4796 ,
         \IDinst/n4795 , \IDinst/n4794 , \IDinst/n4793 , \IDinst/n4792 ,
         \IDinst/n4791 , \IDinst/n4790 , \IDinst/n4789 , \IDinst/n4788 ,
         \IDinst/n4787 , \IDinst/n4786 , \IDinst/n4785 , \IDinst/n4784 ,
         \IDinst/n4783 , \IDinst/n4782 , \IDinst/n4781 , \IDinst/n4780 ,
         \IDinst/n4779 , \IDinst/n4778 , \IDinst/n4777 , \IDinst/n4776 ,
         \IDinst/n4775 , \IDinst/n4774 , \IDinst/n4773 , \IDinst/n4772 ,
         \IDinst/n4771 , \IDinst/n4770 , \IDinst/n4769 , \IDinst/n4768 ,
         \IDinst/n4767 , \IDinst/n4766 , \IDinst/n4765 , \IDinst/n4764 ,
         \IDinst/n4763 , \IDinst/n4762 , \IDinst/n4761 , \IDinst/n4760 ,
         \IDinst/n4759 , \IDinst/n4758 , \IDinst/n4757 , \IDinst/n4756 ,
         \IDinst/n4755 , \IDinst/n4754 , \IDinst/n4753 , \IDinst/n4752 ,
         \IDinst/n4751 , \IDinst/n4750 , \IDinst/n4749 , \IDinst/n4748 ,
         \IDinst/n4747 , \IDinst/n4746 , \IDinst/n4745 , \IDinst/n4744 ,
         \IDinst/n4743 , \IDinst/n4742 , \IDinst/n4741 , \IDinst/n4740 ,
         \IDinst/n4739 , \IDinst/n4738 , \IDinst/n4737 , \IDinst/n4736 ,
         \IDinst/n4735 , \IDinst/n4734 , \IDinst/n4733 , \IDinst/n4732 ,
         \IDinst/n4731 , \IDinst/n4730 , \IDinst/n4729 , \IDinst/n1445 ,
         \IDinst/n1444 , \IDinst/n1440 , \IDinst/n1433 , \IDinst/n1432 ,
         \IDinst/n1431 , \IDinst/n1430 , \IDinst/n1403 , \IDinst/N1055 ,
         \IDinst/N1054 , \IDinst/N1053 , \IDinst/N1052 , \IDinst/N1051 ,
         \IDinst/N1050 , \IDinst/N1049 , \IDinst/N1048 , \IDinst/N1047 ,
         \IDinst/N1046 , \IDinst/N1045 , \IDinst/N1044 , \IDinst/N1043 ,
         \IDinst/N1042 , \IDinst/N1041 , \IDinst/N1040 , \IDinst/N1039 ,
         \IDinst/N1038 , \IDinst/N1037 , \IDinst/N1036 , \IDinst/N1035 ,
         \IDinst/N1034 , \IDinst/N1033 , \IDinst/N1032 , \IDinst/N1031 ,
         \IDinst/N1030 , \IDinst/N1029 , \IDinst/N1028 , \IDinst/N1027 ,
         \IDinst/N1026 , \IDinst/N1025 , \IDinst/N1024 , \IDinst/N1023 ,
         \IDinst/N1022 , \IDinst/N1021 , \IDinst/N1020 , \IDinst/N1019 ,
         \IDinst/N1018 , \IDinst/N1017 , \IDinst/N1016 , \IDinst/N1015 ,
         \IDinst/N1014 , \IDinst/N1013 , \IDinst/N1012 , \IDinst/N1011 ,
         \IDinst/N1010 , \IDinst/N1009 , \IDinst/N1008 , \IDinst/N1007 ,
         \IDinst/N1006 , \IDinst/N1005 , \IDinst/N1004 , \IDinst/N1003 ,
         \IDinst/N1002 , \IDinst/N1001 , \IDinst/N1000 , \IDinst/N999 ,
         \IDinst/N998 , \IDinst/N997 , \IDinst/N996 , \IDinst/N995 ,
         \IDinst/N994 , \IDinst/N993 , \IDinst/N992 , \IDinst/opcode_of_WB[2] ,
         \IDinst/N120 , \IDinst/N119 , \IDinst/N118 , \IDinst/N117 ,
         \IDinst/N116 , \IDinst/N115 , \IDinst/N114 , \IDinst/N113 ,
         \IDinst/N112 , \IDinst/N111 , \IDinst/N110 , \IDinst/N109 ,
         \IDinst/N108 , \IDinst/N107 , \IDinst/N106 , \IDinst/N105 ,
         \IDinst/N104 , \IDinst/N103 , \IDinst/N102 , \IDinst/N101 ,
         \IDinst/N100 , \IDinst/N99 , \IDinst/N98 , \IDinst/N97 , \IDinst/N96 ,
         \IDinst/N95 , \IDinst/N94 , \IDinst/N93 , \IDinst/N92 , \IDinst/N91 ,
         \IDinst/N90 , \IDinst/N89 , \IDinst/N85 , \IDinst/N84 , \IDinst/N83 ,
         \IDinst/N82 , \IDinst/N81 , \IDinst/N80 , \IDinst/N79 , \IDinst/N78 ,
         \IDinst/N77 , \IDinst/N76 , \IDinst/N75 , \IDinst/N74 , \IDinst/N73 ,
         \IDinst/N72 , \IDinst/N71 , \IDinst/N70 , \IDinst/N69 , \IDinst/N68 ,
         \IDinst/N67 , \IDinst/N66 , \IDinst/N65 , \IDinst/N64 , \IDinst/N63 ,
         \IDinst/N62 , \IDinst/N61 , \IDinst/N60 , \IDinst/N59 , \IDinst/N58 ,
         \IDinst/N57 , \IDinst/N56 , \IDinst/N55 , \IDinst/N54 ,
         \IDinst/RegFile[0][31] , \IDinst/RegFile[0][30] ,
         \IDinst/RegFile[0][29] , \IDinst/RegFile[0][28] ,
         \IDinst/RegFile[0][27] , \IDinst/RegFile[0][26] ,
         \IDinst/RegFile[0][25] , \IDinst/RegFile[0][24] ,
         \IDinst/RegFile[0][23] , \IDinst/RegFile[0][22] ,
         \IDinst/RegFile[0][21] , \IDinst/RegFile[0][20] ,
         \IDinst/RegFile[0][19] , \IDinst/RegFile[0][18] ,
         \IDinst/RegFile[0][17] , \IDinst/RegFile[0][16] ,
         \IDinst/RegFile[0][15] , \IDinst/RegFile[0][14] ,
         \IDinst/RegFile[0][13] , \IDinst/RegFile[0][12] ,
         \IDinst/RegFile[0][11] , \IDinst/RegFile[0][10] ,
         \IDinst/RegFile[0][9] , \IDinst/RegFile[0][8] ,
         \IDinst/RegFile[0][7] , \IDinst/RegFile[0][6] ,
         \IDinst/RegFile[0][5] , \IDinst/RegFile[0][4] ,
         \IDinst/RegFile[0][3] , \IDinst/RegFile[0][2] ,
         \IDinst/RegFile[0][1] , \IDinst/RegFile[0][0] ,
         \IDinst/RegFile[1][31] , \IDinst/RegFile[1][30] ,
         \IDinst/RegFile[1][29] , \IDinst/RegFile[1][28] ,
         \IDinst/RegFile[1][27] , \IDinst/RegFile[1][26] ,
         \IDinst/RegFile[1][25] , \IDinst/RegFile[1][24] ,
         \IDinst/RegFile[1][23] , \IDinst/RegFile[1][22] ,
         \IDinst/RegFile[1][21] , \IDinst/RegFile[1][20] ,
         \IDinst/RegFile[1][19] , \IDinst/RegFile[1][18] ,
         \IDinst/RegFile[1][17] , \IDinst/RegFile[1][16] ,
         \IDinst/RegFile[1][15] , \IDinst/RegFile[1][14] ,
         \IDinst/RegFile[1][13] , \IDinst/RegFile[1][12] ,
         \IDinst/RegFile[1][11] , \IDinst/RegFile[1][10] ,
         \IDinst/RegFile[1][9] , \IDinst/RegFile[1][8] ,
         \IDinst/RegFile[1][7] , \IDinst/RegFile[1][6] ,
         \IDinst/RegFile[1][5] , \IDinst/RegFile[1][4] ,
         \IDinst/RegFile[1][3] , \IDinst/RegFile[1][2] ,
         \IDinst/RegFile[1][1] , \IDinst/RegFile[1][0] ,
         \IDinst/RegFile[2][31] , \IDinst/RegFile[2][30] ,
         \IDinst/RegFile[2][29] , \IDinst/RegFile[2][28] ,
         \IDinst/RegFile[2][27] , \IDinst/RegFile[2][26] ,
         \IDinst/RegFile[2][25] , \IDinst/RegFile[2][24] ,
         \IDinst/RegFile[2][23] , \IDinst/RegFile[2][22] ,
         \IDinst/RegFile[2][21] , \IDinst/RegFile[2][20] ,
         \IDinst/RegFile[2][19] , \IDinst/RegFile[2][18] ,
         \IDinst/RegFile[2][17] , \IDinst/RegFile[2][16] ,
         \IDinst/RegFile[2][15] , \IDinst/RegFile[2][14] ,
         \IDinst/RegFile[2][13] , \IDinst/RegFile[2][12] ,
         \IDinst/RegFile[2][11] , \IDinst/RegFile[2][10] ,
         \IDinst/RegFile[2][9] , \IDinst/RegFile[2][8] ,
         \IDinst/RegFile[2][7] , \IDinst/RegFile[2][6] ,
         \IDinst/RegFile[2][5] , \IDinst/RegFile[2][4] ,
         \IDinst/RegFile[2][3] , \IDinst/RegFile[2][2] ,
         \IDinst/RegFile[2][1] , \IDinst/RegFile[2][0] ,
         \IDinst/RegFile[3][31] , \IDinst/RegFile[3][30] ,
         \IDinst/RegFile[3][29] , \IDinst/RegFile[3][28] ,
         \IDinst/RegFile[3][27] , \IDinst/RegFile[3][26] ,
         \IDinst/RegFile[3][25] , \IDinst/RegFile[3][24] ,
         \IDinst/RegFile[3][23] , \IDinst/RegFile[3][22] ,
         \IDinst/RegFile[3][21] , \IDinst/RegFile[3][20] ,
         \IDinst/RegFile[3][19] , \IDinst/RegFile[3][18] ,
         \IDinst/RegFile[3][17] , \IDinst/RegFile[3][16] ,
         \IDinst/RegFile[3][15] , \IDinst/RegFile[3][14] ,
         \IDinst/RegFile[3][13] , \IDinst/RegFile[3][12] ,
         \IDinst/RegFile[3][11] , \IDinst/RegFile[3][10] ,
         \IDinst/RegFile[3][9] , \IDinst/RegFile[3][8] ,
         \IDinst/RegFile[3][7] , \IDinst/RegFile[3][6] ,
         \IDinst/RegFile[3][5] , \IDinst/RegFile[3][4] ,
         \IDinst/RegFile[3][3] , \IDinst/RegFile[3][2] ,
         \IDinst/RegFile[3][1] , \IDinst/RegFile[3][0] ,
         \IDinst/RegFile[4][31] , \IDinst/RegFile[4][30] ,
         \IDinst/RegFile[4][29] , \IDinst/RegFile[4][28] ,
         \IDinst/RegFile[4][27] , \IDinst/RegFile[4][26] ,
         \IDinst/RegFile[4][25] , \IDinst/RegFile[4][24] ,
         \IDinst/RegFile[4][23] , \IDinst/RegFile[4][22] ,
         \IDinst/RegFile[4][21] , \IDinst/RegFile[4][20] ,
         \IDinst/RegFile[4][19] , \IDinst/RegFile[4][18] ,
         \IDinst/RegFile[4][17] , \IDinst/RegFile[4][16] ,
         \IDinst/RegFile[4][15] , \IDinst/RegFile[4][14] ,
         \IDinst/RegFile[4][13] , \IDinst/RegFile[4][12] ,
         \IDinst/RegFile[4][11] , \IDinst/RegFile[4][10] ,
         \IDinst/RegFile[4][9] , \IDinst/RegFile[4][8] ,
         \IDinst/RegFile[4][7] , \IDinst/RegFile[4][6] ,
         \IDinst/RegFile[4][5] , \IDinst/RegFile[4][4] ,
         \IDinst/RegFile[4][3] , \IDinst/RegFile[4][2] ,
         \IDinst/RegFile[4][1] , \IDinst/RegFile[4][0] ,
         \IDinst/RegFile[5][31] , \IDinst/RegFile[5][30] ,
         \IDinst/RegFile[5][29] , \IDinst/RegFile[5][28] ,
         \IDinst/RegFile[5][27] , \IDinst/RegFile[5][26] ,
         \IDinst/RegFile[5][25] , \IDinst/RegFile[5][24] ,
         \IDinst/RegFile[5][23] , \IDinst/RegFile[5][22] ,
         \IDinst/RegFile[5][21] , \IDinst/RegFile[5][20] ,
         \IDinst/RegFile[5][19] , \IDinst/RegFile[5][18] ,
         \IDinst/RegFile[5][17] , \IDinst/RegFile[5][16] ,
         \IDinst/RegFile[5][15] , \IDinst/RegFile[5][14] ,
         \IDinst/RegFile[5][13] , \IDinst/RegFile[5][12] ,
         \IDinst/RegFile[5][11] , \IDinst/RegFile[5][10] ,
         \IDinst/RegFile[5][9] , \IDinst/RegFile[5][8] ,
         \IDinst/RegFile[5][7] , \IDinst/RegFile[5][6] ,
         \IDinst/RegFile[5][5] , \IDinst/RegFile[5][4] ,
         \IDinst/RegFile[5][3] , \IDinst/RegFile[5][2] ,
         \IDinst/RegFile[5][1] , \IDinst/RegFile[5][0] ,
         \IDinst/RegFile[6][31] , \IDinst/RegFile[6][30] ,
         \IDinst/RegFile[6][29] , \IDinst/RegFile[6][28] ,
         \IDinst/RegFile[6][27] , \IDinst/RegFile[6][26] ,
         \IDinst/RegFile[6][25] , \IDinst/RegFile[6][24] ,
         \IDinst/RegFile[6][23] , \IDinst/RegFile[6][22] ,
         \IDinst/RegFile[6][21] , \IDinst/RegFile[6][20] ,
         \IDinst/RegFile[6][19] , \IDinst/RegFile[6][18] ,
         \IDinst/RegFile[6][17] , \IDinst/RegFile[6][16] ,
         \IDinst/RegFile[6][15] , \IDinst/RegFile[6][14] ,
         \IDinst/RegFile[6][13] , \IDinst/RegFile[6][12] ,
         \IDinst/RegFile[6][11] , \IDinst/RegFile[6][10] ,
         \IDinst/RegFile[6][9] , \IDinst/RegFile[6][8] ,
         \IDinst/RegFile[6][7] , \IDinst/RegFile[6][6] ,
         \IDinst/RegFile[6][5] , \IDinst/RegFile[6][4] ,
         \IDinst/RegFile[6][3] , \IDinst/RegFile[6][2] ,
         \IDinst/RegFile[6][1] , \IDinst/RegFile[6][0] ,
         \IDinst/RegFile[7][31] , \IDinst/RegFile[7][30] ,
         \IDinst/RegFile[7][29] , \IDinst/RegFile[7][28] ,
         \IDinst/RegFile[7][27] , \IDinst/RegFile[7][26] ,
         \IDinst/RegFile[7][25] , \IDinst/RegFile[7][24] ,
         \IDinst/RegFile[7][23] , \IDinst/RegFile[7][22] ,
         \IDinst/RegFile[7][21] , \IDinst/RegFile[7][20] ,
         \IDinst/RegFile[7][19] , \IDinst/RegFile[7][18] ,
         \IDinst/RegFile[7][17] , \IDinst/RegFile[7][16] ,
         \IDinst/RegFile[7][15] , \IDinst/RegFile[7][14] ,
         \IDinst/RegFile[7][13] , \IDinst/RegFile[7][12] ,
         \IDinst/RegFile[7][11] , \IDinst/RegFile[7][10] ,
         \IDinst/RegFile[7][9] , \IDinst/RegFile[7][8] ,
         \IDinst/RegFile[7][7] , \IDinst/RegFile[7][6] ,
         \IDinst/RegFile[7][5] , \IDinst/RegFile[7][4] ,
         \IDinst/RegFile[7][3] , \IDinst/RegFile[7][2] ,
         \IDinst/RegFile[7][1] , \IDinst/RegFile[7][0] ,
         \IDinst/RegFile[8][31] , \IDinst/RegFile[8][30] ,
         \IDinst/RegFile[8][29] , \IDinst/RegFile[8][28] ,
         \IDinst/RegFile[8][27] , \IDinst/RegFile[8][26] ,
         \IDinst/RegFile[8][25] , \IDinst/RegFile[8][24] ,
         \IDinst/RegFile[8][23] , \IDinst/RegFile[8][22] ,
         \IDinst/RegFile[8][21] , \IDinst/RegFile[8][20] ,
         \IDinst/RegFile[8][19] , \IDinst/RegFile[8][18] ,
         \IDinst/RegFile[8][17] , \IDinst/RegFile[8][16] ,
         \IDinst/RegFile[8][15] , \IDinst/RegFile[8][14] ,
         \IDinst/RegFile[8][13] , \IDinst/RegFile[8][12] ,
         \IDinst/RegFile[8][11] , \IDinst/RegFile[8][10] ,
         \IDinst/RegFile[8][9] , \IDinst/RegFile[8][8] ,
         \IDinst/RegFile[8][7] , \IDinst/RegFile[8][6] ,
         \IDinst/RegFile[8][5] , \IDinst/RegFile[8][4] ,
         \IDinst/RegFile[8][3] , \IDinst/RegFile[8][2] ,
         \IDinst/RegFile[8][1] , \IDinst/RegFile[8][0] ,
         \IDinst/RegFile[9][31] , \IDinst/RegFile[9][30] ,
         \IDinst/RegFile[9][29] , \IDinst/RegFile[9][28] ,
         \IDinst/RegFile[9][27] , \IDinst/RegFile[9][26] ,
         \IDinst/RegFile[9][25] , \IDinst/RegFile[9][24] ,
         \IDinst/RegFile[9][23] , \IDinst/RegFile[9][22] ,
         \IDinst/RegFile[9][21] , \IDinst/RegFile[9][20] ,
         \IDinst/RegFile[9][19] , \IDinst/RegFile[9][18] ,
         \IDinst/RegFile[9][17] , \IDinst/RegFile[9][16] ,
         \IDinst/RegFile[9][15] , \IDinst/RegFile[9][14] ,
         \IDinst/RegFile[9][13] , \IDinst/RegFile[9][12] ,
         \IDinst/RegFile[9][11] , \IDinst/RegFile[9][10] ,
         \IDinst/RegFile[9][9] , \IDinst/RegFile[9][8] ,
         \IDinst/RegFile[9][7] , \IDinst/RegFile[9][6] ,
         \IDinst/RegFile[9][5] , \IDinst/RegFile[9][4] ,
         \IDinst/RegFile[9][3] , \IDinst/RegFile[9][2] ,
         \IDinst/RegFile[9][1] , \IDinst/RegFile[9][0] ,
         \IDinst/RegFile[10][31] , \IDinst/RegFile[10][30] ,
         \IDinst/RegFile[10][29] , \IDinst/RegFile[10][28] ,
         \IDinst/RegFile[10][27] , \IDinst/RegFile[10][26] ,
         \IDinst/RegFile[10][25] , \IDinst/RegFile[10][24] ,
         \IDinst/RegFile[10][23] , \IDinst/RegFile[10][22] ,
         \IDinst/RegFile[10][21] , \IDinst/RegFile[10][20] ,
         \IDinst/RegFile[10][19] , \IDinst/RegFile[10][18] ,
         \IDinst/RegFile[10][17] , \IDinst/RegFile[10][16] ,
         \IDinst/RegFile[10][15] , \IDinst/RegFile[10][14] ,
         \IDinst/RegFile[10][13] , \IDinst/RegFile[10][12] ,
         \IDinst/RegFile[10][11] , \IDinst/RegFile[10][10] ,
         \IDinst/RegFile[10][9] , \IDinst/RegFile[10][8] ,
         \IDinst/RegFile[10][7] , \IDinst/RegFile[10][6] ,
         \IDinst/RegFile[10][5] , \IDinst/RegFile[10][4] ,
         \IDinst/RegFile[10][3] , \IDinst/RegFile[10][2] ,
         \IDinst/RegFile[10][1] , \IDinst/RegFile[10][0] ,
         \IDinst/RegFile[11][31] , \IDinst/RegFile[11][30] ,
         \IDinst/RegFile[11][29] , \IDinst/RegFile[11][28] ,
         \IDinst/RegFile[11][27] , \IDinst/RegFile[11][26] ,
         \IDinst/RegFile[11][25] , \IDinst/RegFile[11][24] ,
         \IDinst/RegFile[11][23] , \IDinst/RegFile[11][22] ,
         \IDinst/RegFile[11][21] , \IDinst/RegFile[11][20] ,
         \IDinst/RegFile[11][19] , \IDinst/RegFile[11][18] ,
         \IDinst/RegFile[11][17] , \IDinst/RegFile[11][16] ,
         \IDinst/RegFile[11][15] , \IDinst/RegFile[11][14] ,
         \IDinst/RegFile[11][13] , \IDinst/RegFile[11][12] ,
         \IDinst/RegFile[11][11] , \IDinst/RegFile[11][10] ,
         \IDinst/RegFile[11][9] , \IDinst/RegFile[11][8] ,
         \IDinst/RegFile[11][7] , \IDinst/RegFile[11][6] ,
         \IDinst/RegFile[11][5] , \IDinst/RegFile[11][4] ,
         \IDinst/RegFile[11][3] , \IDinst/RegFile[11][2] ,
         \IDinst/RegFile[11][1] , \IDinst/RegFile[11][0] ,
         \IDinst/RegFile[12][31] , \IDinst/RegFile[12][30] ,
         \IDinst/RegFile[12][29] , \IDinst/RegFile[12][28] ,
         \IDinst/RegFile[12][27] , \IDinst/RegFile[12][26] ,
         \IDinst/RegFile[12][25] , \IDinst/RegFile[12][24] ,
         \IDinst/RegFile[12][23] , \IDinst/RegFile[12][22] ,
         \IDinst/RegFile[12][21] , \IDinst/RegFile[12][20] ,
         \IDinst/RegFile[12][19] , \IDinst/RegFile[12][18] ,
         \IDinst/RegFile[12][17] , \IDinst/RegFile[12][16] ,
         \IDinst/RegFile[12][15] , \IDinst/RegFile[12][14] ,
         \IDinst/RegFile[12][13] , \IDinst/RegFile[12][12] ,
         \IDinst/RegFile[12][11] , \IDinst/RegFile[12][10] ,
         \IDinst/RegFile[12][9] , \IDinst/RegFile[12][8] ,
         \IDinst/RegFile[12][7] , \IDinst/RegFile[12][6] ,
         \IDinst/RegFile[12][5] , \IDinst/RegFile[12][4] ,
         \IDinst/RegFile[12][3] , \IDinst/RegFile[12][2] ,
         \IDinst/RegFile[12][1] , \IDinst/RegFile[12][0] ,
         \IDinst/RegFile[13][31] , \IDinst/RegFile[13][30] ,
         \IDinst/RegFile[13][29] , \IDinst/RegFile[13][28] ,
         \IDinst/RegFile[13][27] , \IDinst/RegFile[13][26] ,
         \IDinst/RegFile[13][25] , \IDinst/RegFile[13][24] ,
         \IDinst/RegFile[13][23] , \IDinst/RegFile[13][22] ,
         \IDinst/RegFile[13][21] , \IDinst/RegFile[13][20] ,
         \IDinst/RegFile[13][19] , \IDinst/RegFile[13][18] ,
         \IDinst/RegFile[13][17] , \IDinst/RegFile[13][16] ,
         \IDinst/RegFile[13][15] , \IDinst/RegFile[13][14] ,
         \IDinst/RegFile[13][13] , \IDinst/RegFile[13][12] ,
         \IDinst/RegFile[13][11] , \IDinst/RegFile[13][10] ,
         \IDinst/RegFile[13][9] , \IDinst/RegFile[13][8] ,
         \IDinst/RegFile[13][7] , \IDinst/RegFile[13][6] ,
         \IDinst/RegFile[13][5] , \IDinst/RegFile[13][4] ,
         \IDinst/RegFile[13][3] , \IDinst/RegFile[13][2] ,
         \IDinst/RegFile[13][1] , \IDinst/RegFile[13][0] ,
         \IDinst/RegFile[14][31] , \IDinst/RegFile[14][30] ,
         \IDinst/RegFile[14][29] , \IDinst/RegFile[14][28] ,
         \IDinst/RegFile[14][27] , \IDinst/RegFile[14][26] ,
         \IDinst/RegFile[14][25] , \IDinst/RegFile[14][24] ,
         \IDinst/RegFile[14][23] , \IDinst/RegFile[14][22] ,
         \IDinst/RegFile[14][21] , \IDinst/RegFile[14][20] ,
         \IDinst/RegFile[14][19] , \IDinst/RegFile[14][18] ,
         \IDinst/RegFile[14][17] , \IDinst/RegFile[14][16] ,
         \IDinst/RegFile[14][15] , \IDinst/RegFile[14][14] ,
         \IDinst/RegFile[14][13] , \IDinst/RegFile[14][12] ,
         \IDinst/RegFile[14][11] , \IDinst/RegFile[14][10] ,
         \IDinst/RegFile[14][9] , \IDinst/RegFile[14][8] ,
         \IDinst/RegFile[14][7] , \IDinst/RegFile[14][6] ,
         \IDinst/RegFile[14][5] , \IDinst/RegFile[14][4] ,
         \IDinst/RegFile[14][3] , \IDinst/RegFile[14][2] ,
         \IDinst/RegFile[14][1] , \IDinst/RegFile[14][0] ,
         \IDinst/RegFile[15][31] , \IDinst/RegFile[15][30] ,
         \IDinst/RegFile[15][29] , \IDinst/RegFile[15][28] ,
         \IDinst/RegFile[15][27] , \IDinst/RegFile[15][26] ,
         \IDinst/RegFile[15][25] , \IDinst/RegFile[15][24] ,
         \IDinst/RegFile[15][23] , \IDinst/RegFile[15][22] ,
         \IDinst/RegFile[15][21] , \IDinst/RegFile[15][20] ,
         \IDinst/RegFile[15][19] , \IDinst/RegFile[15][18] ,
         \IDinst/RegFile[15][17] , \IDinst/RegFile[15][16] ,
         \IDinst/RegFile[15][15] , \IDinst/RegFile[15][14] ,
         \IDinst/RegFile[15][13] , \IDinst/RegFile[15][12] ,
         \IDinst/RegFile[15][11] , \IDinst/RegFile[15][10] ,
         \IDinst/RegFile[15][9] , \IDinst/RegFile[15][8] ,
         \IDinst/RegFile[15][7] , \IDinst/RegFile[15][6] ,
         \IDinst/RegFile[15][5] , \IDinst/RegFile[15][4] ,
         \IDinst/RegFile[15][3] , \IDinst/RegFile[15][2] ,
         \IDinst/RegFile[15][1] , \IDinst/RegFile[15][0] ,
         \IDinst/RegFile[16][31] , \IDinst/RegFile[16][30] ,
         \IDinst/RegFile[16][29] , \IDinst/RegFile[16][28] ,
         \IDinst/RegFile[16][27] , \IDinst/RegFile[16][26] ,
         \IDinst/RegFile[16][25] , \IDinst/RegFile[16][24] ,
         \IDinst/RegFile[16][23] , \IDinst/RegFile[16][22] ,
         \IDinst/RegFile[16][21] , \IDinst/RegFile[16][20] ,
         \IDinst/RegFile[16][19] , \IDinst/RegFile[16][18] ,
         \IDinst/RegFile[16][17] , \IDinst/RegFile[16][16] ,
         \IDinst/RegFile[16][15] , \IDinst/RegFile[16][14] ,
         \IDinst/RegFile[16][13] , \IDinst/RegFile[16][12] ,
         \IDinst/RegFile[16][11] , \IDinst/RegFile[16][10] ,
         \IDinst/RegFile[16][9] , \IDinst/RegFile[16][8] ,
         \IDinst/RegFile[16][7] , \IDinst/RegFile[16][6] ,
         \IDinst/RegFile[16][5] , \IDinst/RegFile[16][4] ,
         \IDinst/RegFile[16][3] , \IDinst/RegFile[16][2] ,
         \IDinst/RegFile[16][1] , \IDinst/RegFile[16][0] ,
         \IDinst/RegFile[17][31] , \IDinst/RegFile[17][30] ,
         \IDinst/RegFile[17][29] , \IDinst/RegFile[17][28] ,
         \IDinst/RegFile[17][27] , \IDinst/RegFile[17][26] ,
         \IDinst/RegFile[17][25] , \IDinst/RegFile[17][24] ,
         \IDinst/RegFile[17][23] , \IDinst/RegFile[17][22] ,
         \IDinst/RegFile[17][21] , \IDinst/RegFile[17][20] ,
         \IDinst/RegFile[17][19] , \IDinst/RegFile[17][18] ,
         \IDinst/RegFile[17][17] , \IDinst/RegFile[17][16] ,
         \IDinst/RegFile[17][15] , \IDinst/RegFile[17][14] ,
         \IDinst/RegFile[17][13] , \IDinst/RegFile[17][12] ,
         \IDinst/RegFile[17][11] , \IDinst/RegFile[17][10] ,
         \IDinst/RegFile[17][9] , \IDinst/RegFile[17][8] ,
         \IDinst/RegFile[17][7] , \IDinst/RegFile[17][6] ,
         \IDinst/RegFile[17][5] , \IDinst/RegFile[17][4] ,
         \IDinst/RegFile[17][3] , \IDinst/RegFile[17][2] ,
         \IDinst/RegFile[17][1] , \IDinst/RegFile[17][0] ,
         \IDinst/RegFile[18][31] , \IDinst/RegFile[18][30] ,
         \IDinst/RegFile[18][29] , \IDinst/RegFile[18][28] ,
         \IDinst/RegFile[18][27] , \IDinst/RegFile[18][26] ,
         \IDinst/RegFile[18][25] , \IDinst/RegFile[18][24] ,
         \IDinst/RegFile[18][23] , \IDinst/RegFile[18][22] ,
         \IDinst/RegFile[18][21] , \IDinst/RegFile[18][20] ,
         \IDinst/RegFile[18][19] , \IDinst/RegFile[18][18] ,
         \IDinst/RegFile[18][17] , \IDinst/RegFile[18][16] ,
         \IDinst/RegFile[18][15] , \IDinst/RegFile[18][14] ,
         \IDinst/RegFile[18][13] , \IDinst/RegFile[18][12] ,
         \IDinst/RegFile[18][11] , \IDinst/RegFile[18][10] ,
         \IDinst/RegFile[18][9] , \IDinst/RegFile[18][8] ,
         \IDinst/RegFile[18][7] , \IDinst/RegFile[18][6] ,
         \IDinst/RegFile[18][5] , \IDinst/RegFile[18][4] ,
         \IDinst/RegFile[18][3] , \IDinst/RegFile[18][2] ,
         \IDinst/RegFile[18][1] , \IDinst/RegFile[18][0] ,
         \IDinst/RegFile[19][31] , \IDinst/RegFile[19][30] ,
         \IDinst/RegFile[19][29] , \IDinst/RegFile[19][28] ,
         \IDinst/RegFile[19][27] , \IDinst/RegFile[19][26] ,
         \IDinst/RegFile[19][25] , \IDinst/RegFile[19][24] ,
         \IDinst/RegFile[19][23] , \IDinst/RegFile[19][22] ,
         \IDinst/RegFile[19][21] , \IDinst/RegFile[19][20] ,
         \IDinst/RegFile[19][19] , \IDinst/RegFile[19][18] ,
         \IDinst/RegFile[19][17] , \IDinst/RegFile[19][16] ,
         \IDinst/RegFile[19][15] , \IDinst/RegFile[19][14] ,
         \IDinst/RegFile[19][13] , \IDinst/RegFile[19][12] ,
         \IDinst/RegFile[19][11] , \IDinst/RegFile[19][10] ,
         \IDinst/RegFile[19][9] , \IDinst/RegFile[19][8] ,
         \IDinst/RegFile[19][7] , \IDinst/RegFile[19][6] ,
         \IDinst/RegFile[19][5] , \IDinst/RegFile[19][4] ,
         \IDinst/RegFile[19][3] , \IDinst/RegFile[19][2] ,
         \IDinst/RegFile[19][1] , \IDinst/RegFile[19][0] ,
         \IDinst/RegFile[20][31] , \IDinst/RegFile[20][30] ,
         \IDinst/RegFile[20][29] , \IDinst/RegFile[20][28] ,
         \IDinst/RegFile[20][27] , \IDinst/RegFile[20][26] ,
         \IDinst/RegFile[20][25] , \IDinst/RegFile[20][24] ,
         \IDinst/RegFile[20][23] , \IDinst/RegFile[20][22] ,
         \IDinst/RegFile[20][21] , \IDinst/RegFile[20][20] ,
         \IDinst/RegFile[20][19] , \IDinst/RegFile[20][18] ,
         \IDinst/RegFile[20][17] , \IDinst/RegFile[20][16] ,
         \IDinst/RegFile[20][15] , \IDinst/RegFile[20][14] ,
         \IDinst/RegFile[20][13] , \IDinst/RegFile[20][12] ,
         \IDinst/RegFile[20][11] , \IDinst/RegFile[20][10] ,
         \IDinst/RegFile[20][9] , \IDinst/RegFile[20][8] ,
         \IDinst/RegFile[20][7] , \IDinst/RegFile[20][6] ,
         \IDinst/RegFile[20][5] , \IDinst/RegFile[20][4] ,
         \IDinst/RegFile[20][3] , \IDinst/RegFile[20][2] ,
         \IDinst/RegFile[20][1] , \IDinst/RegFile[20][0] ,
         \IDinst/RegFile[21][31] , \IDinst/RegFile[21][30] ,
         \IDinst/RegFile[21][29] , \IDinst/RegFile[21][28] ,
         \IDinst/RegFile[21][27] , \IDinst/RegFile[21][26] ,
         \IDinst/RegFile[21][25] , \IDinst/RegFile[21][24] ,
         \IDinst/RegFile[21][23] , \IDinst/RegFile[21][22] ,
         \IDinst/RegFile[21][21] , \IDinst/RegFile[21][20] ,
         \IDinst/RegFile[21][19] , \IDinst/RegFile[21][18] ,
         \IDinst/RegFile[21][17] , \IDinst/RegFile[21][16] ,
         \IDinst/RegFile[21][15] , \IDinst/RegFile[21][14] ,
         \IDinst/RegFile[21][13] , \IDinst/RegFile[21][12] ,
         \IDinst/RegFile[21][11] , \IDinst/RegFile[21][10] ,
         \IDinst/RegFile[21][9] , \IDinst/RegFile[21][8] ,
         \IDinst/RegFile[21][7] , \IDinst/RegFile[21][6] ,
         \IDinst/RegFile[21][5] , \IDinst/RegFile[21][4] ,
         \IDinst/RegFile[21][3] , \IDinst/RegFile[21][2] ,
         \IDinst/RegFile[21][1] , \IDinst/RegFile[21][0] ,
         \IDinst/RegFile[22][31] , \IDinst/RegFile[22][30] ,
         \IDinst/RegFile[22][29] , \IDinst/RegFile[22][28] ,
         \IDinst/RegFile[22][27] , \IDinst/RegFile[22][26] ,
         \IDinst/RegFile[22][25] , \IDinst/RegFile[22][24] ,
         \IDinst/RegFile[22][23] , \IDinst/RegFile[22][22] ,
         \IDinst/RegFile[22][21] , \IDinst/RegFile[22][20] ,
         \IDinst/RegFile[22][19] , \IDinst/RegFile[22][18] ,
         \IDinst/RegFile[22][17] , \IDinst/RegFile[22][16] ,
         \IDinst/RegFile[22][15] , \IDinst/RegFile[22][14] ,
         \IDinst/RegFile[22][13] , \IDinst/RegFile[22][12] ,
         \IDinst/RegFile[22][11] , \IDinst/RegFile[22][10] ,
         \IDinst/RegFile[22][9] , \IDinst/RegFile[22][8] ,
         \IDinst/RegFile[22][7] , \IDinst/RegFile[22][6] ,
         \IDinst/RegFile[22][5] , \IDinst/RegFile[22][4] ,
         \IDinst/RegFile[22][3] , \IDinst/RegFile[22][2] ,
         \IDinst/RegFile[22][1] , \IDinst/RegFile[22][0] ,
         \IDinst/RegFile[23][31] , \IDinst/RegFile[23][30] ,
         \IDinst/RegFile[23][29] , \IDinst/RegFile[23][28] ,
         \IDinst/RegFile[23][27] , \IDinst/RegFile[23][26] ,
         \IDinst/RegFile[23][25] , \IDinst/RegFile[23][24] ,
         \IDinst/RegFile[23][23] , \IDinst/RegFile[23][22] ,
         \IDinst/RegFile[23][21] , \IDinst/RegFile[23][20] ,
         \IDinst/RegFile[23][19] , \IDinst/RegFile[23][18] ,
         \IDinst/RegFile[23][17] , \IDinst/RegFile[23][16] ,
         \IDinst/RegFile[23][15] , \IDinst/RegFile[23][14] ,
         \IDinst/RegFile[23][13] , \IDinst/RegFile[23][12] ,
         \IDinst/RegFile[23][11] , \IDinst/RegFile[23][10] ,
         \IDinst/RegFile[23][9] , \IDinst/RegFile[23][8] ,
         \IDinst/RegFile[23][7] , \IDinst/RegFile[23][6] ,
         \IDinst/RegFile[23][5] , \IDinst/RegFile[23][4] ,
         \IDinst/RegFile[23][3] , \IDinst/RegFile[23][2] ,
         \IDinst/RegFile[23][1] , \IDinst/RegFile[23][0] ,
         \IDinst/RegFile[24][31] , \IDinst/RegFile[24][30] ,
         \IDinst/RegFile[24][29] , \IDinst/RegFile[24][28] ,
         \IDinst/RegFile[24][27] , \IDinst/RegFile[24][26] ,
         \IDinst/RegFile[24][25] , \IDinst/RegFile[24][24] ,
         \IDinst/RegFile[24][23] , \IDinst/RegFile[24][22] ,
         \IDinst/RegFile[24][21] , \IDinst/RegFile[24][20] ,
         \IDinst/RegFile[24][19] , \IDinst/RegFile[24][18] ,
         \IDinst/RegFile[24][17] , \IDinst/RegFile[24][16] ,
         \IDinst/RegFile[24][15] , \IDinst/RegFile[24][14] ,
         \IDinst/RegFile[24][13] , \IDinst/RegFile[24][12] ,
         \IDinst/RegFile[24][11] , \IDinst/RegFile[24][10] ,
         \IDinst/RegFile[24][9] , \IDinst/RegFile[24][8] ,
         \IDinst/RegFile[24][7] , \IDinst/RegFile[24][6] ,
         \IDinst/RegFile[24][5] , \IDinst/RegFile[24][4] ,
         \IDinst/RegFile[24][3] , \IDinst/RegFile[24][2] ,
         \IDinst/RegFile[24][1] , \IDinst/RegFile[24][0] ,
         \IDinst/RegFile[25][31] , \IDinst/RegFile[25][30] ,
         \IDinst/RegFile[25][29] , \IDinst/RegFile[25][28] ,
         \IDinst/RegFile[25][27] , \IDinst/RegFile[25][26] ,
         \IDinst/RegFile[25][25] , \IDinst/RegFile[25][24] ,
         \IDinst/RegFile[25][23] , \IDinst/RegFile[25][22] ,
         \IDinst/RegFile[25][21] , \IDinst/RegFile[25][20] ,
         \IDinst/RegFile[25][19] , \IDinst/RegFile[25][18] ,
         \IDinst/RegFile[25][17] , \IDinst/RegFile[25][16] ,
         \IDinst/RegFile[25][15] , \IDinst/RegFile[25][14] ,
         \IDinst/RegFile[25][13] , \IDinst/RegFile[25][12] ,
         \IDinst/RegFile[25][11] , \IDinst/RegFile[25][10] ,
         \IDinst/RegFile[25][9] , \IDinst/RegFile[25][8] ,
         \IDinst/RegFile[25][7] , \IDinst/RegFile[25][6] ,
         \IDinst/RegFile[25][5] , \IDinst/RegFile[25][4] ,
         \IDinst/RegFile[25][3] , \IDinst/RegFile[25][2] ,
         \IDinst/RegFile[25][1] , \IDinst/RegFile[25][0] ,
         \IDinst/RegFile[26][31] , \IDinst/RegFile[26][30] ,
         \IDinst/RegFile[26][29] , \IDinst/RegFile[26][28] ,
         \IDinst/RegFile[26][27] , \IDinst/RegFile[26][26] ,
         \IDinst/RegFile[26][25] , \IDinst/RegFile[26][24] ,
         \IDinst/RegFile[26][23] , \IDinst/RegFile[26][22] ,
         \IDinst/RegFile[26][21] , \IDinst/RegFile[26][20] ,
         \IDinst/RegFile[26][19] , \IDinst/RegFile[26][18] ,
         \IDinst/RegFile[26][17] , \IDinst/RegFile[26][16] ,
         \IDinst/RegFile[26][15] , \IDinst/RegFile[26][14] ,
         \IDinst/RegFile[26][13] , \IDinst/RegFile[26][12] ,
         \IDinst/RegFile[26][11] , \IDinst/RegFile[26][10] ,
         \IDinst/RegFile[26][9] , \IDinst/RegFile[26][8] ,
         \IDinst/RegFile[26][7] , \IDinst/RegFile[26][6] ,
         \IDinst/RegFile[26][5] , \IDinst/RegFile[26][4] ,
         \IDinst/RegFile[26][3] , \IDinst/RegFile[26][2] ,
         \IDinst/RegFile[26][1] , \IDinst/RegFile[26][0] ,
         \IDinst/RegFile[27][31] , \IDinst/RegFile[27][30] ,
         \IDinst/RegFile[27][29] , \IDinst/RegFile[27][28] ,
         \IDinst/RegFile[27][27] , \IDinst/RegFile[27][26] ,
         \IDinst/RegFile[27][25] , \IDinst/RegFile[27][24] ,
         \IDinst/RegFile[27][23] , \IDinst/RegFile[27][22] ,
         \IDinst/RegFile[27][21] , \IDinst/RegFile[27][20] ,
         \IDinst/RegFile[27][19] , \IDinst/RegFile[27][18] ,
         \IDinst/RegFile[27][17] , \IDinst/RegFile[27][16] ,
         \IDinst/RegFile[27][15] , \IDinst/RegFile[27][14] ,
         \IDinst/RegFile[27][13] , \IDinst/RegFile[27][12] ,
         \IDinst/RegFile[27][11] , \IDinst/RegFile[27][10] ,
         \IDinst/RegFile[27][9] , \IDinst/RegFile[27][8] ,
         \IDinst/RegFile[27][7] , \IDinst/RegFile[27][6] ,
         \IDinst/RegFile[27][5] , \IDinst/RegFile[27][4] ,
         \IDinst/RegFile[27][3] , \IDinst/RegFile[27][2] ,
         \IDinst/RegFile[27][1] , \IDinst/RegFile[27][0] ,
         \IDinst/RegFile[28][31] , \IDinst/RegFile[28][30] ,
         \IDinst/RegFile[28][29] , \IDinst/RegFile[28][28] ,
         \IDinst/RegFile[28][27] , \IDinst/RegFile[28][26] ,
         \IDinst/RegFile[28][25] , \IDinst/RegFile[28][24] ,
         \IDinst/RegFile[28][23] , \IDinst/RegFile[28][22] ,
         \IDinst/RegFile[28][21] , \IDinst/RegFile[28][20] ,
         \IDinst/RegFile[28][19] , \IDinst/RegFile[28][18] ,
         \IDinst/RegFile[28][17] , \IDinst/RegFile[28][16] ,
         \IDinst/RegFile[28][15] , \IDinst/RegFile[28][14] ,
         \IDinst/RegFile[28][13] , \IDinst/RegFile[28][12] ,
         \IDinst/RegFile[28][11] , \IDinst/RegFile[28][10] ,
         \IDinst/RegFile[28][9] , \IDinst/RegFile[28][8] ,
         \IDinst/RegFile[28][7] , \IDinst/RegFile[28][6] ,
         \IDinst/RegFile[28][5] , \IDinst/RegFile[28][4] ,
         \IDinst/RegFile[28][3] , \IDinst/RegFile[28][2] ,
         \IDinst/RegFile[28][1] , \IDinst/RegFile[28][0] ,
         \IDinst/RegFile[29][31] , \IDinst/RegFile[29][30] ,
         \IDinst/RegFile[29][29] , \IDinst/RegFile[29][28] ,
         \IDinst/RegFile[29][27] , \IDinst/RegFile[29][26] ,
         \IDinst/RegFile[29][25] , \IDinst/RegFile[29][24] ,
         \IDinst/RegFile[29][23] , \IDinst/RegFile[29][22] ,
         \IDinst/RegFile[29][21] , \IDinst/RegFile[29][20] ,
         \IDinst/RegFile[29][19] , \IDinst/RegFile[29][18] ,
         \IDinst/RegFile[29][17] , \IDinst/RegFile[29][16] ,
         \IDinst/RegFile[29][15] , \IDinst/RegFile[29][14] ,
         \IDinst/RegFile[29][13] , \IDinst/RegFile[29][12] ,
         \IDinst/RegFile[29][11] , \IDinst/RegFile[29][10] ,
         \IDinst/RegFile[29][9] , \IDinst/RegFile[29][8] ,
         \IDinst/RegFile[29][7] , \IDinst/RegFile[29][6] ,
         \IDinst/RegFile[29][5] , \IDinst/RegFile[29][4] ,
         \IDinst/RegFile[29][3] , \IDinst/RegFile[29][2] ,
         \IDinst/RegFile[29][1] , \IDinst/RegFile[29][0] ,
         \IDinst/RegFile[30][31] , \IDinst/RegFile[30][30] ,
         \IDinst/RegFile[30][29] , \IDinst/RegFile[30][28] ,
         \IDinst/RegFile[30][27] , \IDinst/RegFile[30][26] ,
         \IDinst/RegFile[30][25] , \IDinst/RegFile[30][24] ,
         \IDinst/RegFile[30][23] , \IDinst/RegFile[30][22] ,
         \IDinst/RegFile[30][21] , \IDinst/RegFile[30][20] ,
         \IDinst/RegFile[30][19] , \IDinst/RegFile[30][18] ,
         \IDinst/RegFile[30][17] , \IDinst/RegFile[30][16] ,
         \IDinst/RegFile[30][15] , \IDinst/RegFile[30][14] ,
         \IDinst/RegFile[30][13] , \IDinst/RegFile[30][12] ,
         \IDinst/RegFile[30][11] , \IDinst/RegFile[30][10] ,
         \IDinst/RegFile[30][9] , \IDinst/RegFile[30][8] ,
         \IDinst/RegFile[30][7] , \IDinst/RegFile[30][6] ,
         \IDinst/RegFile[30][5] , \IDinst/RegFile[30][4] ,
         \IDinst/RegFile[30][3] , \IDinst/RegFile[30][2] ,
         \IDinst/RegFile[30][1] , \IDinst/RegFile[30][0] ,
         \IDinst/RegFile[31][31] , \IDinst/RegFile[31][30] ,
         \IDinst/RegFile[31][29] , \IDinst/RegFile[31][28] ,
         \IDinst/RegFile[31][27] , \IDinst/RegFile[31][26] ,
         \IDinst/RegFile[31][25] , \IDinst/RegFile[31][24] ,
         \IDinst/RegFile[31][23] , \IDinst/RegFile[31][22] ,
         \IDinst/RegFile[31][21] , \IDinst/RegFile[31][20] ,
         \IDinst/RegFile[31][19] , \IDinst/RegFile[31][18] ,
         \IDinst/RegFile[31][17] , \IDinst/RegFile[31][16] ,
         \IDinst/RegFile[31][15] , \IDinst/RegFile[31][14] ,
         \IDinst/RegFile[31][13] , \IDinst/RegFile[31][12] ,
         \IDinst/RegFile[31][11] , \IDinst/RegFile[31][10] ,
         \IDinst/RegFile[31][9] , \IDinst/RegFile[31][8] ,
         \IDinst/RegFile[31][7] , \IDinst/RegFile[31][6] ,
         \IDinst/RegFile[31][5] , \IDinst/RegFile[31][4] ,
         \IDinst/RegFile[31][3] , \IDinst/RegFile[31][2] ,
         \IDinst/RegFile[31][1] , \IDinst/RegFile[31][0] , \IDinst/N48 ,
         \IDinst/N46 , \IDinst/N45 , \IDinst/N44 , \IDinst/N43 , \IDinst/N41 ,
         \IDinst/N40 , \IDinst/N39 , \EXinst/n1463 , \EXinst/n1462 ,
         \EXinst/n1461 , \EXinst/n1460 , \EXinst/n1459 , \EXinst/n1458 ,
         \EXinst/n1457 , \EXinst/n1456 , \EXinst/n1455 , \EXinst/n1454 ,
         \EXinst/n1453 , \EXinst/n1452 , \EXinst/n1451 , \EXinst/n1450 ,
         \EXinst/n1449 , \EXinst/n1448 , \EXinst/n1447 , \EXinst/n1446 ,
         \EXinst/n1445 , \EXinst/n1444 , \EXinst/n1443 , \EXinst/n1442 ,
         \EXinst/n1441 , \EXinst/n1440 , \EXinst/n1439 , \EXinst/n1438 ,
         \EXinst/n1437 , \EXinst/n1436 , \EXinst/n1435 , \EXinst/n1434 ,
         \EXinst/n1433 , \EXinst/n1432 , \EXinst/n1423 , \EXinst/n1387 ,
         \EXinst/N1341 , \EXinst/N1340 , \EXinst/N1339 , \EXinst/N1338 ,
         \EXinst/N1337 , \EXinst/N1336 , \EXinst/N1335 , \EXinst/N1334 ,
         \EXinst/N1333 , \EXinst/N1332 , \EXinst/N1331 , \EXinst/N1330 ,
         \EXinst/N1329 , \EXinst/N1328 , \EXinst/N1327 , \EXinst/N1326 ,
         \EXinst/N1325 , \EXinst/N1324 , \EXinst/N1323 , \EXinst/N1322 ,
         \EXinst/N1321 , \EXinst/N1320 , \EXinst/N1319 , \EXinst/N1318 ,
         \EXinst/N1317 , \EXinst/N1316 , \EXinst/N1315 , \EXinst/N1314 ,
         \EXinst/N1313 , \EXinst/N1312 , \EXinst/N1311 , \EXinst/N1310 ,
         \EXinst/N1309 , \EXinst/N1308 , \EXinst/N1307 , \EXinst/N1306 ,
         \EXinst/N1305 , \MEMinst/N88 , \MEMinst/N87 , \MEMinst/N86 ,
         \MEMinst/N85 , \MEMinst/N84 , \MEMinst/N83 , \MEMinst/N82 ,
         \MEMinst/N81 , \MEMinst/N80 , \MEMinst/N79 , \MEMinst/N78 ,
         \MEMinst/N77 , \MEMinst/N76 , \MEMinst/N75 , \MEMinst/N74 ,
         \MEMinst/N73 , \MEMinst/N72 , \MEMinst/N71 , \MEMinst/N70 ,
         \MEMinst/N69 , \MEMinst/N68 , \MEMinst/N67 , \MEMinst/N66 ,
         \MEMinst/N65 , \MEMinst/N64 , \MEMinst/N63 , \MEMinst/N62 ,
         \MEMinst/N61 , \MEMinst/N60 , \MEMinst/N59 , \MEMinst/N58 ,
         \MEMinst/N57 , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588;

  assign \NPC[1]  = \IFinst/N8 ;
  assign \NPC[0]  = \IFinst/N7 ;

  dffascs1 \IFinst/IR_previous_reg[0]  ( .DIN(\IFinst/n591 ), .CLK(clk), 
        .CLRB(n1018), .SETB(1'b1), .Q(n9587) );
  dffascs1 \IFinst/IR_latched_reg[0]  ( .DIN(\IFinst/N104 ), .CLK(clk), 
        .CLRB(n1018), .SETB(1'b1), .Q(n41), .QN(n9384) );
  dffascs1 \IFinst/IR_curr_reg[0]  ( .DIN(\IFinst/n594 ), .CLK(clk), 
        .CLRB(n962), .SETB(1'b1), .Q(n9586) );
  dffascs1 \IFinst/IR_previous_reg[1]  ( .DIN(\IFinst/n596 ), .CLK(clk), 
        .CLRB(n958), .SETB(1'b1), .Q(n9585) );
  dffascs1 \IFinst/IR_latched_reg[1]  ( .DIN(\IFinst/N105 ), .CLK(clk), 
        .CLRB(n958), .SETB(1'b1), .Q(n42), .QN(n9388) );
  dffascs1 \IFinst/IR_curr_reg[1]  ( .DIN(\IFinst/n599 ), .CLK(clk), 
        .CLRB(n961), .SETB(1'b1), .Q(n9584) );
  dffascs1 \IFinst/IR_previous_reg[2]  ( .DIN(\IFinst/n601 ), .CLK(clk), 
        .CLRB(n958), .SETB(1'b1), .Q(n9583) );
  dffascs1 \IFinst/IR_latched_reg[2]  ( .DIN(\IFinst/N106 ), .CLK(clk), 
        .CLRB(n958), .SETB(1'b1), .Q(n100) );
  dffascs1 \IFinst/IR_curr_reg[2]  ( .DIN(\IFinst/n604 ), .CLK(clk), 
        .CLRB(n961), .SETB(1'b1), .Q(n9582) );
  dffascs1 \IFinst/IR_previous_reg[3]  ( .DIN(\IFinst/n606 ), .CLK(clk), 
        .CLRB(n957), .SETB(1'b1), .Q(n9581) );
  dffascs1 \IFinst/IR_latched_reg[3]  ( .DIN(\IFinst/N107 ), .CLK(clk), 
        .CLRB(n957), .SETB(1'b1), .Q(n116), .QN(n9389) );
  dffascs1 \IFinst/IR_curr_reg[3]  ( .DIN(\IFinst/n609 ), .CLK(clk), 
        .CLRB(n961), .SETB(1'b1), .Q(n9580) );
  dffascs1 \IFinst/IR_previous_reg[4]  ( .DIN(\IFinst/n611 ), .CLK(clk), 
        .CLRB(n957), .SETB(1'b1), .Q(n9579) );
  dffascs1 \IFinst/IR_latched_reg[4]  ( .DIN(\IFinst/N108 ), .CLK(clk), 
        .CLRB(n957), .SETB(1'b1), .Q(n99) );
  dffascs1 \IFinst/IR_curr_reg[4]  ( .DIN(\IFinst/n614 ), .CLK(clk), 
        .CLRB(n961), .SETB(1'b1), .Q(n9578) );
  dffascs1 \IFinst/IR_previous_reg[5]  ( .DIN(\IFinst/n616 ), .CLK(clk), 
        .CLRB(n957), .SETB(1'b1), .Q(n9577) );
  dffascs1 \IFinst/IR_latched_reg[5]  ( .DIN(\IFinst/N109 ), .CLK(clk), 
        .CLRB(n957), .SETB(1'b1), .Q(n115), .QN(n9390) );
  dffascs1 \IFinst/IR_curr_reg[5]  ( .DIN(\IFinst/n619 ), .CLK(clk), 
        .CLRB(n961), .SETB(1'b1), .Q(n9576) );
  dffascs1 \IFinst/IR_previous_reg[6]  ( .DIN(\IFinst/n621 ), .CLK(clk), 
        .CLRB(n957), .SETB(1'b1), .Q(n9575) );
  dffascs1 \IFinst/IR_latched_reg[6]  ( .DIN(\IFinst/N110 ), .CLK(clk), 
        .CLRB(n957), .SETB(1'b1), .Q(n112) );
  dffascs1 \IFinst/IR_curr_reg[6]  ( .DIN(\IFinst/n624 ), .CLK(clk), 
        .CLRB(n961), .SETB(1'b1), .Q(n9574) );
  dffascs1 \IFinst/IR_previous_reg[7]  ( .DIN(\IFinst/n626 ), .CLK(clk), 
        .CLRB(n957), .SETB(1'b1), .Q(n9573) );
  dffascs1 \IFinst/IR_latched_reg[7]  ( .DIN(\IFinst/N111 ), .CLK(clk), 
        .CLRB(n957), .SETB(1'b1), .Q(n126), .QN(n9391) );
  dffascs1 \IFinst/IR_curr_reg[7]  ( .DIN(\IFinst/n629 ), .CLK(clk), 
        .CLRB(n961), .SETB(1'b1), .Q(n9572) );
  dffascs1 \IFinst/IR_previous_reg[8]  ( .DIN(\IFinst/n631 ), .CLK(clk), 
        .CLRB(n956), .SETB(1'b1), .Q(n9571) );
  dffascs1 \IFinst/IR_latched_reg[8]  ( .DIN(\IFinst/N112 ), .CLK(clk), 
        .CLRB(n956), .SETB(1'b1), .Q(n111) );
  dffascs1 \IFinst/IR_curr_reg[8]  ( .DIN(\IFinst/n634 ), .CLK(clk), 
        .CLRB(n961), .SETB(1'b1), .Q(n9570) );
  dffascs1 \IFinst/IR_previous_reg[9]  ( .DIN(\IFinst/n636 ), .CLK(clk), 
        .CLRB(n956), .SETB(1'b1), .Q(n9569) );
  dffascs1 \IFinst/IR_latched_reg[9]  ( .DIN(\IFinst/N113 ), .CLK(clk), 
        .CLRB(n956), .SETB(1'b1), .Q(n125), .QN(n9392) );
  dffascs1 \IFinst/IR_curr_reg[9]  ( .DIN(\IFinst/n639 ), .CLK(clk), 
        .CLRB(n961), .SETB(1'b1), .Q(n9568) );
  dffascs1 \IFinst/IR_previous_reg[10]  ( .DIN(\IFinst/n641 ), .CLK(clk), 
        .CLRB(n956), .SETB(1'b1), .Q(n9567) );
  dffascs1 \IFinst/IR_latched_reg[10]  ( .DIN(\IFinst/N114 ), .CLK(clk), 
        .CLRB(n956), .SETB(1'b1), .Q(n110) );
  dffascs1 \IFinst/IR_curr_reg[10]  ( .DIN(\IFinst/n644 ), .CLK(clk), 
        .CLRB(n961), .SETB(1'b1), .Q(n9566) );
  dffascs1 \IFinst/IR_previous_reg[11]  ( .DIN(\IFinst/n646 ), .CLK(clk), 
        .CLRB(n956), .SETB(1'b1), .Q(n9565) );
  dffascs1 \IFinst/IR_latched_reg[11]  ( .DIN(\IFinst/N115 ), .CLK(clk), 
        .CLRB(n956), .SETB(1'b1), .Q(n114), .QN(n9385) );
  dffascs1 \IFinst/IR_curr_reg[11]  ( .DIN(\IFinst/n649 ), .CLK(clk), 
        .CLRB(n960), .SETB(1'b1), .Q(n9564) );
  dffascs1 \IFinst/IR_previous_reg[12]  ( .DIN(\IFinst/n651 ), .CLK(clk), 
        .CLRB(n956), .SETB(1'b1), .Q(n9563) );
  dffascs1 \IFinst/IR_latched_reg[12]  ( .DIN(\IFinst/N116 ), .CLK(clk), 
        .CLRB(n956), .SETB(1'b1), .Q(n98) );
  dffascs1 \IFinst/IR_curr_reg[12]  ( .DIN(\IFinst/n654 ), .CLK(clk), 
        .CLRB(n960), .SETB(1'b1), .Q(n9562) );
  dffascs1 \IFinst/IR_previous_reg[13]  ( .DIN(\IFinst/n656 ), .CLK(clk), 
        .CLRB(n955), .SETB(1'b1), .Q(n9561) );
  dffascs1 \IFinst/IR_latched_reg[13]  ( .DIN(\IFinst/N117 ), .CLK(clk), 
        .CLRB(n955), .SETB(1'b1), .Q(n113), .QN(n9386) );
  dffascs1 \IFinst/IR_curr_reg[13]  ( .DIN(\IFinst/n659 ), .CLK(clk), 
        .CLRB(n960), .SETB(1'b1), .Q(n9560) );
  dffascs1 \IFinst/IR_previous_reg[14]  ( .DIN(\IFinst/n661 ), .CLK(clk), 
        .CLRB(n955), .SETB(1'b1), .Q(n9559) );
  dffascs1 \IFinst/IR_latched_reg[14]  ( .DIN(\IFinst/N118 ), .CLK(clk), 
        .CLRB(n955), .SETB(1'b1), .Q(n97) );
  dffascs1 \IFinst/IR_curr_reg[14]  ( .DIN(\IFinst/n664 ), .CLK(clk), 
        .CLRB(n960), .SETB(1'b1), .Q(n9558) );
  dffascs1 \IFinst/IR_previous_reg[15]  ( .DIN(\IFinst/n666 ), .CLK(clk), 
        .CLRB(n955), .SETB(1'b1), .Q(n9557) );
  dffascs1 \IFinst/IR_latched_reg[15]  ( .DIN(\IFinst/N119 ), .CLK(clk), 
        .CLRB(n955), .SETB(1'b1), .Q(n92), .QN(n9387) );
  dffascs1 \IFinst/IR_curr_reg[15]  ( .DIN(\IFinst/n669 ), .CLK(clk), 
        .CLRB(n960), .SETB(1'b1), .Q(n9556) );
  dffascs1 \IFinst/IR_previous_reg[16]  ( .DIN(\IFinst/n671 ), .CLK(clk), 
        .CLRB(n955), .SETB(1'b1), .Q(n9555) );
  dffascs1 \IFinst/IR_latched_reg[16]  ( .DIN(\IFinst/N120 ), .CLK(clk), 
        .CLRB(n955), .SETB(1'b1), .Q(n272) );
  dffascs1 \IFinst/IR_curr_reg[16]  ( .DIN(\IFinst/n674 ), .CLK(clk), 
        .CLRB(n960), .SETB(1'b1), .Q(n9554) );
  dffascs1 \IFinst/IR_previous_reg[17]  ( .DIN(\IFinst/n676 ), .CLK(clk), 
        .CLRB(n954), .SETB(1'b1), .Q(n9553) );
  dffascs1 \IFinst/IR_latched_reg[17]  ( .DIN(\IFinst/N121 ), .CLK(clk), 
        .CLRB(n955), .SETB(1'b1), .Q(n274) );
  dffascs1 \IFinst/IR_curr_reg[17]  ( .DIN(\IFinst/n679 ), .CLK(clk), 
        .CLRB(n960), .SETB(1'b1), .Q(n9552) );
  dffascs1 \IFinst/IR_previous_reg[18]  ( .DIN(\IFinst/n681 ), .CLK(clk), 
        .CLRB(n954), .SETB(1'b1), .Q(n9551) );
  dffascs1 \IFinst/IR_latched_reg[18]  ( .DIN(\IFinst/N122 ), .CLK(clk), 
        .CLRB(n954), .SETB(1'b1), .Q(n278) );
  dffascs1 \IFinst/IR_curr_reg[18]  ( .DIN(\IFinst/n684 ), .CLK(clk), 
        .CLRB(n960), .SETB(1'b1), .Q(n9550) );
  dffascs1 \IFinst/IR_previous_reg[19]  ( .DIN(\IFinst/n686 ), .CLK(clk), 
        .CLRB(n954), .SETB(1'b1), .Q(n9549) );
  dffascs1 \IFinst/IR_latched_reg[19]  ( .DIN(\IFinst/N123 ), .CLK(clk), 
        .CLRB(n954), .SETB(1'b1), .Q(n280) );
  dffascs1 \IFinst/IR_curr_reg[19]  ( .DIN(\IFinst/n689 ), .CLK(clk), 
        .CLRB(n960), .SETB(1'b1), .Q(n9548) );
  dffascs1 \IFinst/IR_previous_reg[20]  ( .DIN(\IFinst/n691 ), .CLK(clk), 
        .CLRB(n953), .SETB(1'b1), .Q(n9547) );
  dffascs1 \IFinst/IR_latched_reg[20]  ( .DIN(\IFinst/N124 ), .CLK(clk), 
        .CLRB(n954), .SETB(1'b1), .Q(n276) );
  dffascs1 \IFinst/IR_curr_reg[20]  ( .DIN(\IFinst/n694 ), .CLK(clk), 
        .CLRB(n960), .SETB(1'b1), .Q(n9546) );
  dffascs1 \IFinst/IR_previous_reg[21]  ( .DIN(\IFinst/n696 ), .CLK(clk), 
        .CLRB(n953), .SETB(1'b1), .Q(n9545) );
  dffascs1 \IFinst/IR_latched_reg[21]  ( .DIN(\IFinst/N125 ), .CLK(clk), 
        .CLRB(n953), .SETB(1'b1), .Q(n308) );
  dffascs1 \IFinst/IR_curr_reg[21]  ( .DIN(\IFinst/n699 ), .CLK(clk), 
        .CLRB(n959), .SETB(1'b1), .Q(n9544) );
  dffascs1 \IFinst/IR_previous_reg[22]  ( .DIN(\IFinst/n701 ), .CLK(clk), 
        .CLRB(n953), .SETB(1'b1), .Q(n9543) );
  dffascs1 \IFinst/IR_latched_reg[22]  ( .DIN(\IFinst/N126 ), .CLK(clk), 
        .CLRB(n953), .SETB(1'b1), .Q(n306) );
  dffascs1 \IFinst/IR_curr_reg[22]  ( .DIN(\IFinst/n704 ), .CLK(clk), 
        .CLRB(n959), .SETB(1'b1), .Q(n9542) );
  dffascs1 \IFinst/IR_previous_reg[23]  ( .DIN(\IFinst/n706 ), .CLK(clk), 
        .CLRB(n953), .SETB(1'b1), .Q(n9541) );
  dffascs1 \IFinst/IR_latched_reg[23]  ( .DIN(\IFinst/N127 ), .CLK(clk), 
        .CLRB(n953), .SETB(1'b1), .Q(n312) );
  dffascs1 \IFinst/IR_curr_reg[23]  ( .DIN(\IFinst/n709 ), .CLK(clk), 
        .CLRB(n959), .SETB(1'b1), .Q(n9540) );
  dffascs1 \IFinst/IR_previous_reg[24]  ( .DIN(\IFinst/n711 ), .CLK(clk), 
        .CLRB(n952), .SETB(1'b1), .Q(n9539) );
  dffascs1 \IFinst/IR_latched_reg[24]  ( .DIN(\IFinst/N128 ), .CLK(clk), 
        .CLRB(n952), .SETB(1'b1), .Q(n314) );
  dffascs1 \IFinst/IR_curr_reg[24]  ( .DIN(\IFinst/n714 ), .CLK(clk), 
        .CLRB(n959), .SETB(1'b1), .Q(n9538) );
  dffascs1 \IFinst/IR_previous_reg[25]  ( .DIN(\IFinst/n716 ), .CLK(clk), 
        .CLRB(n952), .SETB(1'b1), .Q(n9537) );
  dffascs1 \IFinst/IR_latched_reg[25]  ( .DIN(\IFinst/N129 ), .CLK(clk), 
        .CLRB(n952), .SETB(1'b1), .Q(n310) );
  dffascs1 \IFinst/IR_curr_reg[25]  ( .DIN(\IFinst/n719 ), .CLK(clk), 
        .CLRB(n959), .SETB(1'b1), .Q(n9536) );
  dffascs1 \IFinst/IR_previous_reg[26]  ( .DIN(\IFinst/n721 ), .CLK(clk), 
        .CLRB(n952), .SETB(1'b1), .Q(n9535) );
  dffascs1 \IFinst/IR_latched_reg[26]  ( .DIN(\IFinst/N130 ), .CLK(clk), 
        .CLRB(n952), .SETB(1'b1), .Q(n318) );
  dffascs1 \IFinst/IR_curr_reg[26]  ( .DIN(\IFinst/n724 ), .CLK(clk), 
        .CLRB(n959), .SETB(1'b1), .Q(n9534) );
  dffascs1 \IFinst/IR_previous_reg[27]  ( .DIN(\IFinst/n726 ), .CLK(clk), 
        .CLRB(n951), .SETB(1'b1), .Q(n9533) );
  dffascs1 \IFinst/IR_latched_reg[27]  ( .DIN(\IFinst/N131 ), .CLK(clk), 
        .CLRB(n952), .SETB(1'b1), .Q(n320) );
  dffascs1 \IFinst/IR_curr_reg[27]  ( .DIN(\IFinst/n729 ), .CLK(clk), 
        .CLRB(n959), .SETB(1'b1), .Q(n9532) );
  dffascs1 \IFinst/IR_previous_reg[28]  ( .DIN(\IFinst/n731 ), .CLK(clk), 
        .CLRB(n951), .SETB(1'b1), .Q(n9531) );
  dffascs1 \IFinst/IR_latched_reg[28]  ( .DIN(\IFinst/N132 ), .CLK(clk), 
        .CLRB(n951), .SETB(1'b1), .Q(n324) );
  dffascs1 \IFinst/IR_curr_reg[28]  ( .DIN(\IFinst/n734 ), .CLK(clk), 
        .CLRB(n959), .SETB(1'b1), .Q(n9530) );
  dffascs1 \IFinst/IR_previous_reg[29]  ( .DIN(\IFinst/n736 ), .CLK(clk), 
        .CLRB(n951), .SETB(1'b1), .Q(n9529) );
  dffascs1 \IFinst/IR_latched_reg[29]  ( .DIN(\IFinst/N133 ), .CLK(clk), 
        .CLRB(n951), .SETB(1'b1), .Q(n326) );
  dffascs1 \IFinst/IR_curr_reg[29]  ( .DIN(\IFinst/n739 ), .CLK(clk), 
        .CLRB(n959), .SETB(1'b1), .Q(n9528) );
  dffascs1 \IFinst/IR_previous_reg[30]  ( .DIN(\IFinst/n741 ), .CLK(clk), 
        .CLRB(n926), .SETB(1'b1), .Q(n9527) );
  dffascs1 \IFinst/IR_latched_reg[30]  ( .DIN(\IFinst/N134 ), .CLK(clk), 
        .CLRB(n951), .SETB(1'b1), .Q(n316) );
  dffascs1 \IFinst/IR_curr_reg[30]  ( .DIN(\IFinst/n744 ), .CLK(clk), 
        .CLRB(n959), .SETB(1'b1), .Q(n9526) );
  dffascs1 \IFinst/IR_previous_reg[31]  ( .DIN(\IFinst/n746 ), .CLK(clk), 
        .CLRB(n809), .SETB(1'b1), .Q(n9525) );
  dffascs1 \IFinst/IR_latched_reg[31]  ( .DIN(\IFinst/N135 ), .CLK(clk), 
        .CLRB(n958), .SETB(1'b1), .Q(n322) );
  dffascs1 \IFinst/IR_curr_reg[31]  ( .DIN(\IFinst/n749 ), .CLK(clk), 
        .CLRB(n958), .SETB(1'b1), .Q(n9524) );
  dffascs1 \IFinst/PC_reg[0]  ( .DIN(\IFinst/n847 ), .CLK(clk), .CLRB(n925), 
        .SETB(1'b1), .Q(n9523) );
  dffascs1 \IFinst/PC_reg[31]  ( .DIN(\IFinst/n816 ), .CLK(clk), .CLRB(n809), 
        .SETB(1'b1), .Q(n9522) );
  dffascs1 \IFinst/NPC_reg[31]  ( .DIN(\IFinst/N103 ), .CLK(clk), .CLRB(n918), 
        .SETB(1'b1), .Q(\NPC[31] ), .QN(n9424) );
  dffascs1 \IFinst/PC_reg[30]  ( .DIN(\IFinst/n817 ), .CLK(clk), .CLRB(n830), 
        .SETB(1'b1), .Q(n9521) );
  dffascs1 \IFinst/NPC_reg[30]  ( .DIN(\IFinst/N102 ), .CLK(clk), .CLRB(n830), 
        .SETB(1'b1), .Q(\NPC[30] ), .QN(n9520) );
  dffascs1 \IFinst/PC_reg[29]  ( .DIN(\IFinst/n818 ), .CLK(clk), .CLRB(n831), 
        .SETB(1'b1), .Q(n9519) );
  dffascs1 \IFinst/NPC_reg[29]  ( .DIN(\IFinst/N101 ), .CLK(clk), .CLRB(n831), 
        .SETB(1'b1), .Q(\NPC[29] ), .QN(n9425) );
  dffascs1 \IFinst/PC_reg[28]  ( .DIN(\IFinst/n819 ), .CLK(clk), .CLRB(n809), 
        .SETB(1'b1), .Q(n9518) );
  dffascs1 \IFinst/NPC_reg[28]  ( .DIN(\IFinst/N100 ), .CLK(clk), .CLRB(n918), 
        .SETB(1'b1), .Q(\NPC[28] ), .QN(n9426) );
  dffascs1 \IFinst/PC_reg[27]  ( .DIN(\IFinst/n820 ), .CLK(clk), .CLRB(n810), 
        .SETB(1'b1), .Q(n9517) );
  dffascs1 \IFinst/NPC_reg[27]  ( .DIN(\IFinst/N99 ), .CLK(clk), .CLRB(n906), 
        .SETB(1'b1), .Q(\NPC[27] ), .QN(n9427) );
  dffascs1 \IFinst/PC_reg[26]  ( .DIN(\IFinst/n821 ), .CLK(clk), .CLRB(n812), 
        .SETB(1'b1), .Q(n9516) );
  dffascs1 \IFinst/NPC_reg[26]  ( .DIN(\IFinst/N98 ), .CLK(clk), .CLRB(n879), 
        .SETB(1'b1), .Q(\NPC[26] ), .QN(n9428) );
  dffascs1 \IFinst/PC_reg[25]  ( .DIN(\IFinst/n822 ), .CLK(clk), .CLRB(n810), 
        .SETB(1'b1), .Q(n9515) );
  dffascs1 \IFinst/NPC_reg[25]  ( .DIN(\IFinst/N97 ), .CLK(clk), .CLRB(n899), 
        .SETB(1'b1), .Q(\NPC[25] ), .QN(n9429) );
  dffascs1 \IFinst/PC_reg[24]  ( .DIN(\IFinst/n823 ), .CLK(clk), .CLRB(n812), 
        .SETB(1'b1), .Q(n9514) );
  dffascs1 \IFinst/NPC_reg[24]  ( .DIN(\IFinst/N96 ), .CLK(clk), .CLRB(n880), 
        .SETB(1'b1), .Q(\NPC[24] ), .QN(n9430) );
  dffascs1 \IFinst/PC_reg[23]  ( .DIN(\IFinst/n824 ), .CLK(clk), .CLRB(n811), 
        .SETB(1'b1), .Q(n9513) );
  dffascs1 \IFinst/NPC_reg[23]  ( .DIN(\IFinst/N95 ), .CLK(clk), .CLRB(n888), 
        .SETB(1'b1), .Q(\NPC[23] ), .QN(n9431) );
  dffascs1 \IFinst/PC_reg[22]  ( .DIN(\IFinst/n825 ), .CLK(clk), .CLRB(n812), 
        .SETB(1'b1), .Q(n9512) );
  dffascs1 \IFinst/NPC_reg[22]  ( .DIN(\IFinst/N94 ), .CLK(clk), .CLRB(n880), 
        .SETB(1'b1), .Q(\NPC[22] ), .QN(n9432) );
  dffascs1 \IFinst/PC_reg[21]  ( .DIN(\IFinst/n826 ), .CLK(clk), .CLRB(n811), 
        .SETB(1'b1), .Q(n9511) );
  dffascs1 \IFinst/NPC_reg[21]  ( .DIN(\IFinst/N93 ), .CLK(clk), .CLRB(n884), 
        .SETB(1'b1), .Q(\NPC[21] ), .QN(n9433) );
  dffascs1 \IFinst/PC_reg[20]  ( .DIN(\IFinst/n827 ), .CLK(clk), .CLRB(n811), 
        .SETB(1'b1), .Q(n9510) );
  dffascs1 \IFinst/NPC_reg[20]  ( .DIN(\IFinst/N92 ), .CLK(clk), .CLRB(n884), 
        .SETB(1'b1), .Q(\NPC[20] ), .QN(n9434) );
  dffascs1 \IFinst/PC_reg[19]  ( .DIN(\IFinst/n828 ), .CLK(clk), .CLRB(n813), 
        .SETB(1'b1), .Q(n9509) );
  dffascs1 \IFinst/NPC_reg[19]  ( .DIN(\IFinst/N91 ), .CLK(clk), .CLRB(n872), 
        .SETB(1'b1), .Q(\NPC[19] ), .QN(n9435) );
  dffascs1 \IFinst/PC_reg[18]  ( .DIN(\IFinst/n829 ), .CLK(clk), .CLRB(n813), 
        .SETB(1'b1), .Q(n9508) );
  dffascs1 \IFinst/NPC_reg[18]  ( .DIN(\IFinst/N90 ), .CLK(clk), .CLRB(n872), 
        .SETB(1'b1), .Q(\NPC[18] ), .QN(n9436) );
  dffascs1 \IFinst/PC_reg[17]  ( .DIN(\IFinst/n830 ), .CLK(clk), .CLRB(n810), 
        .SETB(1'b1), .Q(n9507) );
  dffascs1 \IFinst/NPC_reg[17]  ( .DIN(\IFinst/N89 ), .CLK(clk), .CLRB(n913), 
        .SETB(1'b1), .Q(\NPC[17] ), .QN(n9437) );
  dffascs1 \IFinst/PC_reg[16]  ( .DIN(\IFinst/n831 ), .CLK(clk), .CLRB(n809), 
        .SETB(1'b1), .Q(n9506) );
  dffascs1 \IFinst/NPC_reg[16]  ( .DIN(\IFinst/N88 ), .CLK(clk), .CLRB(n914), 
        .SETB(1'b1), .Q(\NPC[16] ), .QN(n9438) );
  dffascs1 \IFinst/PC_reg[15]  ( .DIN(\IFinst/n832 ), .CLK(clk), .CLRB(n820), 
        .SETB(1'b1), .Q(n9505) );
  dffascs1 \IFinst/NPC_reg[15]  ( .DIN(\IFinst/N87 ), .CLK(clk), .CLRB(n864), 
        .SETB(1'b1), .Q(\NPC[15] ), .QN(n9439) );
  dffascs1 \IFinst/PC_reg[14]  ( .DIN(\IFinst/n833 ), .CLK(clk), .CLRB(n820), 
        .SETB(1'b1), .Q(n9504) );
  dffascs1 \IFinst/NPC_reg[14]  ( .DIN(\IFinst/N86 ), .CLK(clk), .CLRB(n864), 
        .SETB(1'b1), .Q(\NPC[14] ), .QN(n9440) );
  dffascs1 \IFinst/PC_reg[13]  ( .DIN(\IFinst/n834 ), .CLK(clk), .CLRB(n812), 
        .SETB(1'b1), .Q(n9503) );
  dffascs1 \IFinst/NPC_reg[13]  ( .DIN(\IFinst/N85 ), .CLK(clk), .CLRB(n876), 
        .SETB(1'b1), .Q(\NPC[13] ), .QN(n9441) );
  dffascs1 \IFinst/PC_reg[12]  ( .DIN(\IFinst/n835 ), .CLK(clk), .CLRB(n831), 
        .SETB(1'b1), .Q(n9502) );
  dffascs1 \IFinst/NPC_reg[12]  ( .DIN(\IFinst/N84 ), .CLK(clk), .CLRB(n831), 
        .SETB(1'b1), .Q(\NPC[12] ), .QN(n9442) );
  dffascs1 \IFinst/PC_reg[11]  ( .DIN(\IFinst/n836 ), .CLK(clk), .CLRB(n828), 
        .SETB(1'b1), .Q(n9501) );
  dffascs1 \IFinst/NPC_reg[11]  ( .DIN(\IFinst/N83 ), .CLK(clk), .CLRB(n856), 
        .SETB(1'b1), .Q(\NPC[11] ), .QN(n9443) );
  dffascs1 \IFinst/PC_reg[10]  ( .DIN(\IFinst/n837 ), .CLK(clk), .CLRB(n828), 
        .SETB(1'b1), .Q(n9500) );
  dffascs1 \IFinst/NPC_reg[10]  ( .DIN(\IFinst/N82 ), .CLK(clk), .CLRB(n857), 
        .SETB(1'b1), .Q(\NPC[10] ), .QN(n9444) );
  dffascs1 \IFinst/PC_reg[9]  ( .DIN(\IFinst/n838 ), .CLK(clk), .CLRB(n829), 
        .SETB(1'b1), .Q(n9499) );
  dffascs1 \IFinst/NPC_reg[9]  ( .DIN(\IFinst/N81 ), .CLK(clk), .CLRB(n844), 
        .SETB(1'b1), .Q(\NPC[9] ), .QN(n9445) );
  dffascs1 \IFinst/PC_reg[8]  ( .DIN(\IFinst/n839 ), .CLK(clk), .CLRB(n829), 
        .SETB(1'b1), .Q(n9498) );
  dffascs1 \IFinst/NPC_reg[8]  ( .DIN(\IFinst/N80 ), .CLK(clk), .CLRB(n845), 
        .SETB(1'b1), .Q(\NPC[8] ), .QN(n9446) );
  dffascs1 \IFinst/PC_reg[7]  ( .DIN(\IFinst/n840 ), .CLK(clk), .CLRB(n829), 
        .SETB(1'b1), .Q(n9497) );
  dffascs1 \IFinst/NPC_reg[7]  ( .DIN(\IFinst/N79 ), .CLK(clk), .CLRB(n849), 
        .SETB(1'b1), .Q(\NPC[7] ), .QN(n9447) );
  dffascs1 \IFinst/PC_reg[6]  ( .DIN(\IFinst/n841 ), .CLK(clk), .CLRB(n829), 
        .SETB(1'b1), .Q(n9496) );
  dffascs1 \IFinst/NPC_reg[6]  ( .DIN(\IFinst/N78 ), .CLK(clk), .CLRB(n845), 
        .SETB(1'b1), .Q(\NPC[6] ), .QN(n9448) );
  dffascs1 \IFinst/PC_reg[5]  ( .DIN(\IFinst/n842 ), .CLK(clk), .CLRB(n832), 
        .SETB(1'b1), .Q(n9495) );
  dffascs1 \IFinst/NPC_reg[5]  ( .DIN(\IFinst/N77 ), .CLK(clk), .CLRB(n832), 
        .SETB(1'b1), .Q(\NPC[5] ), .QN(n9449) );
  dffascs1 \IFinst/PC_reg[4]  ( .DIN(\IFinst/n843 ), .CLK(clk), .CLRB(n832), 
        .SETB(1'b1), .Q(n9494) );
  dffascs1 \IFinst/NPC_reg[4]  ( .DIN(\IFinst/N76 ), .CLK(clk), .CLRB(n833), 
        .SETB(1'b1), .Q(\NPC[4] ), .QN(n9450) );
  dffascs1 \IFinst/PC_reg[3]  ( .DIN(\IFinst/n844 ), .CLK(clk), .CLRB(n833), 
        .SETB(1'b1), .Q(n9493) );
  dffascs1 \IFinst/NPC_reg[3]  ( .DIN(\IFinst/N75 ), .CLK(clk), .CLRB(n833), 
        .SETB(1'b1), .Q(\NPC[3] ), .QN(n9451) );
  dffascs1 \IFinst/PC_reg[2]  ( .DIN(\IFinst/n845 ), .CLK(clk), .CLRB(n830), 
        .SETB(1'b1), .Q(n9492) );
  dffascs1 \IFinst/NPC_reg[2]  ( .DIN(\IFinst/N74 ), .CLK(clk), .CLRB(n833), 
        .SETB(1'b1), .Q(\NPC[2] ), .QN(n9491) );
  dffascs1 \IFinst/PC_reg[1]  ( .DIN(\IFinst/n846 ), .CLK(clk), .CLRB(n829), 
        .SETB(1'b1), .Q(n9490) );
  dffascs1 \IFinst/NPC_reg[1]  ( .DIN(\IFinst/N73 ), .CLK(clk), .CLRB(n833), 
        .SETB(1'b1), .Q(\IFinst/N8 ), .QN(n9422) );
  dffascs1 \IFinst/NPC_reg[0]  ( .DIN(\IFinst/N72 ), .CLK(clk), .CLRB(n926), 
        .SETB(1'b1), .Q(\IFinst/N7 ), .QN(n9423) );
  dffascs1 \IFinst/stalled_reg  ( .DIN(\IFinst/n848 ), .CLK(clk), .CLRB(n958), 
        .SETB(1'b1), .QN(n9383) );
  nnd2s1 \IDinst/U11930  ( .DIN1(\IDinst/n11835 ), .DIN2(\IDinst/N48 ), 
        .Q(\IDinst/n8954 ) );
  nnd2s1 \IDinst/U11929  ( .DIN1(\IDinst/n11790 ), .DIN2(n533), 
        .Q(\IDinst/n8955 ) );
  nnd2s1 \IDinst/U11928  ( .DIN1(\IDinst/n11834 ), .DIN2(\IDinst/n11833 ), 
        .Q(\IDinst/n11835 ) );
  nnd2s1 \IDinst/U11927  ( .DIN1(\IDinst/n11832 ), .DIN2(n667), 
        .Q(\IDinst/n11834 ) );
  nnd2s1 \IDinst/U11926  ( .DIN1(\IDinst/n11811 ), .DIN2(n680), 
        .Q(\IDinst/n11833 ) );
  nnd2s1 \IDinst/U11925  ( .DIN1(\IDinst/n11831 ), .DIN2(\IDinst/n11830 ), 
        .Q(\IDinst/n11832 ) );
  nnd2s1 \IDinst/U11924  ( .DIN1(\IDinst/n11829 ), .DIN2(n1375), 
        .Q(\IDinst/n11831 ) );
  nnd2s1 \IDinst/U11923  ( .DIN1(\IDinst/n11820 ), .DIN2(n1364), 
        .Q(\IDinst/n11830 ) );
  nnd2s1 \IDinst/U11922  ( .DIN1(\IDinst/n11828 ), .DIN2(\IDinst/n11827 ), 
        .Q(\IDinst/n11829 ) );
  nnd2s1 \IDinst/U11921  ( .DIN1(\IDinst/n11826 ), .DIN2(n1322), 
        .Q(\IDinst/n11828 ) );
  nnd2s1 \IDinst/U11920  ( .DIN1(\IDinst/n11823 ), .DIN2(n1348), 
        .Q(\IDinst/n11827 ) );
  nnd2s1 \IDinst/U11919  ( .DIN1(\IDinst/n11825 ), .DIN2(\IDinst/n11824 ), 
        .Q(\IDinst/n11826 ) );
  nnd2s1 \IDinst/U11918  ( .DIN1(\IDinst/RegFile[31][31] ), .DIN2(n1218), 
        .Q(\IDinst/n11825 ) );
  nnd2s1 \IDinst/U11917  ( .DIN1(\IDinst/RegFile[30][31] ), .DIN2(n1269), 
        .Q(\IDinst/n11824 ) );
  nnd2s1 \IDinst/U11916  ( .DIN1(\IDinst/n11822 ), .DIN2(\IDinst/n11821 ), 
        .Q(\IDinst/n11823 ) );
  nnd2s1 \IDinst/U11915  ( .DIN1(\IDinst/RegFile[29][31] ), .DIN2(n1213), 
        .Q(\IDinst/n11822 ) );
  nnd2s1 \IDinst/U11914  ( .DIN1(\IDinst/RegFile[28][31] ), .DIN2(n1282), 
        .Q(\IDinst/n11821 ) );
  nnd2s1 \IDinst/U11913  ( .DIN1(\IDinst/n11819 ), .DIN2(\IDinst/n11818 ), 
        .Q(\IDinst/n11820 ) );
  nnd2s1 \IDinst/U11912  ( .DIN1(\IDinst/n11817 ), .DIN2(n1322), 
        .Q(\IDinst/n11819 ) );
  nnd2s1 \IDinst/U11911  ( .DIN1(\IDinst/n11814 ), .DIN2(n1348), 
        .Q(\IDinst/n11818 ) );
  nnd2s1 \IDinst/U11910  ( .DIN1(\IDinst/n11816 ), .DIN2(\IDinst/n11815 ), 
        .Q(\IDinst/n11817 ) );
  nnd2s1 \IDinst/U11909  ( .DIN1(\IDinst/RegFile[27][31] ), .DIN2(n1208), 
        .Q(\IDinst/n11816 ) );
  nnd2s1 \IDinst/U11908  ( .DIN1(\IDinst/RegFile[26][31] ), .DIN2(n1282), 
        .Q(\IDinst/n11815 ) );
  nnd2s1 \IDinst/U11907  ( .DIN1(\IDinst/n11813 ), .DIN2(\IDinst/n11812 ), 
        .Q(\IDinst/n11814 ) );
  nnd2s1 \IDinst/U11906  ( .DIN1(\IDinst/RegFile[25][31] ), .DIN2(n1208), 
        .Q(\IDinst/n11813 ) );
  nnd2s1 \IDinst/U11905  ( .DIN1(\IDinst/RegFile[24][31] ), .DIN2(n1282), 
        .Q(\IDinst/n11812 ) );
  nnd2s1 \IDinst/U11904  ( .DIN1(\IDinst/n11810 ), .DIN2(\IDinst/n11809 ), 
        .Q(\IDinst/n11811 ) );
  nnd2s1 \IDinst/U11903  ( .DIN1(\IDinst/n11808 ), .DIN2(n1373), 
        .Q(\IDinst/n11810 ) );
  nnd2s1 \IDinst/U11902  ( .DIN1(\IDinst/n11799 ), .DIN2(n1371), 
        .Q(\IDinst/n11809 ) );
  nnd2s1 \IDinst/U11901  ( .DIN1(\IDinst/n11807 ), .DIN2(\IDinst/n11806 ), 
        .Q(\IDinst/n11808 ) );
  nnd2s1 \IDinst/U11900  ( .DIN1(\IDinst/n11805 ), .DIN2(n1322), 
        .Q(\IDinst/n11807 ) );
  nnd2s1 \IDinst/U11899  ( .DIN1(\IDinst/n11802 ), .DIN2(n1348), 
        .Q(\IDinst/n11806 ) );
  nnd2s1 \IDinst/U11898  ( .DIN1(\IDinst/n11804 ), .DIN2(\IDinst/n11803 ), 
        .Q(\IDinst/n11805 ) );
  nnd2s1 \IDinst/U11897  ( .DIN1(\IDinst/RegFile[23][31] ), .DIN2(n1208), 
        .Q(\IDinst/n11804 ) );
  nnd2s1 \IDinst/U11896  ( .DIN1(\IDinst/RegFile[22][31] ), .DIN2(n1282), 
        .Q(\IDinst/n11803 ) );
  nnd2s1 \IDinst/U11895  ( .DIN1(\IDinst/n11801 ), .DIN2(\IDinst/n11800 ), 
        .Q(\IDinst/n11802 ) );
  nnd2s1 \IDinst/U11894  ( .DIN1(\IDinst/RegFile[21][31] ), .DIN2(n1208), 
        .Q(\IDinst/n11801 ) );
  nnd2s1 \IDinst/U11893  ( .DIN1(\IDinst/RegFile[20][31] ), .DIN2(n1282), 
        .Q(\IDinst/n11800 ) );
  nnd2s1 \IDinst/U11892  ( .DIN1(\IDinst/n11798 ), .DIN2(\IDinst/n11797 ), 
        .Q(\IDinst/n11799 ) );
  nnd2s1 \IDinst/U11891  ( .DIN1(\IDinst/n11796 ), .DIN2(n1322), 
        .Q(\IDinst/n11798 ) );
  nnd2s1 \IDinst/U11890  ( .DIN1(\IDinst/n11793 ), .DIN2(n1348), 
        .Q(\IDinst/n11797 ) );
  nnd2s1 \IDinst/U11889  ( .DIN1(\IDinst/n11795 ), .DIN2(\IDinst/n11794 ), 
        .Q(\IDinst/n11796 ) );
  nnd2s1 \IDinst/U11888  ( .DIN1(\IDinst/RegFile[19][31] ), .DIN2(n1208), 
        .Q(\IDinst/n11795 ) );
  nnd2s1 \IDinst/U11887  ( .DIN1(\IDinst/RegFile[18][31] ), .DIN2(n1282), 
        .Q(\IDinst/n11794 ) );
  nnd2s1 \IDinst/U11886  ( .DIN1(\IDinst/n11792 ), .DIN2(\IDinst/n11791 ), 
        .Q(\IDinst/n11793 ) );
  nnd2s1 \IDinst/U11885  ( .DIN1(\IDinst/RegFile[17][31] ), .DIN2(n1208), 
        .Q(\IDinst/n11792 ) );
  nnd2s1 \IDinst/U11884  ( .DIN1(\IDinst/RegFile[16][31] ), .DIN2(n1281), 
        .Q(\IDinst/n11791 ) );
  nnd2s1 \IDinst/U11883  ( .DIN1(\IDinst/n11789 ), .DIN2(\IDinst/n11788 ), 
        .Q(\IDinst/n11790 ) );
  nnd2s1 \IDinst/U11882  ( .DIN1(\IDinst/n11787 ), .DIN2(n665), 
        .Q(\IDinst/n11789 ) );
  nnd2s1 \IDinst/U11881  ( .DIN1(\IDinst/n11766 ), .DIN2(n680), 
        .Q(\IDinst/n11788 ) );
  nnd2s1 \IDinst/U11880  ( .DIN1(\IDinst/n11786 ), .DIN2(\IDinst/n11785 ), 
        .Q(\IDinst/n11787 ) );
  nnd2s1 \IDinst/U11879  ( .DIN1(\IDinst/n11784 ), .DIN2(n1373), 
        .Q(\IDinst/n11786 ) );
  nnd2s1 \IDinst/U11878  ( .DIN1(\IDinst/n11775 ), .DIN2(n1366), 
        .Q(\IDinst/n11785 ) );
  nnd2s1 \IDinst/U11877  ( .DIN1(\IDinst/n11783 ), .DIN2(\IDinst/n11782 ), 
        .Q(\IDinst/n11784 ) );
  nnd2s1 \IDinst/U11876  ( .DIN1(\IDinst/n11781 ), .DIN2(n1322), 
        .Q(\IDinst/n11783 ) );
  nnd2s1 \IDinst/U11875  ( .DIN1(\IDinst/n11778 ), .DIN2(n1348), 
        .Q(\IDinst/n11782 ) );
  nnd2s1 \IDinst/U11874  ( .DIN1(\IDinst/n11780 ), .DIN2(\IDinst/n11779 ), 
        .Q(\IDinst/n11781 ) );
  nnd2s1 \IDinst/U11873  ( .DIN1(\IDinst/RegFile[15][31] ), .DIN2(n1209), 
        .Q(\IDinst/n11780 ) );
  nnd2s1 \IDinst/U11872  ( .DIN1(\IDinst/RegFile[14][31] ), .DIN2(n1281), 
        .Q(\IDinst/n11779 ) );
  nnd2s1 \IDinst/U11871  ( .DIN1(\IDinst/n11777 ), .DIN2(\IDinst/n11776 ), 
        .Q(\IDinst/n11778 ) );
  nnd2s1 \IDinst/U11870  ( .DIN1(\IDinst/RegFile[13][31] ), .DIN2(n1209), 
        .Q(\IDinst/n11777 ) );
  nnd2s1 \IDinst/U11869  ( .DIN1(\IDinst/RegFile[12][31] ), .DIN2(n1281), 
        .Q(\IDinst/n11776 ) );
  nnd2s1 \IDinst/U11868  ( .DIN1(\IDinst/n11774 ), .DIN2(\IDinst/n11773 ), 
        .Q(\IDinst/n11775 ) );
  nnd2s1 \IDinst/U11867  ( .DIN1(\IDinst/n11772 ), .DIN2(n1322), 
        .Q(\IDinst/n11774 ) );
  nnd2s1 \IDinst/U11866  ( .DIN1(\IDinst/n11769 ), .DIN2(n1348), 
        .Q(\IDinst/n11773 ) );
  nnd2s1 \IDinst/U11865  ( .DIN1(\IDinst/n11771 ), .DIN2(\IDinst/n11770 ), 
        .Q(\IDinst/n11772 ) );
  nnd2s1 \IDinst/U11864  ( .DIN1(\IDinst/RegFile[11][31] ), .DIN2(n1209), 
        .Q(\IDinst/n11771 ) );
  nnd2s1 \IDinst/U11863  ( .DIN1(\IDinst/RegFile[10][31] ), .DIN2(n1281), 
        .Q(\IDinst/n11770 ) );
  nnd2s1 \IDinst/U11862  ( .DIN1(\IDinst/n11768 ), .DIN2(\IDinst/n11767 ), 
        .Q(\IDinst/n11769 ) );
  nnd2s1 \IDinst/U11861  ( .DIN1(\IDinst/RegFile[9][31] ), .DIN2(n1209), 
        .Q(\IDinst/n11768 ) );
  nnd2s1 \IDinst/U11860  ( .DIN1(\IDinst/RegFile[8][31] ), .DIN2(n1281), 
        .Q(\IDinst/n11767 ) );
  nnd2s1 \IDinst/U11859  ( .DIN1(\IDinst/n11765 ), .DIN2(\IDinst/n11764 ), 
        .Q(\IDinst/n11766 ) );
  nnd2s1 \IDinst/U11858  ( .DIN1(\IDinst/n11763 ), .DIN2(n1373), 
        .Q(\IDinst/n11765 ) );
  nnd2s1 \IDinst/U11857  ( .DIN1(\IDinst/n11754 ), .DIN2(n1370), 
        .Q(\IDinst/n11764 ) );
  nnd2s1 \IDinst/U11856  ( .DIN1(\IDinst/n11762 ), .DIN2(\IDinst/n11761 ), 
        .Q(\IDinst/n11763 ) );
  nnd2s1 \IDinst/U11855  ( .DIN1(\IDinst/n11760 ), .DIN2(n1322), 
        .Q(\IDinst/n11762 ) );
  nnd2s1 \IDinst/U11854  ( .DIN1(\IDinst/n11757 ), .DIN2(n1349), 
        .Q(\IDinst/n11761 ) );
  nnd2s1 \IDinst/U11853  ( .DIN1(\IDinst/n11759 ), .DIN2(\IDinst/n11758 ), 
        .Q(\IDinst/n11760 ) );
  nnd2s1 \IDinst/U11852  ( .DIN1(\IDinst/RegFile[7][31] ), .DIN2(n1209), 
        .Q(\IDinst/n11759 ) );
  nnd2s1 \IDinst/U11851  ( .DIN1(\IDinst/RegFile[6][31] ), .DIN2(n1281), 
        .Q(\IDinst/n11758 ) );
  nnd2s1 \IDinst/U11850  ( .DIN1(\IDinst/n11756 ), .DIN2(\IDinst/n11755 ), 
        .Q(\IDinst/n11757 ) );
  nnd2s1 \IDinst/U11849  ( .DIN1(\IDinst/RegFile[5][31] ), .DIN2(n1209), 
        .Q(\IDinst/n11756 ) );
  nnd2s1 \IDinst/U11848  ( .DIN1(\IDinst/RegFile[4][31] ), .DIN2(n1281), 
        .Q(\IDinst/n11755 ) );
  nnd2s1 \IDinst/U11847  ( .DIN1(\IDinst/n11753 ), .DIN2(\IDinst/n11752 ), 
        .Q(\IDinst/n11754 ) );
  nnd2s1 \IDinst/U11846  ( .DIN1(\IDinst/n11751 ), .DIN2(n1321), 
        .Q(\IDinst/n11753 ) );
  nnd2s1 \IDinst/U11845  ( .DIN1(\IDinst/n11748 ), .DIN2(n1349), 
        .Q(\IDinst/n11752 ) );
  nnd2s1 \IDinst/U11844  ( .DIN1(\IDinst/n11750 ), .DIN2(\IDinst/n11749 ), 
        .Q(\IDinst/n11751 ) );
  nnd2s1 \IDinst/U11843  ( .DIN1(\IDinst/RegFile[3][31] ), .DIN2(n1209), 
        .Q(\IDinst/n11750 ) );
  nnd2s1 \IDinst/U11842  ( .DIN1(\IDinst/RegFile[2][31] ), .DIN2(n1281), 
        .Q(\IDinst/n11749 ) );
  nnd2s1 \IDinst/U11841  ( .DIN1(\IDinst/n11747 ), .DIN2(\IDinst/n11746 ), 
        .Q(\IDinst/n11748 ) );
  nnd2s1 \IDinst/U11840  ( .DIN1(\IDinst/RegFile[1][31] ), .DIN2(n1209), 
        .Q(\IDinst/n11747 ) );
  nnd2s1 \IDinst/U11839  ( .DIN1(\IDinst/RegFile[0][31] ), .DIN2(n1281), 
        .Q(\IDinst/n11746 ) );
  nnd2s1 \IDinst/U11838  ( .DIN1(\IDinst/n11745 ), .DIN2(n535), 
        .Q(\IDinst/n8952 ) );
  nnd2s1 \IDinst/U11837  ( .DIN1(\IDinst/n11700 ), .DIN2(n634), 
        .Q(\IDinst/n8953 ) );
  nnd2s1 \IDinst/U11836  ( .DIN1(\IDinst/n11744 ), .DIN2(\IDinst/n11743 ), 
        .Q(\IDinst/n11745 ) );
  nnd2s1 \IDinst/U11835  ( .DIN1(\IDinst/n11742 ), .DIN2(n668), 
        .Q(\IDinst/n11744 ) );
  nnd2s1 \IDinst/U11834  ( .DIN1(\IDinst/n11721 ), .DIN2(n683), 
        .Q(\IDinst/n11743 ) );
  nnd2s1 \IDinst/U11833  ( .DIN1(\IDinst/n11741 ), .DIN2(\IDinst/n11740 ), 
        .Q(\IDinst/n11742 ) );
  nnd2s1 \IDinst/U11832  ( .DIN1(\IDinst/n11739 ), .DIN2(n1373), 
        .Q(\IDinst/n11741 ) );
  nnd2s1 \IDinst/U11831  ( .DIN1(\IDinst/n11730 ), .DIN2(n1365), 
        .Q(\IDinst/n11740 ) );
  nnd2s1 \IDinst/U11830  ( .DIN1(\IDinst/n11738 ), .DIN2(\IDinst/n11737 ), 
        .Q(\IDinst/n11739 ) );
  nnd2s1 \IDinst/U11829  ( .DIN1(\IDinst/n11736 ), .DIN2(n1321), 
        .Q(\IDinst/n11738 ) );
  nnd2s1 \IDinst/U11828  ( .DIN1(\IDinst/n11733 ), .DIN2(n1349), 
        .Q(\IDinst/n11737 ) );
  nnd2s1 \IDinst/U11827  ( .DIN1(\IDinst/n11735 ), .DIN2(\IDinst/n11734 ), 
        .Q(\IDinst/n11736 ) );
  nnd2s1 \IDinst/U11826  ( .DIN1(\IDinst/RegFile[31][30] ), .DIN2(n1209), 
        .Q(\IDinst/n11735 ) );
  nnd2s1 \IDinst/U11825  ( .DIN1(\IDinst/RegFile[30][30] ), .DIN2(n1280), 
        .Q(\IDinst/n11734 ) );
  nnd2s1 \IDinst/U11824  ( .DIN1(\IDinst/n11732 ), .DIN2(\IDinst/n11731 ), 
        .Q(\IDinst/n11733 ) );
  nnd2s1 \IDinst/U11823  ( .DIN1(\IDinst/RegFile[29][30] ), .DIN2(n1209), 
        .Q(\IDinst/n11732 ) );
  nnd2s1 \IDinst/U11822  ( .DIN1(\IDinst/RegFile[28][30] ), .DIN2(n1280), 
        .Q(\IDinst/n11731 ) );
  nnd2s1 \IDinst/U11821  ( .DIN1(\IDinst/n11729 ), .DIN2(\IDinst/n11728 ), 
        .Q(\IDinst/n11730 ) );
  nnd2s1 \IDinst/U11820  ( .DIN1(\IDinst/n11727 ), .DIN2(n1321), 
        .Q(\IDinst/n11729 ) );
  nnd2s1 \IDinst/U11819  ( .DIN1(\IDinst/n11724 ), .DIN2(n1349), 
        .Q(\IDinst/n11728 ) );
  nnd2s1 \IDinst/U11818  ( .DIN1(\IDinst/n11726 ), .DIN2(\IDinst/n11725 ), 
        .Q(\IDinst/n11727 ) );
  nnd2s1 \IDinst/U11817  ( .DIN1(\IDinst/RegFile[27][30] ), .DIN2(n1209), 
        .Q(\IDinst/n11726 ) );
  nnd2s1 \IDinst/U11816  ( .DIN1(\IDinst/RegFile[26][30] ), .DIN2(n1280), 
        .Q(\IDinst/n11725 ) );
  nnd2s1 \IDinst/U11815  ( .DIN1(\IDinst/n11723 ), .DIN2(\IDinst/n11722 ), 
        .Q(\IDinst/n11724 ) );
  nnd2s1 \IDinst/U11814  ( .DIN1(\IDinst/RegFile[25][30] ), .DIN2(n1209), 
        .Q(\IDinst/n11723 ) );
  nnd2s1 \IDinst/U11813  ( .DIN1(\IDinst/RegFile[24][30] ), .DIN2(n1280), 
        .Q(\IDinst/n11722 ) );
  nnd2s1 \IDinst/U11812  ( .DIN1(\IDinst/n11720 ), .DIN2(\IDinst/n11719 ), 
        .Q(\IDinst/n11721 ) );
  nnd2s1 \IDinst/U11811  ( .DIN1(\IDinst/n11718 ), .DIN2(n1373), 
        .Q(\IDinst/n11720 ) );
  nnd2s1 \IDinst/U11810  ( .DIN1(\IDinst/n11709 ), .DIN2(n1369), 
        .Q(\IDinst/n11719 ) );
  nnd2s1 \IDinst/U11809  ( .DIN1(\IDinst/n11717 ), .DIN2(\IDinst/n11716 ), 
        .Q(\IDinst/n11718 ) );
  nnd2s1 \IDinst/U11808  ( .DIN1(\IDinst/n11715 ), .DIN2(n1321), 
        .Q(\IDinst/n11717 ) );
  nnd2s1 \IDinst/U11807  ( .DIN1(\IDinst/n11712 ), .DIN2(n1349), 
        .Q(\IDinst/n11716 ) );
  nnd2s1 \IDinst/U11806  ( .DIN1(\IDinst/n11714 ), .DIN2(\IDinst/n11713 ), 
        .Q(\IDinst/n11715 ) );
  nnd2s1 \IDinst/U11805  ( .DIN1(\IDinst/RegFile[23][30] ), .DIN2(n1209), 
        .Q(\IDinst/n11714 ) );
  nnd2s1 \IDinst/U11804  ( .DIN1(\IDinst/RegFile[22][30] ), .DIN2(n1280), 
        .Q(\IDinst/n11713 ) );
  nnd2s1 \IDinst/U11803  ( .DIN1(\IDinst/n11711 ), .DIN2(\IDinst/n11710 ), 
        .Q(\IDinst/n11712 ) );
  nnd2s1 \IDinst/U11802  ( .DIN1(\IDinst/RegFile[21][30] ), .DIN2(n1210), 
        .Q(\IDinst/n11711 ) );
  nnd2s1 \IDinst/U11801  ( .DIN1(\IDinst/RegFile[20][30] ), .DIN2(n1280), 
        .Q(\IDinst/n11710 ) );
  nnd2s1 \IDinst/U11800  ( .DIN1(\IDinst/n11708 ), .DIN2(\IDinst/n11707 ), 
        .Q(\IDinst/n11709 ) );
  nnd2s1 \IDinst/U11799  ( .DIN1(\IDinst/n11706 ), .DIN2(n1321), 
        .Q(\IDinst/n11708 ) );
  nnd2s1 \IDinst/U11798  ( .DIN1(\IDinst/n11703 ), .DIN2(n1349), 
        .Q(\IDinst/n11707 ) );
  nnd2s1 \IDinst/U11797  ( .DIN1(\IDinst/n11705 ), .DIN2(\IDinst/n11704 ), 
        .Q(\IDinst/n11706 ) );
  nnd2s1 \IDinst/U11796  ( .DIN1(\IDinst/RegFile[19][30] ), .DIN2(n1210), 
        .Q(\IDinst/n11705 ) );
  nnd2s1 \IDinst/U11795  ( .DIN1(\IDinst/RegFile[18][30] ), .DIN2(n1280), 
        .Q(\IDinst/n11704 ) );
  nnd2s1 \IDinst/U11794  ( .DIN1(\IDinst/n11702 ), .DIN2(\IDinst/n11701 ), 
        .Q(\IDinst/n11703 ) );
  nnd2s1 \IDinst/U11793  ( .DIN1(\IDinst/RegFile[17][30] ), .DIN2(n1210), 
        .Q(\IDinst/n11702 ) );
  nnd2s1 \IDinst/U11792  ( .DIN1(\IDinst/RegFile[16][30] ), .DIN2(n1280), 
        .Q(\IDinst/n11701 ) );
  nnd2s1 \IDinst/U11791  ( .DIN1(\IDinst/n11699 ), .DIN2(\IDinst/n11698 ), 
        .Q(\IDinst/n11700 ) );
  nnd2s1 \IDinst/U11790  ( .DIN1(\IDinst/n11697 ), .DIN2(n666), 
        .Q(\IDinst/n11699 ) );
  nnd2s1 \IDinst/U11789  ( .DIN1(\IDinst/n11676 ), .DIN2(n682), 
        .Q(\IDinst/n11698 ) );
  nnd2s1 \IDinst/U11788  ( .DIN1(\IDinst/n11696 ), .DIN2(\IDinst/n11695 ), 
        .Q(\IDinst/n11697 ) );
  nnd2s1 \IDinst/U11787  ( .DIN1(\IDinst/n11694 ), .DIN2(n1373), 
        .Q(\IDinst/n11696 ) );
  nnd2s1 \IDinst/U11786  ( .DIN1(\IDinst/n11685 ), .DIN2(n1365), 
        .Q(\IDinst/n11695 ) );
  nnd2s1 \IDinst/U11785  ( .DIN1(\IDinst/n11693 ), .DIN2(\IDinst/n11692 ), 
        .Q(\IDinst/n11694 ) );
  nnd2s1 \IDinst/U11784  ( .DIN1(\IDinst/n11691 ), .DIN2(n1321), 
        .Q(\IDinst/n11693 ) );
  nnd2s1 \IDinst/U11783  ( .DIN1(\IDinst/n11688 ), .DIN2(n1349), 
        .Q(\IDinst/n11692 ) );
  nnd2s1 \IDinst/U11782  ( .DIN1(\IDinst/n11690 ), .DIN2(\IDinst/n11689 ), 
        .Q(\IDinst/n11691 ) );
  nnd2s1 \IDinst/U11781  ( .DIN1(\IDinst/RegFile[15][30] ), .DIN2(n1210), 
        .Q(\IDinst/n11690 ) );
  nnd2s1 \IDinst/U11780  ( .DIN1(\IDinst/RegFile[14][30] ), .DIN2(n1280), 
        .Q(\IDinst/n11689 ) );
  nnd2s1 \IDinst/U11779  ( .DIN1(\IDinst/n11687 ), .DIN2(\IDinst/n11686 ), 
        .Q(\IDinst/n11688 ) );
  nnd2s1 \IDinst/U11778  ( .DIN1(\IDinst/RegFile[13][30] ), .DIN2(n1210), 
        .Q(\IDinst/n11687 ) );
  nnd2s1 \IDinst/U11777  ( .DIN1(\IDinst/RegFile[12][30] ), .DIN2(n1279), 
        .Q(\IDinst/n11686 ) );
  nnd2s1 \IDinst/U11776  ( .DIN1(\IDinst/n11684 ), .DIN2(\IDinst/n11683 ), 
        .Q(\IDinst/n11685 ) );
  nnd2s1 \IDinst/U11775  ( .DIN1(\IDinst/n11682 ), .DIN2(n1321), 
        .Q(\IDinst/n11684 ) );
  nnd2s1 \IDinst/U11774  ( .DIN1(\IDinst/n11679 ), .DIN2(n1349), 
        .Q(\IDinst/n11683 ) );
  nnd2s1 \IDinst/U11773  ( .DIN1(\IDinst/n11681 ), .DIN2(\IDinst/n11680 ), 
        .Q(\IDinst/n11682 ) );
  nnd2s1 \IDinst/U11772  ( .DIN1(\IDinst/RegFile[11][30] ), .DIN2(n1210), 
        .Q(\IDinst/n11681 ) );
  nnd2s1 \IDinst/U11771  ( .DIN1(\IDinst/RegFile[10][30] ), .DIN2(n1279), 
        .Q(\IDinst/n11680 ) );
  nnd2s1 \IDinst/U11770  ( .DIN1(\IDinst/n11678 ), .DIN2(\IDinst/n11677 ), 
        .Q(\IDinst/n11679 ) );
  nnd2s1 \IDinst/U11769  ( .DIN1(\IDinst/RegFile[9][30] ), .DIN2(n1210), 
        .Q(\IDinst/n11678 ) );
  nnd2s1 \IDinst/U11768  ( .DIN1(\IDinst/RegFile[8][30] ), .DIN2(n1279), 
        .Q(\IDinst/n11677 ) );
  nnd2s1 \IDinst/U11767  ( .DIN1(\IDinst/n11675 ), .DIN2(\IDinst/n11674 ), 
        .Q(\IDinst/n11676 ) );
  nnd2s1 \IDinst/U11766  ( .DIN1(\IDinst/n11673 ), .DIN2(n1376), 
        .Q(\IDinst/n11675 ) );
  nnd2s1 \IDinst/U11765  ( .DIN1(\IDinst/n11664 ), .DIN2(n1368), 
        .Q(\IDinst/n11674 ) );
  nnd2s1 \IDinst/U11764  ( .DIN1(\IDinst/n11672 ), .DIN2(\IDinst/n11671 ), 
        .Q(\IDinst/n11673 ) );
  nnd2s1 \IDinst/U11763  ( .DIN1(\IDinst/n11670 ), .DIN2(n1321), 
        .Q(\IDinst/n11672 ) );
  nnd2s1 \IDinst/U11762  ( .DIN1(\IDinst/n11667 ), .DIN2(n1349), 
        .Q(\IDinst/n11671 ) );
  nnd2s1 \IDinst/U11761  ( .DIN1(\IDinst/n11669 ), .DIN2(\IDinst/n11668 ), 
        .Q(\IDinst/n11670 ) );
  nnd2s1 \IDinst/U11760  ( .DIN1(\IDinst/RegFile[7][30] ), .DIN2(n1210), 
        .Q(\IDinst/n11669 ) );
  nnd2s1 \IDinst/U11759  ( .DIN1(\IDinst/RegFile[6][30] ), .DIN2(n1279), 
        .Q(\IDinst/n11668 ) );
  nnd2s1 \IDinst/U11758  ( .DIN1(\IDinst/n11666 ), .DIN2(\IDinst/n11665 ), 
        .Q(\IDinst/n11667 ) );
  nnd2s1 \IDinst/U11757  ( .DIN1(\IDinst/RegFile[5][30] ), .DIN2(n1210), 
        .Q(\IDinst/n11666 ) );
  nnd2s1 \IDinst/U11756  ( .DIN1(\IDinst/RegFile[4][30] ), .DIN2(n1279), 
        .Q(\IDinst/n11665 ) );
  nnd2s1 \IDinst/U11755  ( .DIN1(\IDinst/n11663 ), .DIN2(\IDinst/n11662 ), 
        .Q(\IDinst/n11664 ) );
  nnd2s1 \IDinst/U11754  ( .DIN1(\IDinst/n11661 ), .DIN2(n1321), 
        .Q(\IDinst/n11663 ) );
  nnd2s1 \IDinst/U11753  ( .DIN1(\IDinst/n11658 ), .DIN2(n1350), 
        .Q(\IDinst/n11662 ) );
  nnd2s1 \IDinst/U11752  ( .DIN1(\IDinst/n11660 ), .DIN2(\IDinst/n11659 ), 
        .Q(\IDinst/n11661 ) );
  nnd2s1 \IDinst/U11751  ( .DIN1(\IDinst/RegFile[3][30] ), .DIN2(n1210), 
        .Q(\IDinst/n11660 ) );
  nnd2s1 \IDinst/U11750  ( .DIN1(\IDinst/RegFile[2][30] ), .DIN2(n1279), 
        .Q(\IDinst/n11659 ) );
  nnd2s1 \IDinst/U11749  ( .DIN1(\IDinst/n11657 ), .DIN2(\IDinst/n11656 ), 
        .Q(\IDinst/n11658 ) );
  nnd2s1 \IDinst/U11748  ( .DIN1(\IDinst/RegFile[1][30] ), .DIN2(n1210), 
        .Q(\IDinst/n11657 ) );
  nnd2s1 \IDinst/U11747  ( .DIN1(\IDinst/RegFile[0][30] ), .DIN2(n1279), 
        .Q(\IDinst/n11656 ) );
  nnd2s1 \IDinst/U11746  ( .DIN1(\IDinst/n11655 ), .DIN2(n534), 
        .Q(\IDinst/n8950 ) );
  nnd2s1 \IDinst/U11745  ( .DIN1(\IDinst/n11610 ), .DIN2(n533), 
        .Q(\IDinst/n8951 ) );
  nnd2s1 \IDinst/U11744  ( .DIN1(\IDinst/n11654 ), .DIN2(\IDinst/n11653 ), 
        .Q(\IDinst/n11655 ) );
  nnd2s1 \IDinst/U11743  ( .DIN1(\IDinst/n11652 ), .DIN2(n667), 
        .Q(\IDinst/n11654 ) );
  nnd2s1 \IDinst/U11742  ( .DIN1(\IDinst/n11631 ), .DIN2(n680), 
        .Q(\IDinst/n11653 ) );
  nnd2s1 \IDinst/U11741  ( .DIN1(\IDinst/n11651 ), .DIN2(\IDinst/n11650 ), 
        .Q(\IDinst/n11652 ) );
  nnd2s1 \IDinst/U11740  ( .DIN1(\IDinst/n11649 ), .DIN2(n1373), 
        .Q(\IDinst/n11651 ) );
  nnd2s1 \IDinst/U11739  ( .DIN1(\IDinst/n11640 ), .DIN2(n1371), 
        .Q(\IDinst/n11650 ) );
  nnd2s1 \IDinst/U11738  ( .DIN1(\IDinst/n11648 ), .DIN2(\IDinst/n11647 ), 
        .Q(\IDinst/n11649 ) );
  nnd2s1 \IDinst/U11737  ( .DIN1(\IDinst/n11646 ), .DIN2(n1321), 
        .Q(\IDinst/n11648 ) );
  nnd2s1 \IDinst/U11736  ( .DIN1(\IDinst/n11643 ), .DIN2(n1350), 
        .Q(\IDinst/n11647 ) );
  nnd2s1 \IDinst/U11735  ( .DIN1(\IDinst/n11645 ), .DIN2(\IDinst/n11644 ), 
        .Q(\IDinst/n11646 ) );
  nnd2s1 \IDinst/U11734  ( .DIN1(\IDinst/RegFile[31][29] ), .DIN2(n1210), 
        .Q(\IDinst/n11645 ) );
  nnd2s1 \IDinst/U11733  ( .DIN1(\IDinst/RegFile[30][29] ), .DIN2(n1279), 
        .Q(\IDinst/n11644 ) );
  nnd2s1 \IDinst/U11732  ( .DIN1(\IDinst/n11642 ), .DIN2(\IDinst/n11641 ), 
        .Q(\IDinst/n11643 ) );
  nnd2s1 \IDinst/U11731  ( .DIN1(\IDinst/RegFile[29][29] ), .DIN2(n1210), 
        .Q(\IDinst/n11642 ) );
  nnd2s1 \IDinst/U11730  ( .DIN1(\IDinst/RegFile[28][29] ), .DIN2(n1279), 
        .Q(\IDinst/n11641 ) );
  nnd2s1 \IDinst/U11729  ( .DIN1(\IDinst/n11639 ), .DIN2(\IDinst/n11638 ), 
        .Q(\IDinst/n11640 ) );
  nnd2s1 \IDinst/U11728  ( .DIN1(\IDinst/n11637 ), .DIN2(n1321), 
        .Q(\IDinst/n11639 ) );
  nnd2s1 \IDinst/U11727  ( .DIN1(\IDinst/n11634 ), .DIN2(n1350), 
        .Q(\IDinst/n11638 ) );
  nnd2s1 \IDinst/U11726  ( .DIN1(\IDinst/n11636 ), .DIN2(\IDinst/n11635 ), 
        .Q(\IDinst/n11637 ) );
  nnd2s1 \IDinst/U11725  ( .DIN1(\IDinst/RegFile[27][29] ), .DIN2(n1211), 
        .Q(\IDinst/n11636 ) );
  nnd2s1 \IDinst/U11724  ( .DIN1(\IDinst/RegFile[26][29] ), .DIN2(n1278), 
        .Q(\IDinst/n11635 ) );
  nnd2s1 \IDinst/U11723  ( .DIN1(\IDinst/n11633 ), .DIN2(\IDinst/n11632 ), 
        .Q(\IDinst/n11634 ) );
  nnd2s1 \IDinst/U11722  ( .DIN1(\IDinst/RegFile[25][29] ), .DIN2(n1211), 
        .Q(\IDinst/n11633 ) );
  nnd2s1 \IDinst/U11721  ( .DIN1(\IDinst/RegFile[24][29] ), .DIN2(n1278), 
        .Q(\IDinst/n11632 ) );
  nnd2s1 \IDinst/U11720  ( .DIN1(\IDinst/n11630 ), .DIN2(\IDinst/n11629 ), 
        .Q(\IDinst/n11631 ) );
  nnd2s1 \IDinst/U11719  ( .DIN1(\IDinst/n11628 ), .DIN2(n1373), 
        .Q(\IDinst/n11630 ) );
  nnd2s1 \IDinst/U11718  ( .DIN1(\IDinst/n11619 ), .DIN2(n1370), 
        .Q(\IDinst/n11629 ) );
  nnd2s1 \IDinst/U11717  ( .DIN1(\IDinst/n11627 ), .DIN2(\IDinst/n11626 ), 
        .Q(\IDinst/n11628 ) );
  nnd2s1 \IDinst/U11716  ( .DIN1(\IDinst/n11625 ), .DIN2(n1321), 
        .Q(\IDinst/n11627 ) );
  nnd2s1 \IDinst/U11715  ( .DIN1(\IDinst/n11622 ), .DIN2(n1350), 
        .Q(\IDinst/n11626 ) );
  nnd2s1 \IDinst/U11714  ( .DIN1(\IDinst/n11624 ), .DIN2(\IDinst/n11623 ), 
        .Q(\IDinst/n11625 ) );
  nnd2s1 \IDinst/U11713  ( .DIN1(\IDinst/RegFile[23][29] ), .DIN2(n1211), 
        .Q(\IDinst/n11624 ) );
  nnd2s1 \IDinst/U11712  ( .DIN1(\IDinst/RegFile[22][29] ), .DIN2(n1278), 
        .Q(\IDinst/n11623 ) );
  nnd2s1 \IDinst/U11711  ( .DIN1(\IDinst/n11621 ), .DIN2(\IDinst/n11620 ), 
        .Q(\IDinst/n11622 ) );
  nnd2s1 \IDinst/U11710  ( .DIN1(\IDinst/RegFile[21][29] ), .DIN2(n1211), 
        .Q(\IDinst/n11621 ) );
  nnd2s1 \IDinst/U11709  ( .DIN1(\IDinst/RegFile[20][29] ), .DIN2(n1278), 
        .Q(\IDinst/n11620 ) );
  nnd2s1 \IDinst/U11708  ( .DIN1(\IDinst/n11618 ), .DIN2(\IDinst/n11617 ), 
        .Q(\IDinst/n11619 ) );
  nnd2s1 \IDinst/U11707  ( .DIN1(\IDinst/n11616 ), .DIN2(n1321), 
        .Q(\IDinst/n11618 ) );
  nnd2s1 \IDinst/U11706  ( .DIN1(\IDinst/n11613 ), .DIN2(n1350), 
        .Q(\IDinst/n11617 ) );
  nnd2s1 \IDinst/U11705  ( .DIN1(\IDinst/n11615 ), .DIN2(\IDinst/n11614 ), 
        .Q(\IDinst/n11616 ) );
  nnd2s1 \IDinst/U11704  ( .DIN1(\IDinst/RegFile[19][29] ), .DIN2(n1211), 
        .Q(\IDinst/n11615 ) );
  nnd2s1 \IDinst/U11703  ( .DIN1(\IDinst/RegFile[18][29] ), .DIN2(n1278), 
        .Q(\IDinst/n11614 ) );
  nnd2s1 \IDinst/U11702  ( .DIN1(\IDinst/n11612 ), .DIN2(\IDinst/n11611 ), 
        .Q(\IDinst/n11613 ) );
  nnd2s1 \IDinst/U11701  ( .DIN1(\IDinst/RegFile[17][29] ), .DIN2(n1211), 
        .Q(\IDinst/n11612 ) );
  nnd2s1 \IDinst/U11700  ( .DIN1(\IDinst/RegFile[16][29] ), .DIN2(n1278), 
        .Q(\IDinst/n11611 ) );
  nnd2s1 \IDinst/U11699  ( .DIN1(\IDinst/n11609 ), .DIN2(\IDinst/n11608 ), 
        .Q(\IDinst/n11610 ) );
  nnd2s1 \IDinst/U11698  ( .DIN1(\IDinst/n11607 ), .DIN2(n665), 
        .Q(\IDinst/n11609 ) );
  nnd2s1 \IDinst/U11697  ( .DIN1(\IDinst/n11586 ), .DIN2(n683), 
        .Q(\IDinst/n11608 ) );
  nnd2s1 \IDinst/U11696  ( .DIN1(\IDinst/n11606 ), .DIN2(\IDinst/n11605 ), 
        .Q(\IDinst/n11607 ) );
  nnd2s1 \IDinst/U11695  ( .DIN1(\IDinst/n11604 ), .DIN2(n1373), 
        .Q(\IDinst/n11606 ) );
  nnd2s1 \IDinst/U11694  ( .DIN1(\IDinst/n11595 ), .DIN2(n1369), 
        .Q(\IDinst/n11605 ) );
  nnd2s1 \IDinst/U11693  ( .DIN1(\IDinst/n11603 ), .DIN2(\IDinst/n11602 ), 
        .Q(\IDinst/n11604 ) );
  nnd2s1 \IDinst/U11692  ( .DIN1(\IDinst/n11601 ), .DIN2(n1320), 
        .Q(\IDinst/n11603 ) );
  nnd2s1 \IDinst/U11691  ( .DIN1(\IDinst/n11598 ), .DIN2(n1350), 
        .Q(\IDinst/n11602 ) );
  nnd2s1 \IDinst/U11690  ( .DIN1(\IDinst/n11600 ), .DIN2(\IDinst/n11599 ), 
        .Q(\IDinst/n11601 ) );
  nnd2s1 \IDinst/U11689  ( .DIN1(\IDinst/RegFile[15][29] ), .DIN2(n1211), 
        .Q(\IDinst/n11600 ) );
  nnd2s1 \IDinst/U11688  ( .DIN1(\IDinst/RegFile[14][29] ), .DIN2(n1278), 
        .Q(\IDinst/n11599 ) );
  nnd2s1 \IDinst/U11687  ( .DIN1(\IDinst/n11597 ), .DIN2(\IDinst/n11596 ), 
        .Q(\IDinst/n11598 ) );
  nnd2s1 \IDinst/U11686  ( .DIN1(\IDinst/RegFile[13][29] ), .DIN2(n1211), 
        .Q(\IDinst/n11597 ) );
  nnd2s1 \IDinst/U11685  ( .DIN1(\IDinst/RegFile[12][29] ), .DIN2(n1278), 
        .Q(\IDinst/n11596 ) );
  nnd2s1 \IDinst/U11684  ( .DIN1(\IDinst/n11594 ), .DIN2(\IDinst/n11593 ), 
        .Q(\IDinst/n11595 ) );
  nnd2s1 \IDinst/U11683  ( .DIN1(\IDinst/n11592 ), .DIN2(n1320), 
        .Q(\IDinst/n11594 ) );
  nnd2s1 \IDinst/U11682  ( .DIN1(\IDinst/n11589 ), .DIN2(n1350), 
        .Q(\IDinst/n11593 ) );
  nnd2s1 \IDinst/U11681  ( .DIN1(\IDinst/n11591 ), .DIN2(\IDinst/n11590 ), 
        .Q(\IDinst/n11592 ) );
  nnd2s1 \IDinst/U11680  ( .DIN1(\IDinst/RegFile[11][29] ), .DIN2(n1211), 
        .Q(\IDinst/n11591 ) );
  nnd2s1 \IDinst/U11679  ( .DIN1(\IDinst/RegFile[10][29] ), .DIN2(n1278), 
        .Q(\IDinst/n11590 ) );
  nnd2s1 \IDinst/U11678  ( .DIN1(\IDinst/n11588 ), .DIN2(\IDinst/n11587 ), 
        .Q(\IDinst/n11589 ) );
  nnd2s1 \IDinst/U11677  ( .DIN1(\IDinst/RegFile[9][29] ), .DIN2(n1211), 
        .Q(\IDinst/n11588 ) );
  nnd2s1 \IDinst/U11676  ( .DIN1(\IDinst/RegFile[8][29] ), .DIN2(n1277), 
        .Q(\IDinst/n11587 ) );
  nnd2s1 \IDinst/U11675  ( .DIN1(\IDinst/n11585 ), .DIN2(\IDinst/n11584 ), 
        .Q(\IDinst/n11586 ) );
  nnd2s1 \IDinst/U11674  ( .DIN1(\IDinst/n11583 ), .DIN2(n1373), 
        .Q(\IDinst/n11585 ) );
  nnd2s1 \IDinst/U11673  ( .DIN1(\IDinst/n11574 ), .DIN2(n1368), 
        .Q(\IDinst/n11584 ) );
  nnd2s1 \IDinst/U11672  ( .DIN1(\IDinst/n11582 ), .DIN2(\IDinst/n11581 ), 
        .Q(\IDinst/n11583 ) );
  nnd2s1 \IDinst/U11671  ( .DIN1(\IDinst/n11580 ), .DIN2(n1320), 
        .Q(\IDinst/n11582 ) );
  nnd2s1 \IDinst/U11670  ( .DIN1(\IDinst/n11577 ), .DIN2(n1350), 
        .Q(\IDinst/n11581 ) );
  nnd2s1 \IDinst/U11669  ( .DIN1(\IDinst/n11579 ), .DIN2(\IDinst/n11578 ), 
        .Q(\IDinst/n11580 ) );
  nnd2s1 \IDinst/U11668  ( .DIN1(\IDinst/RegFile[7][29] ), .DIN2(n1211), 
        .Q(\IDinst/n11579 ) );
  nnd2s1 \IDinst/U11667  ( .DIN1(\IDinst/RegFile[6][29] ), .DIN2(n1277), 
        .Q(\IDinst/n11578 ) );
  nnd2s1 \IDinst/U11666  ( .DIN1(\IDinst/n11576 ), .DIN2(\IDinst/n11575 ), 
        .Q(\IDinst/n11577 ) );
  nnd2s1 \IDinst/U11665  ( .DIN1(\IDinst/RegFile[5][29] ), .DIN2(n1211), 
        .Q(\IDinst/n11576 ) );
  nnd2s1 \IDinst/U11664  ( .DIN1(\IDinst/RegFile[4][29] ), .DIN2(n1277), 
        .Q(\IDinst/n11575 ) );
  nnd2s1 \IDinst/U11663  ( .DIN1(\IDinst/n11573 ), .DIN2(\IDinst/n11572 ), 
        .Q(\IDinst/n11574 ) );
  nnd2s1 \IDinst/U11662  ( .DIN1(\IDinst/n11571 ), .DIN2(n1320), 
        .Q(\IDinst/n11573 ) );
  nnd2s1 \IDinst/U11661  ( .DIN1(\IDinst/n11568 ), .DIN2(n1350), 
        .Q(\IDinst/n11572 ) );
  nnd2s1 \IDinst/U11660  ( .DIN1(\IDinst/n11570 ), .DIN2(\IDinst/n11569 ), 
        .Q(\IDinst/n11571 ) );
  nnd2s1 \IDinst/U11659  ( .DIN1(\IDinst/RegFile[3][29] ), .DIN2(n1211), 
        .Q(\IDinst/n11570 ) );
  nnd2s1 \IDinst/U11658  ( .DIN1(\IDinst/RegFile[2][29] ), .DIN2(n1277), 
        .Q(\IDinst/n11569 ) );
  nnd2s1 \IDinst/U11657  ( .DIN1(\IDinst/n11567 ), .DIN2(\IDinst/n11566 ), 
        .Q(\IDinst/n11568 ) );
  nnd2s1 \IDinst/U11656  ( .DIN1(\IDinst/RegFile[1][29] ), .DIN2(n1212), 
        .Q(\IDinst/n11567 ) );
  nnd2s1 \IDinst/U11655  ( .DIN1(\IDinst/RegFile[0][29] ), .DIN2(n1277), 
        .Q(\IDinst/n11566 ) );
  nnd2s1 \IDinst/U11654  ( .DIN1(\IDinst/n11565 ), .DIN2(n535), 
        .Q(\IDinst/n8948 ) );
  nnd2s1 \IDinst/U11653  ( .DIN1(\IDinst/n11520 ), .DIN2(n634), 
        .Q(\IDinst/n8949 ) );
  nnd2s1 \IDinst/U11652  ( .DIN1(\IDinst/n11564 ), .DIN2(\IDinst/n11563 ), 
        .Q(\IDinst/n11565 ) );
  nnd2s1 \IDinst/U11651  ( .DIN1(\IDinst/n11562 ), .DIN2(n668), 
        .Q(\IDinst/n11564 ) );
  nnd2s1 \IDinst/U11650  ( .DIN1(\IDinst/n11541 ), .DIN2(n682), 
        .Q(\IDinst/n11563 ) );
  nnd2s1 \IDinst/U11649  ( .DIN1(\IDinst/n11561 ), .DIN2(\IDinst/n11560 ), 
        .Q(\IDinst/n11562 ) );
  nnd2s1 \IDinst/U11648  ( .DIN1(\IDinst/n11559 ), .DIN2(n1377), 
        .Q(\IDinst/n11561 ) );
  nnd2s1 \IDinst/U11647  ( .DIN1(\IDinst/n11550 ), .DIN2(n1367), 
        .Q(\IDinst/n11560 ) );
  nnd2s1 \IDinst/U11646  ( .DIN1(\IDinst/n11558 ), .DIN2(\IDinst/n11557 ), 
        .Q(\IDinst/n11559 ) );
  nnd2s1 \IDinst/U11645  ( .DIN1(\IDinst/n11556 ), .DIN2(n1320), 
        .Q(\IDinst/n11558 ) );
  nnd2s1 \IDinst/U11644  ( .DIN1(\IDinst/n11553 ), .DIN2(n1338), 
        .Q(\IDinst/n11557 ) );
  nnd2s1 \IDinst/U11643  ( .DIN1(\IDinst/n11555 ), .DIN2(\IDinst/n11554 ), 
        .Q(\IDinst/n11556 ) );
  nnd2s1 \IDinst/U11642  ( .DIN1(\IDinst/RegFile[31][28] ), .DIN2(n1212), 
        .Q(\IDinst/n11555 ) );
  nnd2s1 \IDinst/U11641  ( .DIN1(\IDinst/RegFile[30][28] ), .DIN2(n1277), 
        .Q(\IDinst/n11554 ) );
  nnd2s1 \IDinst/U11640  ( .DIN1(\IDinst/n11552 ), .DIN2(\IDinst/n11551 ), 
        .Q(\IDinst/n11553 ) );
  nnd2s1 \IDinst/U11639  ( .DIN1(\IDinst/RegFile[29][28] ), .DIN2(n1212), 
        .Q(\IDinst/n11552 ) );
  nnd2s1 \IDinst/U11638  ( .DIN1(\IDinst/RegFile[28][28] ), .DIN2(n1277), 
        .Q(\IDinst/n11551 ) );
  nnd2s1 \IDinst/U11637  ( .DIN1(\IDinst/n11549 ), .DIN2(\IDinst/n11548 ), 
        .Q(\IDinst/n11550 ) );
  nnd2s1 \IDinst/U11636  ( .DIN1(\IDinst/n11547 ), .DIN2(n1320), 
        .Q(\IDinst/n11549 ) );
  nnd2s1 \IDinst/U11635  ( .DIN1(\IDinst/n11544 ), .DIN2(n1337), 
        .Q(\IDinst/n11548 ) );
  nnd2s1 \IDinst/U11634  ( .DIN1(\IDinst/n11546 ), .DIN2(\IDinst/n11545 ), 
        .Q(\IDinst/n11547 ) );
  nnd2s1 \IDinst/U11633  ( .DIN1(\IDinst/RegFile[27][28] ), .DIN2(n1212), 
        .Q(\IDinst/n11546 ) );
  nnd2s1 \IDinst/U11632  ( .DIN1(\IDinst/RegFile[26][28] ), .DIN2(n1277), 
        .Q(\IDinst/n11545 ) );
  nnd2s1 \IDinst/U11631  ( .DIN1(\IDinst/n11543 ), .DIN2(\IDinst/n11542 ), 
        .Q(\IDinst/n11544 ) );
  nnd2s1 \IDinst/U11630  ( .DIN1(\IDinst/RegFile[25][28] ), .DIN2(n1212), 
        .Q(\IDinst/n11543 ) );
  nnd2s1 \IDinst/U11629  ( .DIN1(\IDinst/RegFile[24][28] ), .DIN2(n1277), 
        .Q(\IDinst/n11542 ) );
  nnd2s1 \IDinst/U11628  ( .DIN1(\IDinst/n11540 ), .DIN2(\IDinst/n11539 ), 
        .Q(\IDinst/n11541 ) );
  nnd2s1 \IDinst/U11627  ( .DIN1(\IDinst/n11538 ), .DIN2(n1378), 
        .Q(\IDinst/n11540 ) );
  nnd2s1 \IDinst/U11626  ( .DIN1(\IDinst/n11529 ), .DIN2(n1366), 
        .Q(\IDinst/n11539 ) );
  nnd2s1 \IDinst/U11625  ( .DIN1(\IDinst/n11537 ), .DIN2(\IDinst/n11536 ), 
        .Q(\IDinst/n11538 ) );
  nnd2s1 \IDinst/U11624  ( .DIN1(\IDinst/n11535 ), .DIN2(n1320), 
        .Q(\IDinst/n11537 ) );
  nnd2s1 \IDinst/U11623  ( .DIN1(\IDinst/n11532 ), .DIN2(n1350), 
        .Q(\IDinst/n11536 ) );
  nnd2s1 \IDinst/U11622  ( .DIN1(\IDinst/n11534 ), .DIN2(\IDinst/n11533 ), 
        .Q(\IDinst/n11535 ) );
  nnd2s1 \IDinst/U11621  ( .DIN1(\IDinst/RegFile[23][28] ), .DIN2(n1212), 
        .Q(\IDinst/n11534 ) );
  nnd2s1 \IDinst/U11620  ( .DIN1(\IDinst/RegFile[22][28] ), .DIN2(n1276), 
        .Q(\IDinst/n11533 ) );
  nnd2s1 \IDinst/U11619  ( .DIN1(\IDinst/n11531 ), .DIN2(\IDinst/n11530 ), 
        .Q(\IDinst/n11532 ) );
  nnd2s1 \IDinst/U11618  ( .DIN1(\IDinst/RegFile[21][28] ), .DIN2(n1212), 
        .Q(\IDinst/n11531 ) );
  nnd2s1 \IDinst/U11617  ( .DIN1(\IDinst/RegFile[20][28] ), .DIN2(n1276), 
        .Q(\IDinst/n11530 ) );
  nnd2s1 \IDinst/U11616  ( .DIN1(\IDinst/n11528 ), .DIN2(\IDinst/n11527 ), 
        .Q(\IDinst/n11529 ) );
  nnd2s1 \IDinst/U11615  ( .DIN1(\IDinst/n11526 ), .DIN2(n1320), 
        .Q(\IDinst/n11528 ) );
  nnd2s1 \IDinst/U11614  ( .DIN1(\IDinst/n11523 ), .DIN2(n1351), 
        .Q(\IDinst/n11527 ) );
  nnd2s1 \IDinst/U11613  ( .DIN1(\IDinst/n11525 ), .DIN2(\IDinst/n11524 ), 
        .Q(\IDinst/n11526 ) );
  nnd2s1 \IDinst/U11612  ( .DIN1(\IDinst/RegFile[19][28] ), .DIN2(n1212), 
        .Q(\IDinst/n11525 ) );
  nnd2s1 \IDinst/U11611  ( .DIN1(\IDinst/RegFile[18][28] ), .DIN2(n1276), 
        .Q(\IDinst/n11524 ) );
  nnd2s1 \IDinst/U11610  ( .DIN1(\IDinst/n11522 ), .DIN2(\IDinst/n11521 ), 
        .Q(\IDinst/n11523 ) );
  nnd2s1 \IDinst/U11609  ( .DIN1(\IDinst/RegFile[17][28] ), .DIN2(n1212), 
        .Q(\IDinst/n11522 ) );
  nnd2s1 \IDinst/U11608  ( .DIN1(\IDinst/RegFile[16][28] ), .DIN2(n1276), 
        .Q(\IDinst/n11521 ) );
  nnd2s1 \IDinst/U11607  ( .DIN1(\IDinst/n11519 ), .DIN2(\IDinst/n11518 ), 
        .Q(\IDinst/n11520 ) );
  nnd2s1 \IDinst/U11606  ( .DIN1(\IDinst/n11517 ), .DIN2(n666), 
        .Q(\IDinst/n11519 ) );
  nnd2s1 \IDinst/U11605  ( .DIN1(\IDinst/n11496 ), .DIN2(n680), 
        .Q(\IDinst/n11518 ) );
  nnd2s1 \IDinst/U11604  ( .DIN1(\IDinst/n11516 ), .DIN2(\IDinst/n11515 ), 
        .Q(\IDinst/n11517 ) );
  nnd2s1 \IDinst/U11603  ( .DIN1(\IDinst/n11514 ), .DIN2(n1380), 
        .Q(\IDinst/n11516 ) );
  nnd2s1 \IDinst/U11602  ( .DIN1(\IDinst/n11505 ), .DIN2(n1371), 
        .Q(\IDinst/n11515 ) );
  nnd2s1 \IDinst/U11601  ( .DIN1(\IDinst/n11513 ), .DIN2(\IDinst/n11512 ), 
        .Q(\IDinst/n11514 ) );
  nnd2s1 \IDinst/U11600  ( .DIN1(\IDinst/n11511 ), .DIN2(n1320), 
        .Q(\IDinst/n11513 ) );
  nnd2s1 \IDinst/U11599  ( .DIN1(\IDinst/n11508 ), .DIN2(n1355), 
        .Q(\IDinst/n11512 ) );
  nnd2s1 \IDinst/U11598  ( .DIN1(\IDinst/n11510 ), .DIN2(\IDinst/n11509 ), 
        .Q(\IDinst/n11511 ) );
  nnd2s1 \IDinst/U11597  ( .DIN1(\IDinst/RegFile[15][28] ), .DIN2(n1212), 
        .Q(\IDinst/n11510 ) );
  nnd2s1 \IDinst/U11596  ( .DIN1(\IDinst/RegFile[14][28] ), .DIN2(n1276), 
        .Q(\IDinst/n11509 ) );
  nnd2s1 \IDinst/U11595  ( .DIN1(\IDinst/n11507 ), .DIN2(\IDinst/n11506 ), 
        .Q(\IDinst/n11508 ) );
  nnd2s1 \IDinst/U11594  ( .DIN1(\IDinst/RegFile[13][28] ), .DIN2(n1212), 
        .Q(\IDinst/n11507 ) );
  nnd2s1 \IDinst/U11593  ( .DIN1(\IDinst/RegFile[12][28] ), .DIN2(n1276), 
        .Q(\IDinst/n11506 ) );
  nnd2s1 \IDinst/U11592  ( .DIN1(\IDinst/n11504 ), .DIN2(\IDinst/n11503 ), 
        .Q(\IDinst/n11505 ) );
  nnd2s1 \IDinst/U11591  ( .DIN1(\IDinst/n11502 ), .DIN2(n1320), 
        .Q(\IDinst/n11504 ) );
  nnd2s1 \IDinst/U11590  ( .DIN1(\IDinst/n11499 ), .DIN2(n1357), 
        .Q(\IDinst/n11503 ) );
  nnd2s1 \IDinst/U11589  ( .DIN1(\IDinst/n11501 ), .DIN2(\IDinst/n11500 ), 
        .Q(\IDinst/n11502 ) );
  nnd2s1 \IDinst/U11588  ( .DIN1(\IDinst/RegFile[11][28] ), .DIN2(n1212), 
        .Q(\IDinst/n11501 ) );
  nnd2s1 \IDinst/U11587  ( .DIN1(\IDinst/RegFile[10][28] ), .DIN2(n1276), 
        .Q(\IDinst/n11500 ) );
  nnd2s1 \IDinst/U11586  ( .DIN1(\IDinst/n11498 ), .DIN2(\IDinst/n11497 ), 
        .Q(\IDinst/n11499 ) );
  nnd2s1 \IDinst/U11585  ( .DIN1(\IDinst/RegFile[9][28] ), .DIN2(n1212), 
        .Q(\IDinst/n11498 ) );
  nnd2s1 \IDinst/U11584  ( .DIN1(\IDinst/RegFile[8][28] ), .DIN2(n1276), 
        .Q(\IDinst/n11497 ) );
  nnd2s1 \IDinst/U11583  ( .DIN1(\IDinst/n11495 ), .DIN2(\IDinst/n11494 ), 
        .Q(\IDinst/n11496 ) );
  nnd2s1 \IDinst/U11582  ( .DIN1(\IDinst/n11493 ), .DIN2(n1377), 
        .Q(\IDinst/n11495 ) );
  nnd2s1 \IDinst/U11581  ( .DIN1(\IDinst/n11484 ), .DIN2(n1365), 
        .Q(\IDinst/n11494 ) );
  nnd2s1 \IDinst/U11580  ( .DIN1(\IDinst/n11492 ), .DIN2(\IDinst/n11491 ), 
        .Q(\IDinst/n11493 ) );
  nnd2s1 \IDinst/U11579  ( .DIN1(\IDinst/n11490 ), .DIN2(n1320), 
        .Q(\IDinst/n11492 ) );
  nnd2s1 \IDinst/U11578  ( .DIN1(\IDinst/n11487 ), .DIN2(n1333), 
        .Q(\IDinst/n11491 ) );
  nnd2s1 \IDinst/U11577  ( .DIN1(\IDinst/n11489 ), .DIN2(\IDinst/n11488 ), 
        .Q(\IDinst/n11490 ) );
  nnd2s1 \IDinst/U11576  ( .DIN1(\IDinst/RegFile[7][28] ), .DIN2(n1213), 
        .Q(\IDinst/n11489 ) );
  nnd2s1 \IDinst/U11575  ( .DIN1(\IDinst/RegFile[6][28] ), .DIN2(n1275), 
        .Q(\IDinst/n11488 ) );
  nnd2s1 \IDinst/U11574  ( .DIN1(\IDinst/n11486 ), .DIN2(\IDinst/n11485 ), 
        .Q(\IDinst/n11487 ) );
  nnd2s1 \IDinst/U11573  ( .DIN1(\IDinst/RegFile[5][28] ), .DIN2(n1213), 
        .Q(\IDinst/n11486 ) );
  nnd2s1 \IDinst/U11572  ( .DIN1(\IDinst/RegFile[4][28] ), .DIN2(n1275), 
        .Q(\IDinst/n11485 ) );
  nnd2s1 \IDinst/U11571  ( .DIN1(\IDinst/n11483 ), .DIN2(\IDinst/n11482 ), 
        .Q(\IDinst/n11484 ) );
  nnd2s1 \IDinst/U11570  ( .DIN1(\IDinst/n11481 ), .DIN2(n1320), 
        .Q(\IDinst/n11483 ) );
  nnd2s1 \IDinst/U11569  ( .DIN1(\IDinst/n11478 ), .DIN2(n1354), 
        .Q(\IDinst/n11482 ) );
  nnd2s1 \IDinst/U11568  ( .DIN1(\IDinst/n11480 ), .DIN2(\IDinst/n11479 ), 
        .Q(\IDinst/n11481 ) );
  nnd2s1 \IDinst/U11567  ( .DIN1(\IDinst/RegFile[3][28] ), .DIN2(n1213), 
        .Q(\IDinst/n11480 ) );
  nnd2s1 \IDinst/U11566  ( .DIN1(\IDinst/RegFile[2][28] ), .DIN2(n1275), 
        .Q(\IDinst/n11479 ) );
  nnd2s1 \IDinst/U11565  ( .DIN1(\IDinst/n11477 ), .DIN2(\IDinst/n11476 ), 
        .Q(\IDinst/n11478 ) );
  nnd2s1 \IDinst/U11564  ( .DIN1(\IDinst/RegFile[1][28] ), .DIN2(n1213), 
        .Q(\IDinst/n11477 ) );
  nnd2s1 \IDinst/U11563  ( .DIN1(\IDinst/RegFile[0][28] ), .DIN2(n1275), 
        .Q(\IDinst/n11476 ) );
  nnd2s1 \IDinst/U11562  ( .DIN1(\IDinst/n11475 ), .DIN2(n535), 
        .Q(\IDinst/n8946 ) );
  nnd2s1 \IDinst/U11561  ( .DIN1(\IDinst/n11430 ), .DIN2(n533), 
        .Q(\IDinst/n8947 ) );
  nnd2s1 \IDinst/U11560  ( .DIN1(\IDinst/n11474 ), .DIN2(\IDinst/n11473 ), 
        .Q(\IDinst/n11475 ) );
  nnd2s1 \IDinst/U11559  ( .DIN1(\IDinst/n11472 ), .DIN2(n667), 
        .Q(\IDinst/n11474 ) );
  nnd2s1 \IDinst/U11558  ( .DIN1(\IDinst/n11451 ), .DIN2(n683), 
        .Q(\IDinst/n11473 ) );
  nnd2s1 \IDinst/U11557  ( .DIN1(\IDinst/n11471 ), .DIN2(\IDinst/n11470 ), 
        .Q(\IDinst/n11472 ) );
  nnd2s1 \IDinst/U11556  ( .DIN1(\IDinst/n11469 ), .DIN2(n1376), 
        .Q(\IDinst/n11471 ) );
  nnd2s1 \IDinst/U11555  ( .DIN1(\IDinst/n11460 ), .DIN2(n1367), 
        .Q(\IDinst/n11470 ) );
  nnd2s1 \IDinst/U11554  ( .DIN1(\IDinst/n11468 ), .DIN2(\IDinst/n11467 ), 
        .Q(\IDinst/n11469 ) );
  nnd2s1 \IDinst/U11553  ( .DIN1(\IDinst/n11466 ), .DIN2(n1320), 
        .Q(\IDinst/n11468 ) );
  nnd2s1 \IDinst/U11552  ( .DIN1(\IDinst/n11463 ), .DIN2(n1360), 
        .Q(\IDinst/n11467 ) );
  nnd2s1 \IDinst/U11551  ( .DIN1(\IDinst/n11465 ), .DIN2(\IDinst/n11464 ), 
        .Q(\IDinst/n11466 ) );
  nnd2s1 \IDinst/U11550  ( .DIN1(\IDinst/RegFile[31][27] ), .DIN2(n1213), 
        .Q(\IDinst/n11465 ) );
  nnd2s1 \IDinst/U11549  ( .DIN1(\IDinst/RegFile[30][27] ), .DIN2(n1275), 
        .Q(\IDinst/n11464 ) );
  nnd2s1 \IDinst/U11548  ( .DIN1(\IDinst/n11462 ), .DIN2(\IDinst/n11461 ), 
        .Q(\IDinst/n11463 ) );
  nnd2s1 \IDinst/U11547  ( .DIN1(\IDinst/RegFile[29][27] ), .DIN2(n1213), 
        .Q(\IDinst/n11462 ) );
  nnd2s1 \IDinst/U11546  ( .DIN1(\IDinst/RegFile[28][27] ), .DIN2(n1275), 
        .Q(\IDinst/n11461 ) );
  nnd2s1 \IDinst/U11545  ( .DIN1(\IDinst/n11459 ), .DIN2(\IDinst/n11458 ), 
        .Q(\IDinst/n11460 ) );
  nnd2s1 \IDinst/U11544  ( .DIN1(\IDinst/n11457 ), .DIN2(n1319), 
        .Q(\IDinst/n11459 ) );
  nnd2s1 \IDinst/U11543  ( .DIN1(\IDinst/n11454 ), .DIN2(n1351), 
        .Q(\IDinst/n11458 ) );
  nnd2s1 \IDinst/U11542  ( .DIN1(\IDinst/n11456 ), .DIN2(\IDinst/n11455 ), 
        .Q(\IDinst/n11457 ) );
  nnd2s1 \IDinst/U11541  ( .DIN1(\IDinst/RegFile[27][27] ), .DIN2(n1213), 
        .Q(\IDinst/n11456 ) );
  nnd2s1 \IDinst/U11540  ( .DIN1(\IDinst/RegFile[26][27] ), .DIN2(n1275), 
        .Q(\IDinst/n11455 ) );
  nnd2s1 \IDinst/U11539  ( .DIN1(\IDinst/n11453 ), .DIN2(\IDinst/n11452 ), 
        .Q(\IDinst/n11454 ) );
  nnd2s1 \IDinst/U11538  ( .DIN1(\IDinst/RegFile[25][27] ), .DIN2(n1213), 
        .Q(\IDinst/n11453 ) );
  nnd2s1 \IDinst/U11537  ( .DIN1(\IDinst/RegFile[24][27] ), .DIN2(n1275), 
        .Q(\IDinst/n11452 ) );
  nnd2s1 \IDinst/U11536  ( .DIN1(\IDinst/n11450 ), .DIN2(\IDinst/n11449 ), 
        .Q(\IDinst/n11451 ) );
  nnd2s1 \IDinst/U11535  ( .DIN1(\IDinst/n11448 ), .DIN2(n1378), 
        .Q(\IDinst/n11450 ) );
  nnd2s1 \IDinst/U11534  ( .DIN1(\IDinst/n11439 ), .DIN2(n1371), 
        .Q(\IDinst/n11449 ) );
  nnd2s1 \IDinst/U11533  ( .DIN1(\IDinst/n11447 ), .DIN2(\IDinst/n11446 ), 
        .Q(\IDinst/n11448 ) );
  nnd2s1 \IDinst/U11532  ( .DIN1(\IDinst/n11445 ), .DIN2(n1319), 
        .Q(\IDinst/n11447 ) );
  nnd2s1 \IDinst/U11531  ( .DIN1(\IDinst/n11442 ), .DIN2(n1351), 
        .Q(\IDinst/n11446 ) );
  nnd2s1 \IDinst/U11530  ( .DIN1(\IDinst/n11444 ), .DIN2(\IDinst/n11443 ), 
        .Q(\IDinst/n11445 ) );
  nnd2s1 \IDinst/U11529  ( .DIN1(\IDinst/RegFile[23][27] ), .DIN2(n1213), 
        .Q(\IDinst/n11444 ) );
  nnd2s1 \IDinst/U11528  ( .DIN1(\IDinst/RegFile[22][27] ), .DIN2(n1275), 
        .Q(\IDinst/n11443 ) );
  nnd2s1 \IDinst/U11527  ( .DIN1(\IDinst/n11441 ), .DIN2(\IDinst/n11440 ), 
        .Q(\IDinst/n11442 ) );
  nnd2s1 \IDinst/U11526  ( .DIN1(\IDinst/RegFile[21][27] ), .DIN2(n1213), 
        .Q(\IDinst/n11441 ) );
  nnd2s1 \IDinst/U11525  ( .DIN1(\IDinst/RegFile[20][27] ), .DIN2(n1274), 
        .Q(\IDinst/n11440 ) );
  nnd2s1 \IDinst/U11524  ( .DIN1(\IDinst/n11438 ), .DIN2(\IDinst/n11437 ), 
        .Q(\IDinst/n11439 ) );
  nnd2s1 \IDinst/U11523  ( .DIN1(\IDinst/n11436 ), .DIN2(n1319), 
        .Q(\IDinst/n11438 ) );
  nnd2s1 \IDinst/U11522  ( .DIN1(\IDinst/n11433 ), .DIN2(n1351), 
        .Q(\IDinst/n11437 ) );
  nnd2s1 \IDinst/U11521  ( .DIN1(\IDinst/n11435 ), .DIN2(\IDinst/n11434 ), 
        .Q(\IDinst/n11436 ) );
  nnd2s1 \IDinst/U11520  ( .DIN1(\IDinst/RegFile[19][27] ), .DIN2(n1213), 
        .Q(\IDinst/n11435 ) );
  nnd2s1 \IDinst/U11519  ( .DIN1(\IDinst/RegFile[18][27] ), .DIN2(n1274), 
        .Q(\IDinst/n11434 ) );
  nnd2s1 \IDinst/U11518  ( .DIN1(\IDinst/n11432 ), .DIN2(\IDinst/n11431 ), 
        .Q(\IDinst/n11433 ) );
  nnd2s1 \IDinst/U11517  ( .DIN1(\IDinst/RegFile[17][27] ), .DIN2(n1213), 
        .Q(\IDinst/n11432 ) );
  nnd2s1 \IDinst/U11516  ( .DIN1(\IDinst/RegFile[16][27] ), .DIN2(n1274), 
        .Q(\IDinst/n11431 ) );
  nnd2s1 \IDinst/U11515  ( .DIN1(\IDinst/n11429 ), .DIN2(\IDinst/n11428 ), 
        .Q(\IDinst/n11430 ) );
  nnd2s1 \IDinst/U11514  ( .DIN1(\IDinst/n11427 ), .DIN2(n665), 
        .Q(\IDinst/n11429 ) );
  nnd2s1 \IDinst/U11513  ( .DIN1(\IDinst/n11406 ), .DIN2(n682), 
        .Q(\IDinst/n11428 ) );
  nnd2s1 \IDinst/U11512  ( .DIN1(\IDinst/n11426 ), .DIN2(\IDinst/n11425 ), 
        .Q(\IDinst/n11427 ) );
  nnd2s1 \IDinst/U11511  ( .DIN1(\IDinst/n11424 ), .DIN2(n1374), 
        .Q(\IDinst/n11426 ) );
  nnd2s1 \IDinst/U11510  ( .DIN1(\IDinst/n11415 ), .DIN2(n1370), 
        .Q(\IDinst/n11425 ) );
  nnd2s1 \IDinst/U11509  ( .DIN1(\IDinst/n11423 ), .DIN2(\IDinst/n11422 ), 
        .Q(\IDinst/n11424 ) );
  nnd2s1 \IDinst/U11508  ( .DIN1(\IDinst/n11421 ), .DIN2(n1319), 
        .Q(\IDinst/n11423 ) );
  nnd2s1 \IDinst/U11507  ( .DIN1(\IDinst/n11418 ), .DIN2(n1351), 
        .Q(\IDinst/n11422 ) );
  nnd2s1 \IDinst/U11506  ( .DIN1(\IDinst/n11420 ), .DIN2(\IDinst/n11419 ), 
        .Q(\IDinst/n11421 ) );
  nnd2s1 \IDinst/U11505  ( .DIN1(\IDinst/RegFile[15][27] ), .DIN2(n1214), 
        .Q(\IDinst/n11420 ) );
  nnd2s1 \IDinst/U11504  ( .DIN1(\IDinst/RegFile[14][27] ), .DIN2(n1274), 
        .Q(\IDinst/n11419 ) );
  nnd2s1 \IDinst/U11503  ( .DIN1(\IDinst/n11417 ), .DIN2(\IDinst/n11416 ), 
        .Q(\IDinst/n11418 ) );
  nnd2s1 \IDinst/U11502  ( .DIN1(\IDinst/RegFile[13][27] ), .DIN2(n1214), 
        .Q(\IDinst/n11417 ) );
  nnd2s1 \IDinst/U11501  ( .DIN1(\IDinst/RegFile[12][27] ), .DIN2(n1274), 
        .Q(\IDinst/n11416 ) );
  nnd2s1 \IDinst/U11500  ( .DIN1(\IDinst/n11414 ), .DIN2(\IDinst/n11413 ), 
        .Q(\IDinst/n11415 ) );
  nnd2s1 \IDinst/U11499  ( .DIN1(\IDinst/n11412 ), .DIN2(n1319), 
        .Q(\IDinst/n11414 ) );
  nnd2s1 \IDinst/U11498  ( .DIN1(\IDinst/n11409 ), .DIN2(n1351), 
        .Q(\IDinst/n11413 ) );
  nnd2s1 \IDinst/U11497  ( .DIN1(\IDinst/n11411 ), .DIN2(\IDinst/n11410 ), 
        .Q(\IDinst/n11412 ) );
  nnd2s1 \IDinst/U11496  ( .DIN1(\IDinst/RegFile[11][27] ), .DIN2(n1214), 
        .Q(\IDinst/n11411 ) );
  nnd2s1 \IDinst/U11495  ( .DIN1(\IDinst/RegFile[10][27] ), .DIN2(n1274), 
        .Q(\IDinst/n11410 ) );
  nnd2s1 \IDinst/U11494  ( .DIN1(\IDinst/n11408 ), .DIN2(\IDinst/n11407 ), 
        .Q(\IDinst/n11409 ) );
  nnd2s1 \IDinst/U11493  ( .DIN1(\IDinst/RegFile[9][27] ), .DIN2(n1214), 
        .Q(\IDinst/n11408 ) );
  nnd2s1 \IDinst/U11492  ( .DIN1(\IDinst/RegFile[8][27] ), .DIN2(n1274), 
        .Q(\IDinst/n11407 ) );
  nnd2s1 \IDinst/U11491  ( .DIN1(\IDinst/n11405 ), .DIN2(\IDinst/n11404 ), 
        .Q(\IDinst/n11406 ) );
  nnd2s1 \IDinst/U11490  ( .DIN1(\IDinst/n11403 ), .DIN2(n1378), 
        .Q(\IDinst/n11405 ) );
  nnd2s1 \IDinst/U11489  ( .DIN1(\IDinst/n11394 ), .DIN2(n1369), 
        .Q(\IDinst/n11404 ) );
  nnd2s1 \IDinst/U11488  ( .DIN1(\IDinst/n11402 ), .DIN2(\IDinst/n11401 ), 
        .Q(\IDinst/n11403 ) );
  nnd2s1 \IDinst/U11487  ( .DIN1(\IDinst/n11400 ), .DIN2(n1319), 
        .Q(\IDinst/n11402 ) );
  nnd2s1 \IDinst/U11486  ( .DIN1(\IDinst/n11397 ), .DIN2(n1351), 
        .Q(\IDinst/n11401 ) );
  nnd2s1 \IDinst/U11485  ( .DIN1(\IDinst/n11399 ), .DIN2(\IDinst/n11398 ), 
        .Q(\IDinst/n11400 ) );
  nnd2s1 \IDinst/U11484  ( .DIN1(\IDinst/RegFile[7][27] ), .DIN2(n1214), 
        .Q(\IDinst/n11399 ) );
  nnd2s1 \IDinst/U11483  ( .DIN1(\IDinst/RegFile[6][27] ), .DIN2(n1274), 
        .Q(\IDinst/n11398 ) );
  nnd2s1 \IDinst/U11482  ( .DIN1(\IDinst/n11396 ), .DIN2(\IDinst/n11395 ), 
        .Q(\IDinst/n11397 ) );
  nnd2s1 \IDinst/U11481  ( .DIN1(\IDinst/RegFile[5][27] ), .DIN2(n1214), 
        .Q(\IDinst/n11396 ) );
  nnd2s1 \IDinst/U11480  ( .DIN1(\IDinst/RegFile[4][27] ), .DIN2(n1274), 
        .Q(\IDinst/n11395 ) );
  nnd2s1 \IDinst/U11479  ( .DIN1(\IDinst/n11393 ), .DIN2(\IDinst/n11392 ), 
        .Q(\IDinst/n11394 ) );
  nnd2s1 \IDinst/U11478  ( .DIN1(\IDinst/n11391 ), .DIN2(n1319), 
        .Q(\IDinst/n11393 ) );
  nnd2s1 \IDinst/U11477  ( .DIN1(\IDinst/n11388 ), .DIN2(n1351), 
        .Q(\IDinst/n11392 ) );
  nnd2s1 \IDinst/U11476  ( .DIN1(\IDinst/n11390 ), .DIN2(\IDinst/n11389 ), 
        .Q(\IDinst/n11391 ) );
  nnd2s1 \IDinst/U11475  ( .DIN1(\IDinst/RegFile[3][27] ), .DIN2(n1214), 
        .Q(\IDinst/n11390 ) );
  nnd2s1 \IDinst/U11474  ( .DIN1(\IDinst/RegFile[2][27] ), .DIN2(n1273), 
        .Q(\IDinst/n11389 ) );
  nnd2s1 \IDinst/U11473  ( .DIN1(\IDinst/n11387 ), .DIN2(\IDinst/n11386 ), 
        .Q(\IDinst/n11388 ) );
  nnd2s1 \IDinst/U11472  ( .DIN1(\IDinst/RegFile[1][27] ), .DIN2(n1214), 
        .Q(\IDinst/n11387 ) );
  nnd2s1 \IDinst/U11471  ( .DIN1(\IDinst/RegFile[0][27] ), .DIN2(n1273), 
        .Q(\IDinst/n11386 ) );
  nnd2s1 \IDinst/U11470  ( .DIN1(\IDinst/n11385 ), .DIN2(n534), 
        .Q(\IDinst/n8944 ) );
  nnd2s1 \IDinst/U11469  ( .DIN1(\IDinst/n11340 ), .DIN2(n634), 
        .Q(\IDinst/n8945 ) );
  nnd2s1 \IDinst/U11468  ( .DIN1(\IDinst/n11384 ), .DIN2(\IDinst/n11383 ), 
        .Q(\IDinst/n11385 ) );
  nnd2s1 \IDinst/U11467  ( .DIN1(\IDinst/n11382 ), .DIN2(n668), 
        .Q(\IDinst/n11384 ) );
  nnd2s1 \IDinst/U11466  ( .DIN1(\IDinst/n11361 ), .DIN2(n680), 
        .Q(\IDinst/n11383 ) );
  nnd2s1 \IDinst/U11465  ( .DIN1(\IDinst/n11381 ), .DIN2(\IDinst/n11380 ), 
        .Q(\IDinst/n11382 ) );
  nnd2s1 \IDinst/U11464  ( .DIN1(\IDinst/n11379 ), .DIN2(n1378), 
        .Q(\IDinst/n11381 ) );
  nnd2s1 \IDinst/U11463  ( .DIN1(\IDinst/n11370 ), .DIN2(n1368), 
        .Q(\IDinst/n11380 ) );
  nnd2s1 \IDinst/U11462  ( .DIN1(\IDinst/n11378 ), .DIN2(\IDinst/n11377 ), 
        .Q(\IDinst/n11379 ) );
  nnd2s1 \IDinst/U11461  ( .DIN1(\IDinst/n11376 ), .DIN2(n1319), 
        .Q(\IDinst/n11378 ) );
  nnd2s1 \IDinst/U11460  ( .DIN1(\IDinst/n11373 ), .DIN2(n1351), 
        .Q(\IDinst/n11377 ) );
  nnd2s1 \IDinst/U11459  ( .DIN1(\IDinst/n11375 ), .DIN2(\IDinst/n11374 ), 
        .Q(\IDinst/n11376 ) );
  nnd2s1 \IDinst/U11458  ( .DIN1(\IDinst/RegFile[31][26] ), .DIN2(n1214), 
        .Q(\IDinst/n11375 ) );
  nnd2s1 \IDinst/U11457  ( .DIN1(\IDinst/RegFile[30][26] ), .DIN2(n1273), 
        .Q(\IDinst/n11374 ) );
  nnd2s1 \IDinst/U11456  ( .DIN1(\IDinst/n11372 ), .DIN2(\IDinst/n11371 ), 
        .Q(\IDinst/n11373 ) );
  nnd2s1 \IDinst/U11455  ( .DIN1(\IDinst/RegFile[29][26] ), .DIN2(n1214), 
        .Q(\IDinst/n11372 ) );
  nnd2s1 \IDinst/U11454  ( .DIN1(\IDinst/RegFile[28][26] ), .DIN2(n1273), 
        .Q(\IDinst/n11371 ) );
  nnd2s1 \IDinst/U11453  ( .DIN1(\IDinst/n11369 ), .DIN2(\IDinst/n11368 ), 
        .Q(\IDinst/n11370 ) );
  nnd2s1 \IDinst/U11452  ( .DIN1(\IDinst/n11367 ), .DIN2(n1319), 
        .Q(\IDinst/n11369 ) );
  nnd2s1 \IDinst/U11451  ( .DIN1(\IDinst/n11364 ), .DIN2(n1351), 
        .Q(\IDinst/n11368 ) );
  nnd2s1 \IDinst/U11450  ( .DIN1(\IDinst/n11366 ), .DIN2(\IDinst/n11365 ), 
        .Q(\IDinst/n11367 ) );
  nnd2s1 \IDinst/U11449  ( .DIN1(\IDinst/RegFile[27][26] ), .DIN2(n1214), 
        .Q(\IDinst/n11366 ) );
  nnd2s1 \IDinst/U11448  ( .DIN1(\IDinst/RegFile[26][26] ), .DIN2(n1273), 
        .Q(\IDinst/n11365 ) );
  nnd2s1 \IDinst/U11447  ( .DIN1(\IDinst/n11363 ), .DIN2(\IDinst/n11362 ), 
        .Q(\IDinst/n11364 ) );
  nnd2s1 \IDinst/U11446  ( .DIN1(\IDinst/RegFile[25][26] ), .DIN2(n1214), 
        .Q(\IDinst/n11363 ) );
  nnd2s1 \IDinst/U11445  ( .DIN1(\IDinst/RegFile[24][26] ), .DIN2(n1273), 
        .Q(\IDinst/n11362 ) );
  nnd2s1 \IDinst/U11444  ( .DIN1(\IDinst/n11360 ), .DIN2(\IDinst/n11359 ), 
        .Q(\IDinst/n11361 ) );
  nnd2s1 \IDinst/U11443  ( .DIN1(\IDinst/n11358 ), .DIN2(n1378), 
        .Q(\IDinst/n11360 ) );
  nnd2s1 \IDinst/U11442  ( .DIN1(\IDinst/n11349 ), .DIN2(n1371), 
        .Q(\IDinst/n11359 ) );
  nnd2s1 \IDinst/U11441  ( .DIN1(\IDinst/n11357 ), .DIN2(\IDinst/n11356 ), 
        .Q(\IDinst/n11358 ) );
  nnd2s1 \IDinst/U11440  ( .DIN1(\IDinst/n11355 ), .DIN2(n1319), 
        .Q(\IDinst/n11357 ) );
  nnd2s1 \IDinst/U11439  ( .DIN1(\IDinst/n11352 ), .DIN2(n1352), 
        .Q(\IDinst/n11356 ) );
  nnd2s1 \IDinst/U11438  ( .DIN1(\IDinst/n11354 ), .DIN2(\IDinst/n11353 ), 
        .Q(\IDinst/n11355 ) );
  nnd2s1 \IDinst/U11437  ( .DIN1(\IDinst/RegFile[23][26] ), .DIN2(n1214), 
        .Q(\IDinst/n11354 ) );
  nnd2s1 \IDinst/U11436  ( .DIN1(\IDinst/RegFile[22][26] ), .DIN2(n1273), 
        .Q(\IDinst/n11353 ) );
  nnd2s1 \IDinst/U11435  ( .DIN1(\IDinst/n11351 ), .DIN2(\IDinst/n11350 ), 
        .Q(\IDinst/n11352 ) );
  nnd2s1 \IDinst/U11434  ( .DIN1(\IDinst/RegFile[21][26] ), .DIN2(n1215), 
        .Q(\IDinst/n11351 ) );
  nnd2s1 \IDinst/U11433  ( .DIN1(\IDinst/RegFile[20][26] ), .DIN2(n1273), 
        .Q(\IDinst/n11350 ) );
  nnd2s1 \IDinst/U11432  ( .DIN1(\IDinst/n11348 ), .DIN2(\IDinst/n11347 ), 
        .Q(\IDinst/n11349 ) );
  nnd2s1 \IDinst/U11431  ( .DIN1(\IDinst/n11346 ), .DIN2(n1319), 
        .Q(\IDinst/n11348 ) );
  nnd2s1 \IDinst/U11430  ( .DIN1(\IDinst/n11343 ), .DIN2(n1352), 
        .Q(\IDinst/n11347 ) );
  nnd2s1 \IDinst/U11429  ( .DIN1(\IDinst/n11345 ), .DIN2(\IDinst/n11344 ), 
        .Q(\IDinst/n11346 ) );
  nnd2s1 \IDinst/U11428  ( .DIN1(\IDinst/RegFile[19][26] ), .DIN2(n1215), 
        .Q(\IDinst/n11345 ) );
  nnd2s1 \IDinst/U11427  ( .DIN1(\IDinst/RegFile[18][26] ), .DIN2(n1273), 
        .Q(\IDinst/n11344 ) );
  nnd2s1 \IDinst/U11426  ( .DIN1(\IDinst/n11342 ), .DIN2(\IDinst/n11341 ), 
        .Q(\IDinst/n11343 ) );
  nnd2s1 \IDinst/U11425  ( .DIN1(\IDinst/RegFile[17][26] ), .DIN2(n1215), 
        .Q(\IDinst/n11342 ) );
  nnd2s1 \IDinst/U11424  ( .DIN1(\IDinst/RegFile[16][26] ), .DIN2(n1272), 
        .Q(\IDinst/n11341 ) );
  nnd2s1 \IDinst/U11423  ( .DIN1(\IDinst/n11339 ), .DIN2(\IDinst/n11338 ), 
        .Q(\IDinst/n11340 ) );
  nnd2s1 \IDinst/U11422  ( .DIN1(\IDinst/n11337 ), .DIN2(n666), 
        .Q(\IDinst/n11339 ) );
  nnd2s1 \IDinst/U11421  ( .DIN1(\IDinst/n11316 ), .DIN2(n681), 
        .Q(\IDinst/n11338 ) );
  nnd2s1 \IDinst/U11420  ( .DIN1(\IDinst/n11336 ), .DIN2(\IDinst/n11335 ), 
        .Q(\IDinst/n11337 ) );
  nnd2s1 \IDinst/U11419  ( .DIN1(\IDinst/n11334 ), .DIN2(n1374), 
        .Q(\IDinst/n11336 ) );
  nnd2s1 \IDinst/U11418  ( .DIN1(\IDinst/n11325 ), .DIN2(n1371), 
        .Q(\IDinst/n11335 ) );
  nnd2s1 \IDinst/U11417  ( .DIN1(\IDinst/n11333 ), .DIN2(\IDinst/n11332 ), 
        .Q(\IDinst/n11334 ) );
  nnd2s1 \IDinst/U11416  ( .DIN1(\IDinst/n11331 ), .DIN2(n1319), 
        .Q(\IDinst/n11333 ) );
  nnd2s1 \IDinst/U11415  ( .DIN1(\IDinst/n11328 ), .DIN2(n1352), 
        .Q(\IDinst/n11332 ) );
  nnd2s1 \IDinst/U11414  ( .DIN1(\IDinst/n11330 ), .DIN2(\IDinst/n11329 ), 
        .Q(\IDinst/n11331 ) );
  nnd2s1 \IDinst/U11413  ( .DIN1(\IDinst/RegFile[15][26] ), .DIN2(n1215), 
        .Q(\IDinst/n11330 ) );
  nnd2s1 \IDinst/U11412  ( .DIN1(\IDinst/RegFile[14][26] ), .DIN2(n1272), 
        .Q(\IDinst/n11329 ) );
  nnd2s1 \IDinst/U11411  ( .DIN1(\IDinst/n11327 ), .DIN2(\IDinst/n11326 ), 
        .Q(\IDinst/n11328 ) );
  nnd2s1 \IDinst/U11410  ( .DIN1(\IDinst/RegFile[13][26] ), .DIN2(n1215), 
        .Q(\IDinst/n11327 ) );
  nnd2s1 \IDinst/U11409  ( .DIN1(\IDinst/RegFile[12][26] ), .DIN2(n1272), 
        .Q(\IDinst/n11326 ) );
  nnd2s1 \IDinst/U11408  ( .DIN1(\IDinst/n11324 ), .DIN2(\IDinst/n11323 ), 
        .Q(\IDinst/n11325 ) );
  nnd2s1 \IDinst/U11407  ( .DIN1(\IDinst/n11322 ), .DIN2(n1319), 
        .Q(\IDinst/n11324 ) );
  nnd2s1 \IDinst/U11406  ( .DIN1(\IDinst/n11319 ), .DIN2(n1352), 
        .Q(\IDinst/n11323 ) );
  nnd2s1 \IDinst/U11405  ( .DIN1(\IDinst/n11321 ), .DIN2(\IDinst/n11320 ), 
        .Q(\IDinst/n11322 ) );
  nnd2s1 \IDinst/U11404  ( .DIN1(\IDinst/RegFile[11][26] ), .DIN2(n1215), 
        .Q(\IDinst/n11321 ) );
  nnd2s1 \IDinst/U11403  ( .DIN1(\IDinst/RegFile[10][26] ), .DIN2(n1272), 
        .Q(\IDinst/n11320 ) );
  nnd2s1 \IDinst/U11402  ( .DIN1(\IDinst/n11318 ), .DIN2(\IDinst/n11317 ), 
        .Q(\IDinst/n11319 ) );
  nnd2s1 \IDinst/U11401  ( .DIN1(\IDinst/RegFile[9][26] ), .DIN2(n1215), 
        .Q(\IDinst/n11318 ) );
  nnd2s1 \IDinst/U11400  ( .DIN1(\IDinst/RegFile[8][26] ), .DIN2(n1272), 
        .Q(\IDinst/n11317 ) );
  nnd2s1 \IDinst/U11399  ( .DIN1(\IDinst/n11315 ), .DIN2(\IDinst/n11314 ), 
        .Q(\IDinst/n11316 ) );
  nnd2s1 \IDinst/U11398  ( .DIN1(\IDinst/n11313 ), .DIN2(\IDinst/N46 ), 
        .Q(\IDinst/n11315 ) );
  nnd2s1 \IDinst/U11397  ( .DIN1(\IDinst/n11304 ), .DIN2(n1371), 
        .Q(\IDinst/n11314 ) );
  nnd2s1 \IDinst/U11396  ( .DIN1(\IDinst/n11312 ), .DIN2(\IDinst/n11311 ), 
        .Q(\IDinst/n11313 ) );
  nnd2s1 \IDinst/U11395  ( .DIN1(\IDinst/n11310 ), .DIN2(n1318), 
        .Q(\IDinst/n11312 ) );
  nnd2s1 \IDinst/U11394  ( .DIN1(\IDinst/n11307 ), .DIN2(n1352), 
        .Q(\IDinst/n11311 ) );
  nnd2s1 \IDinst/U11393  ( .DIN1(\IDinst/n11309 ), .DIN2(\IDinst/n11308 ), 
        .Q(\IDinst/n11310 ) );
  nnd2s1 \IDinst/U11392  ( .DIN1(\IDinst/RegFile[7][26] ), .DIN2(n1215), 
        .Q(\IDinst/n11309 ) );
  nnd2s1 \IDinst/U11391  ( .DIN1(\IDinst/RegFile[6][26] ), .DIN2(n1272), 
        .Q(\IDinst/n11308 ) );
  nnd2s1 \IDinst/U11390  ( .DIN1(\IDinst/n11306 ), .DIN2(\IDinst/n11305 ), 
        .Q(\IDinst/n11307 ) );
  nnd2s1 \IDinst/U11389  ( .DIN1(\IDinst/RegFile[5][26] ), .DIN2(n1215), 
        .Q(\IDinst/n11306 ) );
  nnd2s1 \IDinst/U11388  ( .DIN1(\IDinst/RegFile[4][26] ), .DIN2(n1272), 
        .Q(\IDinst/n11305 ) );
  nnd2s1 \IDinst/U11387  ( .DIN1(\IDinst/n11303 ), .DIN2(\IDinst/n11302 ), 
        .Q(\IDinst/n11304 ) );
  nnd2s1 \IDinst/U11386  ( .DIN1(\IDinst/n11301 ), .DIN2(n1318), 
        .Q(\IDinst/n11303 ) );
  nnd2s1 \IDinst/U11385  ( .DIN1(\IDinst/n11298 ), .DIN2(n1352), 
        .Q(\IDinst/n11302 ) );
  nnd2s1 \IDinst/U11384  ( .DIN1(\IDinst/n11300 ), .DIN2(\IDinst/n11299 ), 
        .Q(\IDinst/n11301 ) );
  nnd2s1 \IDinst/U11383  ( .DIN1(\IDinst/RegFile[3][26] ), .DIN2(n1215), 
        .Q(\IDinst/n11300 ) );
  nnd2s1 \IDinst/U11382  ( .DIN1(\IDinst/RegFile[2][26] ), .DIN2(n1272), 
        .Q(\IDinst/n11299 ) );
  nnd2s1 \IDinst/U11381  ( .DIN1(\IDinst/n11297 ), .DIN2(\IDinst/n11296 ), 
        .Q(\IDinst/n11298 ) );
  nnd2s1 \IDinst/U11380  ( .DIN1(\IDinst/RegFile[1][26] ), .DIN2(n1215), 
        .Q(\IDinst/n11297 ) );
  nnd2s1 \IDinst/U11379  ( .DIN1(\IDinst/RegFile[0][26] ), .DIN2(n1272), 
        .Q(\IDinst/n11296 ) );
  nnd2s1 \IDinst/U11378  ( .DIN1(\IDinst/n11295 ), .DIN2(\IDinst/N48 ), 
        .Q(\IDinst/n8942 ) );
  nnd2s1 \IDinst/U11377  ( .DIN1(\IDinst/n11250 ), .DIN2(n533), 
        .Q(\IDinst/n8943 ) );
  nnd2s1 \IDinst/U11376  ( .DIN1(\IDinst/n11294 ), .DIN2(\IDinst/n11293 ), 
        .Q(\IDinst/n11295 ) );
  nnd2s1 \IDinst/U11375  ( .DIN1(\IDinst/n11292 ), .DIN2(n667), 
        .Q(\IDinst/n11294 ) );
  nnd2s1 \IDinst/U11374  ( .DIN1(\IDinst/n11271 ), .DIN2(n683), 
        .Q(\IDinst/n11293 ) );
  nnd2s1 \IDinst/U11373  ( .DIN1(\IDinst/n11291 ), .DIN2(\IDinst/n11290 ), 
        .Q(\IDinst/n11292 ) );
  nnd2s1 \IDinst/U11372  ( .DIN1(\IDinst/n11289 ), .DIN2(n1372), 
        .Q(\IDinst/n11291 ) );
  nnd2s1 \IDinst/U11371  ( .DIN1(\IDinst/n11280 ), .DIN2(n1371), 
        .Q(\IDinst/n11290 ) );
  nnd2s1 \IDinst/U11370  ( .DIN1(\IDinst/n11288 ), .DIN2(\IDinst/n11287 ), 
        .Q(\IDinst/n11289 ) );
  nnd2s1 \IDinst/U11369  ( .DIN1(\IDinst/n11286 ), .DIN2(n1318), 
        .Q(\IDinst/n11288 ) );
  nnd2s1 \IDinst/U11368  ( .DIN1(\IDinst/n11283 ), .DIN2(n1352), 
        .Q(\IDinst/n11287 ) );
  nnd2s1 \IDinst/U11367  ( .DIN1(\IDinst/n11285 ), .DIN2(\IDinst/n11284 ), 
        .Q(\IDinst/n11286 ) );
  nnd2s1 \IDinst/U11366  ( .DIN1(\IDinst/RegFile[31][25] ), .DIN2(n1215), 
        .Q(\IDinst/n11285 ) );
  nnd2s1 \IDinst/U11365  ( .DIN1(\IDinst/RegFile[30][25] ), .DIN2(n1271), 
        .Q(\IDinst/n11284 ) );
  nnd2s1 \IDinst/U11364  ( .DIN1(\IDinst/n11282 ), .DIN2(\IDinst/n11281 ), 
        .Q(\IDinst/n11283 ) );
  nnd2s1 \IDinst/U11363  ( .DIN1(\IDinst/RegFile[29][25] ), .DIN2(n1215), 
        .Q(\IDinst/n11282 ) );
  nnd2s1 \IDinst/U11362  ( .DIN1(\IDinst/RegFile[28][25] ), .DIN2(n1271), 
        .Q(\IDinst/n11281 ) );
  nnd2s1 \IDinst/U11361  ( .DIN1(\IDinst/n11279 ), .DIN2(\IDinst/n11278 ), 
        .Q(\IDinst/n11280 ) );
  nnd2s1 \IDinst/U11360  ( .DIN1(\IDinst/n11277 ), .DIN2(n1318), 
        .Q(\IDinst/n11279 ) );
  nnd2s1 \IDinst/U11359  ( .DIN1(\IDinst/n11274 ), .DIN2(n1352), 
        .Q(\IDinst/n11278 ) );
  nnd2s1 \IDinst/U11358  ( .DIN1(\IDinst/n11276 ), .DIN2(\IDinst/n11275 ), 
        .Q(\IDinst/n11277 ) );
  nnd2s1 \IDinst/U11357  ( .DIN1(\IDinst/RegFile[27][25] ), .DIN2(n1216), 
        .Q(\IDinst/n11276 ) );
  nnd2s1 \IDinst/U11356  ( .DIN1(\IDinst/RegFile[26][25] ), .DIN2(n1271), 
        .Q(\IDinst/n11275 ) );
  nnd2s1 \IDinst/U11355  ( .DIN1(\IDinst/n11273 ), .DIN2(\IDinst/n11272 ), 
        .Q(\IDinst/n11274 ) );
  nnd2s1 \IDinst/U11354  ( .DIN1(\IDinst/RegFile[25][25] ), .DIN2(n1216), 
        .Q(\IDinst/n11273 ) );
  nnd2s1 \IDinst/U11353  ( .DIN1(\IDinst/RegFile[24][25] ), .DIN2(n1271), 
        .Q(\IDinst/n11272 ) );
  nnd2s1 \IDinst/U11352  ( .DIN1(\IDinst/n11270 ), .DIN2(\IDinst/n11269 ), 
        .Q(\IDinst/n11271 ) );
  nnd2s1 \IDinst/U11351  ( .DIN1(\IDinst/n11268 ), .DIN2(n1380), 
        .Q(\IDinst/n11270 ) );
  nnd2s1 \IDinst/U11350  ( .DIN1(\IDinst/n11259 ), .DIN2(n1371), 
        .Q(\IDinst/n11269 ) );
  nnd2s1 \IDinst/U11349  ( .DIN1(\IDinst/n11267 ), .DIN2(\IDinst/n11266 ), 
        .Q(\IDinst/n11268 ) );
  nnd2s1 \IDinst/U11348  ( .DIN1(\IDinst/n11265 ), .DIN2(n1318), 
        .Q(\IDinst/n11267 ) );
  nnd2s1 \IDinst/U11347  ( .DIN1(\IDinst/n11262 ), .DIN2(n1352), 
        .Q(\IDinst/n11266 ) );
  nnd2s1 \IDinst/U11346  ( .DIN1(\IDinst/n11264 ), .DIN2(\IDinst/n11263 ), 
        .Q(\IDinst/n11265 ) );
  nnd2s1 \IDinst/U11345  ( .DIN1(\IDinst/RegFile[23][25] ), .DIN2(n1216), 
        .Q(\IDinst/n11264 ) );
  nnd2s1 \IDinst/U11344  ( .DIN1(\IDinst/RegFile[22][25] ), .DIN2(n1271), 
        .Q(\IDinst/n11263 ) );
  nnd2s1 \IDinst/U11343  ( .DIN1(\IDinst/n11261 ), .DIN2(\IDinst/n11260 ), 
        .Q(\IDinst/n11262 ) );
  nnd2s1 \IDinst/U11342  ( .DIN1(\IDinst/RegFile[21][25] ), .DIN2(n1216), 
        .Q(\IDinst/n11261 ) );
  nnd2s1 \IDinst/U11341  ( .DIN1(\IDinst/RegFile[20][25] ), .DIN2(n1271), 
        .Q(\IDinst/n11260 ) );
  nnd2s1 \IDinst/U11340  ( .DIN1(\IDinst/n11258 ), .DIN2(\IDinst/n11257 ), 
        .Q(\IDinst/n11259 ) );
  nnd2s1 \IDinst/U11339  ( .DIN1(\IDinst/n11256 ), .DIN2(n1318), 
        .Q(\IDinst/n11258 ) );
  nnd2s1 \IDinst/U11338  ( .DIN1(\IDinst/n11253 ), .DIN2(n1353), 
        .Q(\IDinst/n11257 ) );
  nnd2s1 \IDinst/U11337  ( .DIN1(\IDinst/n11255 ), .DIN2(\IDinst/n11254 ), 
        .Q(\IDinst/n11256 ) );
  nnd2s1 \IDinst/U11336  ( .DIN1(\IDinst/RegFile[19][25] ), .DIN2(n1216), 
        .Q(\IDinst/n11255 ) );
  nnd2s1 \IDinst/U11335  ( .DIN1(\IDinst/RegFile[18][25] ), .DIN2(n1271), 
        .Q(\IDinst/n11254 ) );
  nnd2s1 \IDinst/U11334  ( .DIN1(\IDinst/n11252 ), .DIN2(\IDinst/n11251 ), 
        .Q(\IDinst/n11253 ) );
  nnd2s1 \IDinst/U11333  ( .DIN1(\IDinst/RegFile[17][25] ), .DIN2(n1216), 
        .Q(\IDinst/n11252 ) );
  nnd2s1 \IDinst/U11332  ( .DIN1(\IDinst/RegFile[16][25] ), .DIN2(n1271), 
        .Q(\IDinst/n11251 ) );
  nnd2s1 \IDinst/U11331  ( .DIN1(\IDinst/n11249 ), .DIN2(\IDinst/n11248 ), 
        .Q(\IDinst/n11250 ) );
  nnd2s1 \IDinst/U11330  ( .DIN1(\IDinst/n11247 ), .DIN2(n665), 
        .Q(\IDinst/n11249 ) );
  nnd2s1 \IDinst/U11329  ( .DIN1(\IDinst/n11226 ), .DIN2(n682), 
        .Q(\IDinst/n11248 ) );
  nnd2s1 \IDinst/U11328  ( .DIN1(\IDinst/n11246 ), .DIN2(\IDinst/n11245 ), 
        .Q(\IDinst/n11247 ) );
  nnd2s1 \IDinst/U11327  ( .DIN1(\IDinst/n11244 ), .DIN2(n1379), 
        .Q(\IDinst/n11246 ) );
  nnd2s1 \IDinst/U11326  ( .DIN1(\IDinst/n11235 ), .DIN2(n1371), 
        .Q(\IDinst/n11245 ) );
  nnd2s1 \IDinst/U11325  ( .DIN1(\IDinst/n11243 ), .DIN2(\IDinst/n11242 ), 
        .Q(\IDinst/n11244 ) );
  nnd2s1 \IDinst/U11324  ( .DIN1(\IDinst/n11241 ), .DIN2(n1318), 
        .Q(\IDinst/n11243 ) );
  nnd2s1 \IDinst/U11323  ( .DIN1(\IDinst/n11238 ), .DIN2(n1353), 
        .Q(\IDinst/n11242 ) );
  nnd2s1 \IDinst/U11322  ( .DIN1(\IDinst/n11240 ), .DIN2(\IDinst/n11239 ), 
        .Q(\IDinst/n11241 ) );
  nnd2s1 \IDinst/U11321  ( .DIN1(\IDinst/RegFile[15][25] ), .DIN2(n1216), 
        .Q(\IDinst/n11240 ) );
  nnd2s1 \IDinst/U11320  ( .DIN1(\IDinst/RegFile[14][25] ), .DIN2(n1271), 
        .Q(\IDinst/n11239 ) );
  nnd2s1 \IDinst/U11319  ( .DIN1(\IDinst/n11237 ), .DIN2(\IDinst/n11236 ), 
        .Q(\IDinst/n11238 ) );
  nnd2s1 \IDinst/U11318  ( .DIN1(\IDinst/RegFile[13][25] ), .DIN2(n1216), 
        .Q(\IDinst/n11237 ) );
  nnd2s1 \IDinst/U11317  ( .DIN1(\IDinst/RegFile[12][25] ), .DIN2(n1270), 
        .Q(\IDinst/n11236 ) );
  nnd2s1 \IDinst/U11316  ( .DIN1(\IDinst/n11234 ), .DIN2(\IDinst/n11233 ), 
        .Q(\IDinst/n11235 ) );
  nnd2s1 \IDinst/U11315  ( .DIN1(\IDinst/n11232 ), .DIN2(n1318), 
        .Q(\IDinst/n11234 ) );
  nnd2s1 \IDinst/U11314  ( .DIN1(\IDinst/n11229 ), .DIN2(n1353), 
        .Q(\IDinst/n11233 ) );
  nnd2s1 \IDinst/U11313  ( .DIN1(\IDinst/n11231 ), .DIN2(\IDinst/n11230 ), 
        .Q(\IDinst/n11232 ) );
  nnd2s1 \IDinst/U11312  ( .DIN1(\IDinst/RegFile[11][25] ), .DIN2(n1216), 
        .Q(\IDinst/n11231 ) );
  nnd2s1 \IDinst/U11311  ( .DIN1(\IDinst/RegFile[10][25] ), .DIN2(n1270), 
        .Q(\IDinst/n11230 ) );
  nnd2s1 \IDinst/U11310  ( .DIN1(\IDinst/n11228 ), .DIN2(\IDinst/n11227 ), 
        .Q(\IDinst/n11229 ) );
  nnd2s1 \IDinst/U11309  ( .DIN1(\IDinst/RegFile[9][25] ), .DIN2(n1216), 
        .Q(\IDinst/n11228 ) );
  nnd2s1 \IDinst/U11308  ( .DIN1(\IDinst/RegFile[8][25] ), .DIN2(n1270), 
        .Q(\IDinst/n11227 ) );
  nnd2s1 \IDinst/U11307  ( .DIN1(\IDinst/n11225 ), .DIN2(\IDinst/n11224 ), 
        .Q(\IDinst/n11226 ) );
  nnd2s1 \IDinst/U11306  ( .DIN1(\IDinst/n11223 ), .DIN2(n1375), 
        .Q(\IDinst/n11225 ) );
  nnd2s1 \IDinst/U11305  ( .DIN1(\IDinst/n11214 ), .DIN2(n1371), 
        .Q(\IDinst/n11224 ) );
  nnd2s1 \IDinst/U11304  ( .DIN1(\IDinst/n11222 ), .DIN2(\IDinst/n11221 ), 
        .Q(\IDinst/n11223 ) );
  nnd2s1 \IDinst/U11303  ( .DIN1(\IDinst/n11220 ), .DIN2(n1318), 
        .Q(\IDinst/n11222 ) );
  nnd2s1 \IDinst/U11302  ( .DIN1(\IDinst/n11217 ), .DIN2(n1353), 
        .Q(\IDinst/n11221 ) );
  nnd2s1 \IDinst/U11301  ( .DIN1(\IDinst/n11219 ), .DIN2(\IDinst/n11218 ), 
        .Q(\IDinst/n11220 ) );
  nnd2s1 \IDinst/U11300  ( .DIN1(\IDinst/RegFile[7][25] ), .DIN2(n1216), 
        .Q(\IDinst/n11219 ) );
  nnd2s1 \IDinst/U11299  ( .DIN1(\IDinst/RegFile[6][25] ), .DIN2(n1270), 
        .Q(\IDinst/n11218 ) );
  nnd2s1 \IDinst/U11298  ( .DIN1(\IDinst/n11216 ), .DIN2(\IDinst/n11215 ), 
        .Q(\IDinst/n11217 ) );
  nnd2s1 \IDinst/U11297  ( .DIN1(\IDinst/RegFile[5][25] ), .DIN2(n1216), 
        .Q(\IDinst/n11216 ) );
  nnd2s1 \IDinst/U11296  ( .DIN1(\IDinst/RegFile[4][25] ), .DIN2(n1270), 
        .Q(\IDinst/n11215 ) );
  nnd2s1 \IDinst/U11295  ( .DIN1(\IDinst/n11213 ), .DIN2(\IDinst/n11212 ), 
        .Q(\IDinst/n11214 ) );
  nnd2s1 \IDinst/U11294  ( .DIN1(\IDinst/n11211 ), .DIN2(n1318), 
        .Q(\IDinst/n11213 ) );
  nnd2s1 \IDinst/U11293  ( .DIN1(\IDinst/n11208 ), .DIN2(n1353), 
        .Q(\IDinst/n11212 ) );
  nnd2s1 \IDinst/U11292  ( .DIN1(\IDinst/n11210 ), .DIN2(\IDinst/n11209 ), 
        .Q(\IDinst/n11211 ) );
  nnd2s1 \IDinst/U11291  ( .DIN1(\IDinst/RegFile[3][25] ), .DIN2(n1216), 
        .Q(\IDinst/n11210 ) );
  nnd2s1 \IDinst/U11290  ( .DIN1(\IDinst/RegFile[2][25] ), .DIN2(n1270), 
        .Q(\IDinst/n11209 ) );
  nnd2s1 \IDinst/U11289  ( .DIN1(\IDinst/n11207 ), .DIN2(\IDinst/n11206 ), 
        .Q(\IDinst/n11208 ) );
  nnd2s1 \IDinst/U11288  ( .DIN1(\IDinst/RegFile[1][25] ), .DIN2(n1217), 
        .Q(\IDinst/n11207 ) );
  nnd2s1 \IDinst/U11287  ( .DIN1(\IDinst/RegFile[0][25] ), .DIN2(n1270), 
        .Q(\IDinst/n11206 ) );
  nnd2s1 \IDinst/U11286  ( .DIN1(\IDinst/n11205 ), .DIN2(n535), 
        .Q(\IDinst/n8940 ) );
  nnd2s1 \IDinst/U11285  ( .DIN1(\IDinst/n11160 ), .DIN2(n634), 
        .Q(\IDinst/n8941 ) );
  nnd2s1 \IDinst/U11284  ( .DIN1(\IDinst/n11204 ), .DIN2(\IDinst/n11203 ), 
        .Q(\IDinst/n11205 ) );
  nnd2s1 \IDinst/U11283  ( .DIN1(\IDinst/n11202 ), .DIN2(n668), 
        .Q(\IDinst/n11204 ) );
  nnd2s1 \IDinst/U11282  ( .DIN1(\IDinst/n11181 ), .DIN2(n680), 
        .Q(\IDinst/n11203 ) );
  nnd2s1 \IDinst/U11281  ( .DIN1(\IDinst/n11201 ), .DIN2(\IDinst/n11200 ), 
        .Q(\IDinst/n11202 ) );
  nnd2s1 \IDinst/U11280  ( .DIN1(\IDinst/n11199 ), .DIN2(n1374), 
        .Q(\IDinst/n11201 ) );
  nnd2s1 \IDinst/U11279  ( .DIN1(\IDinst/n11190 ), .DIN2(n1371), 
        .Q(\IDinst/n11200 ) );
  nnd2s1 \IDinst/U11278  ( .DIN1(\IDinst/n11198 ), .DIN2(\IDinst/n11197 ), 
        .Q(\IDinst/n11199 ) );
  nnd2s1 \IDinst/U11277  ( .DIN1(\IDinst/n11196 ), .DIN2(n1318), 
        .Q(\IDinst/n11198 ) );
  nnd2s1 \IDinst/U11276  ( .DIN1(\IDinst/n11193 ), .DIN2(n1353), 
        .Q(\IDinst/n11197 ) );
  nnd2s1 \IDinst/U11275  ( .DIN1(\IDinst/n11195 ), .DIN2(\IDinst/n11194 ), 
        .Q(\IDinst/n11196 ) );
  nnd2s1 \IDinst/U11274  ( .DIN1(\IDinst/RegFile[31][24] ), .DIN2(n1217), 
        .Q(\IDinst/n11195 ) );
  nnd2s1 \IDinst/U11273  ( .DIN1(\IDinst/RegFile[30][24] ), .DIN2(n1270), 
        .Q(\IDinst/n11194 ) );
  nnd2s1 \IDinst/U11272  ( .DIN1(\IDinst/n11192 ), .DIN2(\IDinst/n11191 ), 
        .Q(\IDinst/n11193 ) );
  nnd2s1 \IDinst/U11271  ( .DIN1(\IDinst/RegFile[29][24] ), .DIN2(n1217), 
        .Q(\IDinst/n11192 ) );
  nnd2s1 \IDinst/U11270  ( .DIN1(\IDinst/RegFile[28][24] ), .DIN2(n1270), 
        .Q(\IDinst/n11191 ) );
  nnd2s1 \IDinst/U11269  ( .DIN1(\IDinst/n11189 ), .DIN2(\IDinst/n11188 ), 
        .Q(\IDinst/n11190 ) );
  nnd2s1 \IDinst/U11268  ( .DIN1(\IDinst/n11187 ), .DIN2(n1318), 
        .Q(\IDinst/n11189 ) );
  nnd2s1 \IDinst/U11267  ( .DIN1(\IDinst/n11184 ), .DIN2(n1353), 
        .Q(\IDinst/n11188 ) );
  nnd2s1 \IDinst/U11266  ( .DIN1(\IDinst/n11186 ), .DIN2(\IDinst/n11185 ), 
        .Q(\IDinst/n11187 ) );
  nnd2s1 \IDinst/U11265  ( .DIN1(\IDinst/RegFile[27][24] ), .DIN2(n1217), 
        .Q(\IDinst/n11186 ) );
  nnd2s1 \IDinst/U11264  ( .DIN1(\IDinst/RegFile[26][24] ), .DIN2(n1269), 
        .Q(\IDinst/n11185 ) );
  nnd2s1 \IDinst/U11263  ( .DIN1(\IDinst/n11183 ), .DIN2(\IDinst/n11182 ), 
        .Q(\IDinst/n11184 ) );
  nnd2s1 \IDinst/U11262  ( .DIN1(\IDinst/RegFile[25][24] ), .DIN2(n1217), 
        .Q(\IDinst/n11183 ) );
  nnd2s1 \IDinst/U11261  ( .DIN1(\IDinst/RegFile[24][24] ), .DIN2(n1269), 
        .Q(\IDinst/n11182 ) );
  nnd2s1 \IDinst/U11260  ( .DIN1(\IDinst/n11180 ), .DIN2(\IDinst/n11179 ), 
        .Q(\IDinst/n11181 ) );
  nnd2s1 \IDinst/U11259  ( .DIN1(\IDinst/n11178 ), .DIN2(\IDinst/N46 ), 
        .Q(\IDinst/n11180 ) );
  nnd2s1 \IDinst/U11258  ( .DIN1(\IDinst/n11169 ), .DIN2(n1371), 
        .Q(\IDinst/n11179 ) );
  nnd2s1 \IDinst/U11257  ( .DIN1(\IDinst/n11177 ), .DIN2(\IDinst/n11176 ), 
        .Q(\IDinst/n11178 ) );
  nnd2s1 \IDinst/U11256  ( .DIN1(\IDinst/n11175 ), .DIN2(n1318), 
        .Q(\IDinst/n11177 ) );
  nnd2s1 \IDinst/U11255  ( .DIN1(\IDinst/n11172 ), .DIN2(n1353), 
        .Q(\IDinst/n11176 ) );
  nnd2s1 \IDinst/U11254  ( .DIN1(\IDinst/n11174 ), .DIN2(\IDinst/n11173 ), 
        .Q(\IDinst/n11175 ) );
  nnd2s1 \IDinst/U11253  ( .DIN1(\IDinst/RegFile[23][24] ), .DIN2(n1217), 
        .Q(\IDinst/n11174 ) );
  nnd2s1 \IDinst/U11252  ( .DIN1(\IDinst/RegFile[22][24] ), .DIN2(n1269), 
        .Q(\IDinst/n11173 ) );
  nnd2s1 \IDinst/U11251  ( .DIN1(\IDinst/n11171 ), .DIN2(\IDinst/n11170 ), 
        .Q(\IDinst/n11172 ) );
  nnd2s1 \IDinst/U11250  ( .DIN1(\IDinst/RegFile[21][24] ), .DIN2(n1217), 
        .Q(\IDinst/n11171 ) );
  nnd2s1 \IDinst/U11249  ( .DIN1(\IDinst/RegFile[20][24] ), .DIN2(n1276), 
        .Q(\IDinst/n11170 ) );
  nnd2s1 \IDinst/U11248  ( .DIN1(\IDinst/n11168 ), .DIN2(\IDinst/n11167 ), 
        .Q(\IDinst/n11169 ) );
  nnd2s1 \IDinst/U11247  ( .DIN1(\IDinst/n11166 ), .DIN2(n1317), 
        .Q(\IDinst/n11168 ) );
  nnd2s1 \IDinst/U11246  ( .DIN1(\IDinst/n11163 ), .DIN2(n1354), 
        .Q(\IDinst/n11167 ) );
  nnd2s1 \IDinst/U11245  ( .DIN1(\IDinst/n11165 ), .DIN2(\IDinst/n11164 ), 
        .Q(\IDinst/n11166 ) );
  nnd2s1 \IDinst/U11244  ( .DIN1(\IDinst/RegFile[19][24] ), .DIN2(n1217), 
        .Q(\IDinst/n11165 ) );
  nnd2s1 \IDinst/U11243  ( .DIN1(\IDinst/RegFile[18][24] ), .DIN2(n1289), 
        .Q(\IDinst/n11164 ) );
  nnd2s1 \IDinst/U11242  ( .DIN1(\IDinst/n11162 ), .DIN2(\IDinst/n11161 ), 
        .Q(\IDinst/n11163 ) );
  nnd2s1 \IDinst/U11241  ( .DIN1(\IDinst/RegFile[17][24] ), .DIN2(n1217), 
        .Q(\IDinst/n11162 ) );
  nnd2s1 \IDinst/U11240  ( .DIN1(\IDinst/RegFile[16][24] ), .DIN2(n1289), 
        .Q(\IDinst/n11161 ) );
  nnd2s1 \IDinst/U11239  ( .DIN1(\IDinst/n11159 ), .DIN2(\IDinst/n11158 ), 
        .Q(\IDinst/n11160 ) );
  nnd2s1 \IDinst/U11238  ( .DIN1(\IDinst/n11157 ), .DIN2(n666), 
        .Q(\IDinst/n11159 ) );
  nnd2s1 \IDinst/U11237  ( .DIN1(\IDinst/n11136 ), .DIN2(n681), 
        .Q(\IDinst/n11158 ) );
  nnd2s1 \IDinst/U11236  ( .DIN1(\IDinst/n11156 ), .DIN2(\IDinst/n11155 ), 
        .Q(\IDinst/n11157 ) );
  nnd2s1 \IDinst/U11235  ( .DIN1(\IDinst/n11154 ), .DIN2(n1372), 
        .Q(\IDinst/n11156 ) );
  nnd2s1 \IDinst/U11234  ( .DIN1(\IDinst/n11145 ), .DIN2(n1371), 
        .Q(\IDinst/n11155 ) );
  nnd2s1 \IDinst/U11233  ( .DIN1(\IDinst/n11153 ), .DIN2(\IDinst/n11152 ), 
        .Q(\IDinst/n11154 ) );
  nnd2s1 \IDinst/U11232  ( .DIN1(\IDinst/n11151 ), .DIN2(n1317), 
        .Q(\IDinst/n11153 ) );
  nnd2s1 \IDinst/U11231  ( .DIN1(\IDinst/n11148 ), .DIN2(n1354), 
        .Q(\IDinst/n11152 ) );
  nnd2s1 \IDinst/U11230  ( .DIN1(\IDinst/n11150 ), .DIN2(\IDinst/n11149 ), 
        .Q(\IDinst/n11151 ) );
  nnd2s1 \IDinst/U11229  ( .DIN1(\IDinst/RegFile[15][24] ), .DIN2(n1217), 
        .Q(\IDinst/n11150 ) );
  nnd2s1 \IDinst/U11228  ( .DIN1(\IDinst/RegFile[14][24] ), .DIN2(n1289), 
        .Q(\IDinst/n11149 ) );
  nnd2s1 \IDinst/U11227  ( .DIN1(\IDinst/n11147 ), .DIN2(\IDinst/n11146 ), 
        .Q(\IDinst/n11148 ) );
  nnd2s1 \IDinst/U11226  ( .DIN1(\IDinst/RegFile[13][24] ), .DIN2(n1217), 
        .Q(\IDinst/n11147 ) );
  nnd2s1 \IDinst/U11225  ( .DIN1(\IDinst/RegFile[12][24] ), .DIN2(n1289), 
        .Q(\IDinst/n11146 ) );
  nnd2s1 \IDinst/U11224  ( .DIN1(\IDinst/n11144 ), .DIN2(\IDinst/n11143 ), 
        .Q(\IDinst/n11145 ) );
  nnd2s1 \IDinst/U11223  ( .DIN1(\IDinst/n11142 ), .DIN2(n1317), 
        .Q(\IDinst/n11144 ) );
  nnd2s1 \IDinst/U11222  ( .DIN1(\IDinst/n11139 ), .DIN2(n1354), 
        .Q(\IDinst/n11143 ) );
  nnd2s1 \IDinst/U11221  ( .DIN1(\IDinst/n11141 ), .DIN2(\IDinst/n11140 ), 
        .Q(\IDinst/n11142 ) );
  nnd2s1 \IDinst/U11220  ( .DIN1(\IDinst/RegFile[11][24] ), .DIN2(n1217), 
        .Q(\IDinst/n11141 ) );
  nnd2s1 \IDinst/U11219  ( .DIN1(\IDinst/RegFile[10][24] ), .DIN2(n1289), 
        .Q(\IDinst/n11140 ) );
  nnd2s1 \IDinst/U11218  ( .DIN1(\IDinst/n11138 ), .DIN2(\IDinst/n11137 ), 
        .Q(\IDinst/n11139 ) );
  nnd2s1 \IDinst/U11217  ( .DIN1(\IDinst/RegFile[9][24] ), .DIN2(n1217), 
        .Q(\IDinst/n11138 ) );
  nnd2s1 \IDinst/U11216  ( .DIN1(\IDinst/RegFile[8][24] ), .DIN2(n1289), 
        .Q(\IDinst/n11137 ) );
  nnd2s1 \IDinst/U11215  ( .DIN1(\IDinst/n11135 ), .DIN2(\IDinst/n11134 ), 
        .Q(\IDinst/n11136 ) );
  nnd2s1 \IDinst/U11214  ( .DIN1(\IDinst/n11133 ), .DIN2(n1379), 
        .Q(\IDinst/n11135 ) );
  nnd2s1 \IDinst/U11213  ( .DIN1(\IDinst/n11124 ), .DIN2(n1371), 
        .Q(\IDinst/n11134 ) );
  nnd2s1 \IDinst/U11212  ( .DIN1(\IDinst/n11132 ), .DIN2(\IDinst/n11131 ), 
        .Q(\IDinst/n11133 ) );
  nnd2s1 \IDinst/U11211  ( .DIN1(\IDinst/n11130 ), .DIN2(n1317), 
        .Q(\IDinst/n11132 ) );
  nnd2s1 \IDinst/U11210  ( .DIN1(\IDinst/n11127 ), .DIN2(n1354), 
        .Q(\IDinst/n11131 ) );
  nnd2s1 \IDinst/U11209  ( .DIN1(\IDinst/n11129 ), .DIN2(\IDinst/n11128 ), 
        .Q(\IDinst/n11130 ) );
  nnd2s1 \IDinst/U11208  ( .DIN1(\IDinst/RegFile[7][24] ), .DIN2(n1218), 
        .Q(\IDinst/n11129 ) );
  nnd2s1 \IDinst/U11207  ( .DIN1(\IDinst/RegFile[6][24] ), .DIN2(n1289), 
        .Q(\IDinst/n11128 ) );
  nnd2s1 \IDinst/U11206  ( .DIN1(\IDinst/n11126 ), .DIN2(\IDinst/n11125 ), 
        .Q(\IDinst/n11127 ) );
  nnd2s1 \IDinst/U11205  ( .DIN1(\IDinst/RegFile[5][24] ), .DIN2(n1218), 
        .Q(\IDinst/n11126 ) );
  nnd2s1 \IDinst/U11204  ( .DIN1(\IDinst/RegFile[4][24] ), .DIN2(n1290), 
        .Q(\IDinst/n11125 ) );
  nnd2s1 \IDinst/U11203  ( .DIN1(\IDinst/n11123 ), .DIN2(\IDinst/n11122 ), 
        .Q(\IDinst/n11124 ) );
  nnd2s1 \IDinst/U11202  ( .DIN1(\IDinst/n11121 ), .DIN2(n1317), 
        .Q(\IDinst/n11123 ) );
  nnd2s1 \IDinst/U11201  ( .DIN1(\IDinst/n11118 ), .DIN2(n1354), 
        .Q(\IDinst/n11122 ) );
  nnd2s1 \IDinst/U11200  ( .DIN1(\IDinst/n11120 ), .DIN2(\IDinst/n11119 ), 
        .Q(\IDinst/n11121 ) );
  nnd2s1 \IDinst/U11199  ( .DIN1(\IDinst/RegFile[3][24] ), .DIN2(n1218), 
        .Q(\IDinst/n11120 ) );
  nnd2s1 \IDinst/U11198  ( .DIN1(\IDinst/RegFile[2][24] ), .DIN2(n1290), 
        .Q(\IDinst/n11119 ) );
  nnd2s1 \IDinst/U11197  ( .DIN1(\IDinst/n11117 ), .DIN2(\IDinst/n11116 ), 
        .Q(\IDinst/n11118 ) );
  nnd2s1 \IDinst/U11196  ( .DIN1(\IDinst/RegFile[1][24] ), .DIN2(n1218), 
        .Q(\IDinst/n11117 ) );
  nnd2s1 \IDinst/U11195  ( .DIN1(\IDinst/RegFile[0][24] ), .DIN2(n1290), 
        .Q(\IDinst/n11116 ) );
  nnd2s1 \IDinst/U11194  ( .DIN1(\IDinst/n11115 ), .DIN2(n534), 
        .Q(\IDinst/n8938 ) );
  nnd2s1 \IDinst/U11193  ( .DIN1(\IDinst/n11070 ), .DIN2(n533), 
        .Q(\IDinst/n8939 ) );
  nnd2s1 \IDinst/U11192  ( .DIN1(\IDinst/n11114 ), .DIN2(\IDinst/n11113 ), 
        .Q(\IDinst/n11115 ) );
  nnd2s1 \IDinst/U11191  ( .DIN1(\IDinst/n11112 ), .DIN2(n667), 
        .Q(\IDinst/n11114 ) );
  nnd2s1 \IDinst/U11190  ( .DIN1(\IDinst/n11091 ), .DIN2(n683), 
        .Q(\IDinst/n11113 ) );
  nnd2s1 \IDinst/U11189  ( .DIN1(\IDinst/n11111 ), .DIN2(\IDinst/n11110 ), 
        .Q(\IDinst/n11112 ) );
  nnd2s1 \IDinst/U11188  ( .DIN1(\IDinst/n11109 ), .DIN2(n1375), 
        .Q(\IDinst/n11111 ) );
  nnd2s1 \IDinst/U11187  ( .DIN1(\IDinst/n11100 ), .DIN2(n1371), 
        .Q(\IDinst/n11110 ) );
  nnd2s1 \IDinst/U11186  ( .DIN1(\IDinst/n11108 ), .DIN2(\IDinst/n11107 ), 
        .Q(\IDinst/n11109 ) );
  nnd2s1 \IDinst/U11185  ( .DIN1(\IDinst/n11106 ), .DIN2(n1317), 
        .Q(\IDinst/n11108 ) );
  nnd2s1 \IDinst/U11184  ( .DIN1(\IDinst/n11103 ), .DIN2(n1354), 
        .Q(\IDinst/n11107 ) );
  nnd2s1 \IDinst/U11183  ( .DIN1(\IDinst/n11105 ), .DIN2(\IDinst/n11104 ), 
        .Q(\IDinst/n11106 ) );
  nnd2s1 \IDinst/U11182  ( .DIN1(\IDinst/RegFile[31][23] ), .DIN2(n1203), 
        .Q(\IDinst/n11105 ) );
  nnd2s1 \IDinst/U11181  ( .DIN1(\IDinst/RegFile[30][23] ), .DIN2(n1290), 
        .Q(\IDinst/n11104 ) );
  nnd2s1 \IDinst/U11180  ( .DIN1(\IDinst/n11102 ), .DIN2(\IDinst/n11101 ), 
        .Q(\IDinst/n11103 ) );
  nnd2s1 \IDinst/U11179  ( .DIN1(\IDinst/RegFile[29][23] ), .DIN2(n1198), 
        .Q(\IDinst/n11102 ) );
  nnd2s1 \IDinst/U11178  ( .DIN1(\IDinst/RegFile[28][23] ), .DIN2(n1290), 
        .Q(\IDinst/n11101 ) );
  nnd2s1 \IDinst/U11177  ( .DIN1(\IDinst/n11099 ), .DIN2(\IDinst/n11098 ), 
        .Q(\IDinst/n11100 ) );
  nnd2s1 \IDinst/U11176  ( .DIN1(\IDinst/n11097 ), .DIN2(n1317), 
        .Q(\IDinst/n11099 ) );
  nnd2s1 \IDinst/U11175  ( .DIN1(\IDinst/n11094 ), .DIN2(n1354), 
        .Q(\IDinst/n11098 ) );
  nnd2s1 \IDinst/U11174  ( .DIN1(\IDinst/n11096 ), .DIN2(\IDinst/n11095 ), 
        .Q(\IDinst/n11097 ) );
  nnd2s1 \IDinst/U11173  ( .DIN1(\IDinst/RegFile[27][23] ), .DIN2(n1198), 
        .Q(\IDinst/n11096 ) );
  nnd2s1 \IDinst/U11172  ( .DIN1(\IDinst/RegFile[26][23] ), .DIN2(n1290), 
        .Q(\IDinst/n11095 ) );
  nnd2s1 \IDinst/U11171  ( .DIN1(\IDinst/n11093 ), .DIN2(\IDinst/n11092 ), 
        .Q(\IDinst/n11094 ) );
  nnd2s1 \IDinst/U11170  ( .DIN1(\IDinst/RegFile[25][23] ), .DIN2(n1198), 
        .Q(\IDinst/n11093 ) );
  nnd2s1 \IDinst/U11169  ( .DIN1(\IDinst/RegFile[24][23] ), .DIN2(n1290), 
        .Q(\IDinst/n11092 ) );
  nnd2s1 \IDinst/U11168  ( .DIN1(\IDinst/n11090 ), .DIN2(\IDinst/n11089 ), 
        .Q(\IDinst/n11091 ) );
  nnd2s1 \IDinst/U11167  ( .DIN1(\IDinst/n11088 ), .DIN2(n1373), 
        .Q(\IDinst/n11090 ) );
  nnd2s1 \IDinst/U11166  ( .DIN1(\IDinst/n11079 ), .DIN2(n1371), 
        .Q(\IDinst/n11089 ) );
  nnd2s1 \IDinst/U11165  ( .DIN1(\IDinst/n11087 ), .DIN2(\IDinst/n11086 ), 
        .Q(\IDinst/n11088 ) );
  nnd2s1 \IDinst/U11164  ( .DIN1(\IDinst/n11085 ), .DIN2(n1317), 
        .Q(\IDinst/n11087 ) );
  nnd2s1 \IDinst/U11163  ( .DIN1(\IDinst/n11082 ), .DIN2(n1354), 
        .Q(\IDinst/n11086 ) );
  nnd2s1 \IDinst/U11162  ( .DIN1(\IDinst/n11084 ), .DIN2(\IDinst/n11083 ), 
        .Q(\IDinst/n11085 ) );
  nnd2s1 \IDinst/U11161  ( .DIN1(\IDinst/RegFile[23][23] ), .DIN2(n1198), 
        .Q(\IDinst/n11084 ) );
  nnd2s1 \IDinst/U11160  ( .DIN1(\IDinst/RegFile[22][23] ), .DIN2(n1290), 
        .Q(\IDinst/n11083 ) );
  nnd2s1 \IDinst/U11159  ( .DIN1(\IDinst/n11081 ), .DIN2(\IDinst/n11080 ), 
        .Q(\IDinst/n11082 ) );
  nnd2s1 \IDinst/U11158  ( .DIN1(\IDinst/RegFile[21][23] ), .DIN2(n1199), 
        .Q(\IDinst/n11081 ) );
  nnd2s1 \IDinst/U11157  ( .DIN1(\IDinst/RegFile[20][23] ), .DIN2(n1290), 
        .Q(\IDinst/n11080 ) );
  nnd2s1 \IDinst/U11156  ( .DIN1(\IDinst/n11078 ), .DIN2(\IDinst/n11077 ), 
        .Q(\IDinst/n11079 ) );
  nnd2s1 \IDinst/U11155  ( .DIN1(\IDinst/n11076 ), .DIN2(n1317), 
        .Q(\IDinst/n11078 ) );
  nnd2s1 \IDinst/U11154  ( .DIN1(\IDinst/n11073 ), .DIN2(n1354), 
        .Q(\IDinst/n11077 ) );
  nnd2s1 \IDinst/U11153  ( .DIN1(\IDinst/n11075 ), .DIN2(\IDinst/n11074 ), 
        .Q(\IDinst/n11076 ) );
  nnd2s1 \IDinst/U11152  ( .DIN1(\IDinst/RegFile[19][23] ), .DIN2(n1199), 
        .Q(\IDinst/n11075 ) );
  nnd2s1 \IDinst/U11151  ( .DIN1(\IDinst/RegFile[18][23] ), .DIN2(n1291), 
        .Q(\IDinst/n11074 ) );
  nnd2s1 \IDinst/U11150  ( .DIN1(\IDinst/n11072 ), .DIN2(\IDinst/n11071 ), 
        .Q(\IDinst/n11073 ) );
  nnd2s1 \IDinst/U11149  ( .DIN1(\IDinst/RegFile[17][23] ), .DIN2(n1199), 
        .Q(\IDinst/n11072 ) );
  nnd2s1 \IDinst/U11148  ( .DIN1(\IDinst/RegFile[16][23] ), .DIN2(n1291), 
        .Q(\IDinst/n11071 ) );
  nnd2s1 \IDinst/U11147  ( .DIN1(\IDinst/n11069 ), .DIN2(\IDinst/n11068 ), 
        .Q(\IDinst/n11070 ) );
  nnd2s1 \IDinst/U11146  ( .DIN1(\IDinst/n11067 ), .DIN2(n665), 
        .Q(\IDinst/n11069 ) );
  nnd2s1 \IDinst/U11145  ( .DIN1(\IDinst/n11046 ), .DIN2(n682), 
        .Q(\IDinst/n11068 ) );
  nnd2s1 \IDinst/U11144  ( .DIN1(\IDinst/n11066 ), .DIN2(\IDinst/n11065 ), 
        .Q(\IDinst/n11067 ) );
  nnd2s1 \IDinst/U11143  ( .DIN1(\IDinst/n11064 ), .DIN2(n1376), 
        .Q(\IDinst/n11066 ) );
  nnd2s1 \IDinst/U11142  ( .DIN1(\IDinst/n11055 ), .DIN2(n1370), 
        .Q(\IDinst/n11065 ) );
  nnd2s1 \IDinst/U11141  ( .DIN1(\IDinst/n11063 ), .DIN2(\IDinst/n11062 ), 
        .Q(\IDinst/n11064 ) );
  nnd2s1 \IDinst/U11140  ( .DIN1(\IDinst/n11061 ), .DIN2(n1317), 
        .Q(\IDinst/n11063 ) );
  nnd2s1 \IDinst/U11139  ( .DIN1(\IDinst/n11058 ), .DIN2(n1355), 
        .Q(\IDinst/n11062 ) );
  nnd2s1 \IDinst/U11138  ( .DIN1(\IDinst/n11060 ), .DIN2(\IDinst/n11059 ), 
        .Q(\IDinst/n11061 ) );
  nnd2s1 \IDinst/U11137  ( .DIN1(\IDinst/RegFile[15][23] ), .DIN2(n1199), 
        .Q(\IDinst/n11060 ) );
  nnd2s1 \IDinst/U11136  ( .DIN1(\IDinst/RegFile[14][23] ), .DIN2(n1291), 
        .Q(\IDinst/n11059 ) );
  nnd2s1 \IDinst/U11135  ( .DIN1(\IDinst/n11057 ), .DIN2(\IDinst/n11056 ), 
        .Q(\IDinst/n11058 ) );
  nnd2s1 \IDinst/U11134  ( .DIN1(\IDinst/RegFile[13][23] ), .DIN2(n1199), 
        .Q(\IDinst/n11057 ) );
  nnd2s1 \IDinst/U11133  ( .DIN1(\IDinst/RegFile[12][23] ), .DIN2(n1291), 
        .Q(\IDinst/n11056 ) );
  nnd2s1 \IDinst/U11132  ( .DIN1(\IDinst/n11054 ), .DIN2(\IDinst/n11053 ), 
        .Q(\IDinst/n11055 ) );
  nnd2s1 \IDinst/U11131  ( .DIN1(\IDinst/n11052 ), .DIN2(n1317), 
        .Q(\IDinst/n11054 ) );
  nnd2s1 \IDinst/U11130  ( .DIN1(\IDinst/n11049 ), .DIN2(n1355), 
        .Q(\IDinst/n11053 ) );
  nnd2s1 \IDinst/U11129  ( .DIN1(\IDinst/n11051 ), .DIN2(\IDinst/n11050 ), 
        .Q(\IDinst/n11052 ) );
  nnd2s1 \IDinst/U11128  ( .DIN1(\IDinst/RegFile[11][23] ), .DIN2(n1199), 
        .Q(\IDinst/n11051 ) );
  nnd2s1 \IDinst/U11127  ( .DIN1(\IDinst/RegFile[10][23] ), .DIN2(n1291), 
        .Q(\IDinst/n11050 ) );
  nnd2s1 \IDinst/U11126  ( .DIN1(\IDinst/n11048 ), .DIN2(\IDinst/n11047 ), 
        .Q(\IDinst/n11049 ) );
  nnd2s1 \IDinst/U11125  ( .DIN1(\IDinst/RegFile[9][23] ), .DIN2(n1199), 
        .Q(\IDinst/n11048 ) );
  nnd2s1 \IDinst/U11124  ( .DIN1(\IDinst/RegFile[8][23] ), .DIN2(n1291), 
        .Q(\IDinst/n11047 ) );
  nnd2s1 \IDinst/U11123  ( .DIN1(\IDinst/n11045 ), .DIN2(\IDinst/n11044 ), 
        .Q(\IDinst/n11046 ) );
  nnd2s1 \IDinst/U11122  ( .DIN1(\IDinst/n11043 ), .DIN2(n1377), 
        .Q(\IDinst/n11045 ) );
  nnd2s1 \IDinst/U11121  ( .DIN1(\IDinst/n11034 ), .DIN2(n1370), 
        .Q(\IDinst/n11044 ) );
  nnd2s1 \IDinst/U11120  ( .DIN1(\IDinst/n11042 ), .DIN2(\IDinst/n11041 ), 
        .Q(\IDinst/n11043 ) );
  nnd2s1 \IDinst/U11119  ( .DIN1(\IDinst/n11040 ), .DIN2(n1317), 
        .Q(\IDinst/n11042 ) );
  nnd2s1 \IDinst/U11118  ( .DIN1(\IDinst/n11037 ), .DIN2(n1355), 
        .Q(\IDinst/n11041 ) );
  nnd2s1 \IDinst/U11117  ( .DIN1(\IDinst/n11039 ), .DIN2(\IDinst/n11038 ), 
        .Q(\IDinst/n11040 ) );
  nnd2s1 \IDinst/U11116  ( .DIN1(\IDinst/RegFile[7][23] ), .DIN2(n1199), 
        .Q(\IDinst/n11039 ) );
  nnd2s1 \IDinst/U11115  ( .DIN1(\IDinst/RegFile[6][23] ), .DIN2(n1291), 
        .Q(\IDinst/n11038 ) );
  nnd2s1 \IDinst/U11114  ( .DIN1(\IDinst/n11036 ), .DIN2(\IDinst/n11035 ), 
        .Q(\IDinst/n11037 ) );
  nnd2s1 \IDinst/U11113  ( .DIN1(\IDinst/RegFile[5][23] ), .DIN2(n1199), 
        .Q(\IDinst/n11036 ) );
  nnd2s1 \IDinst/U11112  ( .DIN1(\IDinst/RegFile[4][23] ), .DIN2(n1291), 
        .Q(\IDinst/n11035 ) );
  nnd2s1 \IDinst/U11111  ( .DIN1(\IDinst/n11033 ), .DIN2(\IDinst/n11032 ), 
        .Q(\IDinst/n11034 ) );
  nnd2s1 \IDinst/U11110  ( .DIN1(\IDinst/n11031 ), .DIN2(n1316), 
        .Q(\IDinst/n11033 ) );
  nnd2s1 \IDinst/U11109  ( .DIN1(\IDinst/n11028 ), .DIN2(n1355), 
        .Q(\IDinst/n11032 ) );
  nnd2s1 \IDinst/U11108  ( .DIN1(\IDinst/n11030 ), .DIN2(\IDinst/n11029 ), 
        .Q(\IDinst/n11031 ) );
  nnd2s1 \IDinst/U11107  ( .DIN1(\IDinst/RegFile[3][23] ), .DIN2(n1199), 
        .Q(\IDinst/n11030 ) );
  nnd2s1 \IDinst/U11106  ( .DIN1(\IDinst/RegFile[2][23] ), .DIN2(n1291), 
        .Q(\IDinst/n11029 ) );
  nnd2s1 \IDinst/U11105  ( .DIN1(\IDinst/n11027 ), .DIN2(\IDinst/n11026 ), 
        .Q(\IDinst/n11028 ) );
  nnd2s1 \IDinst/U11104  ( .DIN1(\IDinst/RegFile[1][23] ), .DIN2(n1199), 
        .Q(\IDinst/n11027 ) );
  nnd2s1 \IDinst/U11103  ( .DIN1(\IDinst/RegFile[0][23] ), .DIN2(n1292), 
        .Q(\IDinst/n11026 ) );
  nnd2s1 \IDinst/U11102  ( .DIN1(\IDinst/n11025 ), .DIN2(\IDinst/N48 ), 
        .Q(\IDinst/n8936 ) );
  nnd2s1 \IDinst/U11101  ( .DIN1(\IDinst/n10980 ), .DIN2(n634), 
        .Q(\IDinst/n8937 ) );
  nnd2s1 \IDinst/U11100  ( .DIN1(\IDinst/n11024 ), .DIN2(\IDinst/n11023 ), 
        .Q(\IDinst/n11025 ) );
  nnd2s1 \IDinst/U11099  ( .DIN1(\IDinst/n11022 ), .DIN2(n668), 
        .Q(\IDinst/n11024 ) );
  nnd2s1 \IDinst/U11098  ( .DIN1(\IDinst/n11001 ), .DIN2(n680), 
        .Q(\IDinst/n11023 ) );
  nnd2s1 \IDinst/U11097  ( .DIN1(\IDinst/n11021 ), .DIN2(\IDinst/n11020 ), 
        .Q(\IDinst/n11022 ) );
  nnd2s1 \IDinst/U11096  ( .DIN1(\IDinst/n11019 ), .DIN2(n1374), 
        .Q(\IDinst/n11021 ) );
  nnd2s1 \IDinst/U11095  ( .DIN1(\IDinst/n11010 ), .DIN2(n1370), 
        .Q(\IDinst/n11020 ) );
  nnd2s1 \IDinst/U11094  ( .DIN1(\IDinst/n11018 ), .DIN2(\IDinst/n11017 ), 
        .Q(\IDinst/n11019 ) );
  nnd2s1 \IDinst/U11093  ( .DIN1(\IDinst/n11016 ), .DIN2(n1316), 
        .Q(\IDinst/n11018 ) );
  nnd2s1 \IDinst/U11092  ( .DIN1(\IDinst/n11013 ), .DIN2(n1355), 
        .Q(\IDinst/n11017 ) );
  nnd2s1 \IDinst/U11091  ( .DIN1(\IDinst/n11015 ), .DIN2(\IDinst/n11014 ), 
        .Q(\IDinst/n11016 ) );
  nnd2s1 \IDinst/U11090  ( .DIN1(\IDinst/RegFile[31][22] ), .DIN2(n1199), 
        .Q(\IDinst/n11015 ) );
  nnd2s1 \IDinst/U11089  ( .DIN1(\IDinst/RegFile[30][22] ), .DIN2(n1292), 
        .Q(\IDinst/n11014 ) );
  nnd2s1 \IDinst/U11088  ( .DIN1(\IDinst/n11012 ), .DIN2(\IDinst/n11011 ), 
        .Q(\IDinst/n11013 ) );
  nnd2s1 \IDinst/U11087  ( .DIN1(\IDinst/RegFile[29][22] ), .DIN2(n1199), 
        .Q(\IDinst/n11012 ) );
  nnd2s1 \IDinst/U11086  ( .DIN1(\IDinst/RegFile[28][22] ), .DIN2(n1292), 
        .Q(\IDinst/n11011 ) );
  nnd2s1 \IDinst/U11085  ( .DIN1(\IDinst/n11009 ), .DIN2(\IDinst/n11008 ), 
        .Q(\IDinst/n11010 ) );
  nnd2s1 \IDinst/U11084  ( .DIN1(\IDinst/n11007 ), .DIN2(n1316), 
        .Q(\IDinst/n11009 ) );
  nnd2s1 \IDinst/U11083  ( .DIN1(\IDinst/n11004 ), .DIN2(n1355), 
        .Q(\IDinst/n11008 ) );
  nnd2s1 \IDinst/U11082  ( .DIN1(\IDinst/n11006 ), .DIN2(\IDinst/n11005 ), 
        .Q(\IDinst/n11007 ) );
  nnd2s1 \IDinst/U11081  ( .DIN1(\IDinst/RegFile[27][22] ), .DIN2(n1200), 
        .Q(\IDinst/n11006 ) );
  nnd2s1 \IDinst/U11080  ( .DIN1(\IDinst/RegFile[26][22] ), .DIN2(n1292), 
        .Q(\IDinst/n11005 ) );
  nnd2s1 \IDinst/U11079  ( .DIN1(\IDinst/n11003 ), .DIN2(\IDinst/n11002 ), 
        .Q(\IDinst/n11004 ) );
  nnd2s1 \IDinst/U11078  ( .DIN1(\IDinst/RegFile[25][22] ), .DIN2(n1200), 
        .Q(\IDinst/n11003 ) );
  nnd2s1 \IDinst/U11077  ( .DIN1(\IDinst/RegFile[24][22] ), .DIN2(n1292), 
        .Q(\IDinst/n11002 ) );
  nnd2s1 \IDinst/U11076  ( .DIN1(\IDinst/n11000 ), .DIN2(\IDinst/n10999 ), 
        .Q(\IDinst/n11001 ) );
  nnd2s1 \IDinst/U11075  ( .DIN1(\IDinst/n10998 ), .DIN2(\IDinst/N46 ), 
        .Q(\IDinst/n11000 ) );
  nnd2s1 \IDinst/U11074  ( .DIN1(\IDinst/n10989 ), .DIN2(n1370), 
        .Q(\IDinst/n10999 ) );
  nnd2s1 \IDinst/U11073  ( .DIN1(\IDinst/n10997 ), .DIN2(\IDinst/n10996 ), 
        .Q(\IDinst/n10998 ) );
  nnd2s1 \IDinst/U11072  ( .DIN1(\IDinst/n10995 ), .DIN2(n1316), 
        .Q(\IDinst/n10997 ) );
  nnd2s1 \IDinst/U11071  ( .DIN1(\IDinst/n10992 ), .DIN2(n1355), 
        .Q(\IDinst/n10996 ) );
  nnd2s1 \IDinst/U11070  ( .DIN1(\IDinst/n10994 ), .DIN2(\IDinst/n10993 ), 
        .Q(\IDinst/n10995 ) );
  nnd2s1 \IDinst/U11069  ( .DIN1(\IDinst/RegFile[23][22] ), .DIN2(n1200), 
        .Q(\IDinst/n10994 ) );
  nnd2s1 \IDinst/U11068  ( .DIN1(\IDinst/RegFile[22][22] ), .DIN2(n1292), 
        .Q(\IDinst/n10993 ) );
  nnd2s1 \IDinst/U11067  ( .DIN1(\IDinst/n10991 ), .DIN2(\IDinst/n10990 ), 
        .Q(\IDinst/n10992 ) );
  nnd2s1 \IDinst/U11066  ( .DIN1(\IDinst/RegFile[21][22] ), .DIN2(n1200), 
        .Q(\IDinst/n10991 ) );
  nnd2s1 \IDinst/U11065  ( .DIN1(\IDinst/RegFile[20][22] ), .DIN2(n1292), 
        .Q(\IDinst/n10990 ) );
  nnd2s1 \IDinst/U11064  ( .DIN1(\IDinst/n10988 ), .DIN2(\IDinst/n10987 ), 
        .Q(\IDinst/n10989 ) );
  nnd2s1 \IDinst/U11063  ( .DIN1(\IDinst/n10986 ), .DIN2(n1316), 
        .Q(\IDinst/n10988 ) );
  nnd2s1 \IDinst/U11062  ( .DIN1(\IDinst/n10983 ), .DIN2(n1355), 
        .Q(\IDinst/n10987 ) );
  nnd2s1 \IDinst/U11061  ( .DIN1(\IDinst/n10985 ), .DIN2(\IDinst/n10984 ), 
        .Q(\IDinst/n10986 ) );
  nnd2s1 \IDinst/U11060  ( .DIN1(\IDinst/RegFile[19][22] ), .DIN2(n1200), 
        .Q(\IDinst/n10985 ) );
  nnd2s1 \IDinst/U11059  ( .DIN1(\IDinst/RegFile[18][22] ), .DIN2(n1292), 
        .Q(\IDinst/n10984 ) );
  nnd2s1 \IDinst/U11058  ( .DIN1(\IDinst/n10982 ), .DIN2(\IDinst/n10981 ), 
        .Q(\IDinst/n10983 ) );
  nnd2s1 \IDinst/U11057  ( .DIN1(\IDinst/RegFile[17][22] ), .DIN2(n1200), 
        .Q(\IDinst/n10982 ) );
  nnd2s1 \IDinst/U11056  ( .DIN1(\IDinst/RegFile[16][22] ), .DIN2(n1293), 
        .Q(\IDinst/n10981 ) );
  nnd2s1 \IDinst/U11055  ( .DIN1(\IDinst/n10979 ), .DIN2(\IDinst/n10978 ), 
        .Q(\IDinst/n10980 ) );
  nnd2s1 \IDinst/U11054  ( .DIN1(\IDinst/n10977 ), .DIN2(n666), 
        .Q(\IDinst/n10979 ) );
  nnd2s1 \IDinst/U11053  ( .DIN1(\IDinst/n10956 ), .DIN2(n681), 
        .Q(\IDinst/n10978 ) );
  nnd2s1 \IDinst/U11052  ( .DIN1(\IDinst/n10976 ), .DIN2(\IDinst/n10975 ), 
        .Q(\IDinst/n10977 ) );
  nnd2s1 \IDinst/U11051  ( .DIN1(\IDinst/n10974 ), .DIN2(n1372), 
        .Q(\IDinst/n10976 ) );
  nnd2s1 \IDinst/U11050  ( .DIN1(\IDinst/n10965 ), .DIN2(n1370), 
        .Q(\IDinst/n10975 ) );
  nnd2s1 \IDinst/U11049  ( .DIN1(\IDinst/n10973 ), .DIN2(\IDinst/n10972 ), 
        .Q(\IDinst/n10974 ) );
  nnd2s1 \IDinst/U11048  ( .DIN1(\IDinst/n10971 ), .DIN2(n1316), 
        .Q(\IDinst/n10973 ) );
  nnd2s1 \IDinst/U11047  ( .DIN1(\IDinst/n10968 ), .DIN2(n1355), 
        .Q(\IDinst/n10972 ) );
  nnd2s1 \IDinst/U11046  ( .DIN1(\IDinst/n10970 ), .DIN2(\IDinst/n10969 ), 
        .Q(\IDinst/n10971 ) );
  nnd2s1 \IDinst/U11045  ( .DIN1(\IDinst/RegFile[15][22] ), .DIN2(n1200), 
        .Q(\IDinst/n10970 ) );
  nnd2s1 \IDinst/U11044  ( .DIN1(\IDinst/RegFile[14][22] ), .DIN2(n1293), 
        .Q(\IDinst/n10969 ) );
  nnd2s1 \IDinst/U11043  ( .DIN1(\IDinst/n10967 ), .DIN2(\IDinst/n10966 ), 
        .Q(\IDinst/n10968 ) );
  nnd2s1 \IDinst/U11042  ( .DIN1(\IDinst/RegFile[13][22] ), .DIN2(n1200), 
        .Q(\IDinst/n10967 ) );
  nnd2s1 \IDinst/U11041  ( .DIN1(\IDinst/RegFile[12][22] ), .DIN2(n1293), 
        .Q(\IDinst/n10966 ) );
  nnd2s1 \IDinst/U11040  ( .DIN1(\IDinst/n10964 ), .DIN2(\IDinst/n10963 ), 
        .Q(\IDinst/n10965 ) );
  nnd2s1 \IDinst/U11039  ( .DIN1(\IDinst/n10962 ), .DIN2(n1316), 
        .Q(\IDinst/n10964 ) );
  nnd2s1 \IDinst/U11038  ( .DIN1(\IDinst/n10959 ), .DIN2(n1356), 
        .Q(\IDinst/n10963 ) );
  nnd2s1 \IDinst/U11037  ( .DIN1(\IDinst/n10961 ), .DIN2(\IDinst/n10960 ), 
        .Q(\IDinst/n10962 ) );
  nnd2s1 \IDinst/U11036  ( .DIN1(\IDinst/RegFile[11][22] ), .DIN2(n1200), 
        .Q(\IDinst/n10961 ) );
  nnd2s1 \IDinst/U11035  ( .DIN1(\IDinst/RegFile[10][22] ), .DIN2(n1293), 
        .Q(\IDinst/n10960 ) );
  nnd2s1 \IDinst/U11034  ( .DIN1(\IDinst/n10958 ), .DIN2(\IDinst/n10957 ), 
        .Q(\IDinst/n10959 ) );
  nnd2s1 \IDinst/U11033  ( .DIN1(\IDinst/RegFile[9][22] ), .DIN2(n1200), 
        .Q(\IDinst/n10958 ) );
  nnd2s1 \IDinst/U11032  ( .DIN1(\IDinst/RegFile[8][22] ), .DIN2(n1293), 
        .Q(\IDinst/n10957 ) );
  nnd2s1 \IDinst/U11031  ( .DIN1(\IDinst/n10955 ), .DIN2(\IDinst/n10954 ), 
        .Q(\IDinst/n10956 ) );
  nnd2s1 \IDinst/U11030  ( .DIN1(\IDinst/n10953 ), .DIN2(n1379), 
        .Q(\IDinst/n10955 ) );
  nnd2s1 \IDinst/U11029  ( .DIN1(\IDinst/n10944 ), .DIN2(n1370), 
        .Q(\IDinst/n10954 ) );
  nnd2s1 \IDinst/U11028  ( .DIN1(\IDinst/n10952 ), .DIN2(\IDinst/n10951 ), 
        .Q(\IDinst/n10953 ) );
  nnd2s1 \IDinst/U11027  ( .DIN1(\IDinst/n10950 ), .DIN2(n1316), 
        .Q(\IDinst/n10952 ) );
  nnd2s1 \IDinst/U11026  ( .DIN1(\IDinst/n10947 ), .DIN2(n1356), 
        .Q(\IDinst/n10951 ) );
  nnd2s1 \IDinst/U11025  ( .DIN1(\IDinst/n10949 ), .DIN2(\IDinst/n10948 ), 
        .Q(\IDinst/n10950 ) );
  nnd2s1 \IDinst/U11024  ( .DIN1(\IDinst/RegFile[7][22] ), .DIN2(n1200), 
        .Q(\IDinst/n10949 ) );
  nnd2s1 \IDinst/U11023  ( .DIN1(\IDinst/RegFile[6][22] ), .DIN2(n1293), 
        .Q(\IDinst/n10948 ) );
  nnd2s1 \IDinst/U11022  ( .DIN1(\IDinst/n10946 ), .DIN2(\IDinst/n10945 ), 
        .Q(\IDinst/n10947 ) );
  nnd2s1 \IDinst/U11021  ( .DIN1(\IDinst/RegFile[5][22] ), .DIN2(n1200), 
        .Q(\IDinst/n10946 ) );
  nnd2s1 \IDinst/U11020  ( .DIN1(\IDinst/RegFile[4][22] ), .DIN2(n1293), 
        .Q(\IDinst/n10945 ) );
  nnd2s1 \IDinst/U11019  ( .DIN1(\IDinst/n10943 ), .DIN2(\IDinst/n10942 ), 
        .Q(\IDinst/n10944 ) );
  nnd2s1 \IDinst/U11018  ( .DIN1(\IDinst/n10941 ), .DIN2(n1316), 
        .Q(\IDinst/n10943 ) );
  nnd2s1 \IDinst/U11017  ( .DIN1(\IDinst/n10938 ), .DIN2(n1356), 
        .Q(\IDinst/n10942 ) );
  nnd2s1 \IDinst/U11016  ( .DIN1(\IDinst/n10940 ), .DIN2(\IDinst/n10939 ), 
        .Q(\IDinst/n10941 ) );
  nnd2s1 \IDinst/U11015  ( .DIN1(\IDinst/RegFile[3][22] ), .DIN2(n1200), 
        .Q(\IDinst/n10940 ) );
  nnd2s1 \IDinst/U11014  ( .DIN1(\IDinst/RegFile[2][22] ), .DIN2(n1293), 
        .Q(\IDinst/n10939 ) );
  nnd2s1 \IDinst/U11013  ( .DIN1(\IDinst/n10937 ), .DIN2(\IDinst/n10936 ), 
        .Q(\IDinst/n10938 ) );
  nnd2s1 \IDinst/U11012  ( .DIN1(\IDinst/RegFile[1][22] ), .DIN2(n1201), 
        .Q(\IDinst/n10937 ) );
  nnd2s1 \IDinst/U11011  ( .DIN1(\IDinst/RegFile[0][22] ), .DIN2(n1293), 
        .Q(\IDinst/n10936 ) );
  nnd2s1 \IDinst/U11010  ( .DIN1(\IDinst/n10935 ), .DIN2(n535), 
        .Q(\IDinst/n8934 ) );
  nnd2s1 \IDinst/U11009  ( .DIN1(\IDinst/n10890 ), .DIN2(n533), 
        .Q(\IDinst/n8935 ) );
  nnd2s1 \IDinst/U11008  ( .DIN1(\IDinst/n10934 ), .DIN2(\IDinst/n10933 ), 
        .Q(\IDinst/n10935 ) );
  nnd2s1 \IDinst/U11007  ( .DIN1(\IDinst/n10932 ), .DIN2(n667), 
        .Q(\IDinst/n10934 ) );
  nnd2s1 \IDinst/U11006  ( .DIN1(\IDinst/n10911 ), .DIN2(n683), 
        .Q(\IDinst/n10933 ) );
  nnd2s1 \IDinst/U11005  ( .DIN1(\IDinst/n10931 ), .DIN2(\IDinst/n10930 ), 
        .Q(\IDinst/n10932 ) );
  nnd2s1 \IDinst/U11004  ( .DIN1(\IDinst/n10929 ), .DIN2(n1375), 
        .Q(\IDinst/n10931 ) );
  nnd2s1 \IDinst/U11003  ( .DIN1(\IDinst/n10920 ), .DIN2(n1370), 
        .Q(\IDinst/n10930 ) );
  nnd2s1 \IDinst/U11002  ( .DIN1(\IDinst/n10928 ), .DIN2(\IDinst/n10927 ), 
        .Q(\IDinst/n10929 ) );
  nnd2s1 \IDinst/U11001  ( .DIN1(\IDinst/n10926 ), .DIN2(n1316), 
        .Q(\IDinst/n10928 ) );
  nnd2s1 \IDinst/U11000  ( .DIN1(\IDinst/n10923 ), .DIN2(n1356), 
        .Q(\IDinst/n10927 ) );
  nnd2s1 \IDinst/U10999  ( .DIN1(\IDinst/n10925 ), .DIN2(\IDinst/n10924 ), 
        .Q(\IDinst/n10926 ) );
  nnd2s1 \IDinst/U10998  ( .DIN1(\IDinst/RegFile[31][21] ), .DIN2(n1201), 
        .Q(\IDinst/n10925 ) );
  nnd2s1 \IDinst/U10997  ( .DIN1(\IDinst/RegFile[30][21] ), .DIN2(n1294), 
        .Q(\IDinst/n10924 ) );
  nnd2s1 \IDinst/U10996  ( .DIN1(\IDinst/n10922 ), .DIN2(\IDinst/n10921 ), 
        .Q(\IDinst/n10923 ) );
  nnd2s1 \IDinst/U10995  ( .DIN1(\IDinst/RegFile[29][21] ), .DIN2(n1201), 
        .Q(\IDinst/n10922 ) );
  nnd2s1 \IDinst/U10994  ( .DIN1(\IDinst/RegFile[28][21] ), .DIN2(n1294), 
        .Q(\IDinst/n10921 ) );
  nnd2s1 \IDinst/U10993  ( .DIN1(\IDinst/n10919 ), .DIN2(\IDinst/n10918 ), 
        .Q(\IDinst/n10920 ) );
  nnd2s1 \IDinst/U10992  ( .DIN1(\IDinst/n10917 ), .DIN2(n1316), 
        .Q(\IDinst/n10919 ) );
  nnd2s1 \IDinst/U10991  ( .DIN1(\IDinst/n10914 ), .DIN2(n1356), 
        .Q(\IDinst/n10918 ) );
  nnd2s1 \IDinst/U10990  ( .DIN1(\IDinst/n10916 ), .DIN2(\IDinst/n10915 ), 
        .Q(\IDinst/n10917 ) );
  nnd2s1 \IDinst/U10989  ( .DIN1(\IDinst/RegFile[27][21] ), .DIN2(n1201), 
        .Q(\IDinst/n10916 ) );
  nnd2s1 \IDinst/U10988  ( .DIN1(\IDinst/RegFile[26][21] ), .DIN2(n1294), 
        .Q(\IDinst/n10915 ) );
  nnd2s1 \IDinst/U10987  ( .DIN1(\IDinst/n10913 ), .DIN2(\IDinst/n10912 ), 
        .Q(\IDinst/n10914 ) );
  nnd2s1 \IDinst/U10986  ( .DIN1(\IDinst/RegFile[25][21] ), .DIN2(n1201), 
        .Q(\IDinst/n10913 ) );
  nnd2s1 \IDinst/U10985  ( .DIN1(\IDinst/RegFile[24][21] ), .DIN2(n1294), 
        .Q(\IDinst/n10912 ) );
  nnd2s1 \IDinst/U10984  ( .DIN1(\IDinst/n10910 ), .DIN2(\IDinst/n10909 ), 
        .Q(\IDinst/n10911 ) );
  nnd2s1 \IDinst/U10983  ( .DIN1(\IDinst/n10908 ), .DIN2(n1373), 
        .Q(\IDinst/n10910 ) );
  nnd2s1 \IDinst/U10982  ( .DIN1(\IDinst/n10899 ), .DIN2(n1370), 
        .Q(\IDinst/n10909 ) );
  nnd2s1 \IDinst/U10981  ( .DIN1(\IDinst/n10907 ), .DIN2(\IDinst/n10906 ), 
        .Q(\IDinst/n10908 ) );
  nnd2s1 \IDinst/U10980  ( .DIN1(\IDinst/n10905 ), .DIN2(n1316), 
        .Q(\IDinst/n10907 ) );
  nnd2s1 \IDinst/U10979  ( .DIN1(\IDinst/n10902 ), .DIN2(n1356), 
        .Q(\IDinst/n10906 ) );
  nnd2s1 \IDinst/U10978  ( .DIN1(\IDinst/n10904 ), .DIN2(\IDinst/n10903 ), 
        .Q(\IDinst/n10905 ) );
  nnd2s1 \IDinst/U10977  ( .DIN1(\IDinst/RegFile[23][21] ), .DIN2(n1201), 
        .Q(\IDinst/n10904 ) );
  nnd2s1 \IDinst/U10976  ( .DIN1(\IDinst/RegFile[22][21] ), .DIN2(n1294), 
        .Q(\IDinst/n10903 ) );
  nnd2s1 \IDinst/U10975  ( .DIN1(\IDinst/n10901 ), .DIN2(\IDinst/n10900 ), 
        .Q(\IDinst/n10902 ) );
  nnd2s1 \IDinst/U10974  ( .DIN1(\IDinst/RegFile[21][21] ), .DIN2(n1201), 
        .Q(\IDinst/n10901 ) );
  nnd2s1 \IDinst/U10973  ( .DIN1(\IDinst/RegFile[20][21] ), .DIN2(n1294), 
        .Q(\IDinst/n10900 ) );
  nnd2s1 \IDinst/U10972  ( .DIN1(\IDinst/n10898 ), .DIN2(\IDinst/n10897 ), 
        .Q(\IDinst/n10899 ) );
  nnd2s1 \IDinst/U10971  ( .DIN1(\IDinst/n10896 ), .DIN2(n1316), 
        .Q(\IDinst/n10898 ) );
  nnd2s1 \IDinst/U10970  ( .DIN1(\IDinst/n10893 ), .DIN2(n1356), 
        .Q(\IDinst/n10897 ) );
  nnd2s1 \IDinst/U10969  ( .DIN1(\IDinst/n10895 ), .DIN2(\IDinst/n10894 ), 
        .Q(\IDinst/n10896 ) );
  nnd2s1 \IDinst/U10968  ( .DIN1(\IDinst/RegFile[19][21] ), .DIN2(n1201), 
        .Q(\IDinst/n10895 ) );
  nnd2s1 \IDinst/U10967  ( .DIN1(\IDinst/RegFile[18][21] ), .DIN2(n1294), 
        .Q(\IDinst/n10894 ) );
  nnd2s1 \IDinst/U10966  ( .DIN1(\IDinst/n10892 ), .DIN2(\IDinst/n10891 ), 
        .Q(\IDinst/n10893 ) );
  nnd2s1 \IDinst/U10965  ( .DIN1(\IDinst/RegFile[17][21] ), .DIN2(n1201), 
        .Q(\IDinst/n10892 ) );
  nnd2s1 \IDinst/U10964  ( .DIN1(\IDinst/RegFile[16][21] ), .DIN2(n1294), 
        .Q(\IDinst/n10891 ) );
  nnd2s1 \IDinst/U10963  ( .DIN1(\IDinst/n10889 ), .DIN2(\IDinst/n10888 ), 
        .Q(\IDinst/n10890 ) );
  nnd2s1 \IDinst/U10962  ( .DIN1(\IDinst/n10887 ), .DIN2(n665), 
        .Q(\IDinst/n10889 ) );
  nnd2s1 \IDinst/U10961  ( .DIN1(\IDinst/n10866 ), .DIN2(n682), 
        .Q(\IDinst/n10888 ) );
  nnd2s1 \IDinst/U10960  ( .DIN1(\IDinst/n10886 ), .DIN2(\IDinst/n10885 ), 
        .Q(\IDinst/n10887 ) );
  nnd2s1 \IDinst/U10959  ( .DIN1(\IDinst/n10884 ), .DIN2(n1376), 
        .Q(\IDinst/n10886 ) );
  nnd2s1 \IDinst/U10958  ( .DIN1(\IDinst/n10875 ), .DIN2(n1370), 
        .Q(\IDinst/n10885 ) );
  nnd2s1 \IDinst/U10957  ( .DIN1(\IDinst/n10883 ), .DIN2(\IDinst/n10882 ), 
        .Q(\IDinst/n10884 ) );
  nnd2s1 \IDinst/U10956  ( .DIN1(\IDinst/n10881 ), .DIN2(n1315), 
        .Q(\IDinst/n10883 ) );
  nnd2s1 \IDinst/U10955  ( .DIN1(\IDinst/n10878 ), .DIN2(n1356), 
        .Q(\IDinst/n10882 ) );
  nnd2s1 \IDinst/U10954  ( .DIN1(\IDinst/n10880 ), .DIN2(\IDinst/n10879 ), 
        .Q(\IDinst/n10881 ) );
  nnd2s1 \IDinst/U10953  ( .DIN1(\IDinst/RegFile[15][21] ), .DIN2(n1201), 
        .Q(\IDinst/n10880 ) );
  nnd2s1 \IDinst/U10952  ( .DIN1(\IDinst/RegFile[14][21] ), .DIN2(n1294), 
        .Q(\IDinst/n10879 ) );
  nnd2s1 \IDinst/U10951  ( .DIN1(\IDinst/n10877 ), .DIN2(\IDinst/n10876 ), 
        .Q(\IDinst/n10878 ) );
  nnd2s1 \IDinst/U10950  ( .DIN1(\IDinst/RegFile[13][21] ), .DIN2(n1201), 
        .Q(\IDinst/n10877 ) );
  nnd2s1 \IDinst/U10949  ( .DIN1(\IDinst/RegFile[12][21] ), .DIN2(n1295), 
        .Q(\IDinst/n10876 ) );
  nnd2s1 \IDinst/U10948  ( .DIN1(\IDinst/n10874 ), .DIN2(\IDinst/n10873 ), 
        .Q(\IDinst/n10875 ) );
  nnd2s1 \IDinst/U10947  ( .DIN1(\IDinst/n10872 ), .DIN2(n1315), 
        .Q(\IDinst/n10874 ) );
  nnd2s1 \IDinst/U10946  ( .DIN1(\IDinst/n10869 ), .DIN2(n1356), 
        .Q(\IDinst/n10873 ) );
  nnd2s1 \IDinst/U10945  ( .DIN1(\IDinst/n10871 ), .DIN2(\IDinst/n10870 ), 
        .Q(\IDinst/n10872 ) );
  nnd2s1 \IDinst/U10944  ( .DIN1(\IDinst/RegFile[11][21] ), .DIN2(n1201), 
        .Q(\IDinst/n10871 ) );
  nnd2s1 \IDinst/U10943  ( .DIN1(\IDinst/RegFile[10][21] ), .DIN2(n1295), 
        .Q(\IDinst/n10870 ) );
  nnd2s1 \IDinst/U10942  ( .DIN1(\IDinst/n10868 ), .DIN2(\IDinst/n10867 ), 
        .Q(\IDinst/n10869 ) );
  nnd2s1 \IDinst/U10941  ( .DIN1(\IDinst/RegFile[9][21] ), .DIN2(n1201), 
        .Q(\IDinst/n10868 ) );
  nnd2s1 \IDinst/U10940  ( .DIN1(\IDinst/RegFile[8][21] ), .DIN2(n1295), 
        .Q(\IDinst/n10867 ) );
  nnd2s1 \IDinst/U10939  ( .DIN1(\IDinst/n10865 ), .DIN2(\IDinst/n10864 ), 
        .Q(\IDinst/n10866 ) );
  nnd2s1 \IDinst/U10938  ( .DIN1(\IDinst/n10863 ), .DIN2(n1377), 
        .Q(\IDinst/n10865 ) );
  nnd2s1 \IDinst/U10937  ( .DIN1(\IDinst/n10854 ), .DIN2(n1370), 
        .Q(\IDinst/n10864 ) );
  nnd2s1 \IDinst/U10936  ( .DIN1(\IDinst/n10862 ), .DIN2(\IDinst/n10861 ), 
        .Q(\IDinst/n10863 ) );
  nnd2s1 \IDinst/U10935  ( .DIN1(\IDinst/n10860 ), .DIN2(n1315), 
        .Q(\IDinst/n10862 ) );
  nnd2s1 \IDinst/U10934  ( .DIN1(\IDinst/n10857 ), .DIN2(n1357), 
        .Q(\IDinst/n10861 ) );
  nnd2s1 \IDinst/U10933  ( .DIN1(\IDinst/n10859 ), .DIN2(\IDinst/n10858 ), 
        .Q(\IDinst/n10860 ) );
  nnd2s1 \IDinst/U10932  ( .DIN1(\IDinst/RegFile[7][21] ), .DIN2(n1202), 
        .Q(\IDinst/n10859 ) );
  nnd2s1 \IDinst/U10931  ( .DIN1(\IDinst/RegFile[6][21] ), .DIN2(n1295), 
        .Q(\IDinst/n10858 ) );
  nnd2s1 \IDinst/U10930  ( .DIN1(\IDinst/n10856 ), .DIN2(\IDinst/n10855 ), 
        .Q(\IDinst/n10857 ) );
  nnd2s1 \IDinst/U10929  ( .DIN1(\IDinst/RegFile[5][21] ), .DIN2(n1202), 
        .Q(\IDinst/n10856 ) );
  nnd2s1 \IDinst/U10928  ( .DIN1(\IDinst/RegFile[4][21] ), .DIN2(n1295), 
        .Q(\IDinst/n10855 ) );
  nnd2s1 \IDinst/U10927  ( .DIN1(\IDinst/n10853 ), .DIN2(\IDinst/n10852 ), 
        .Q(\IDinst/n10854 ) );
  nnd2s1 \IDinst/U10926  ( .DIN1(\IDinst/n10851 ), .DIN2(n1315), 
        .Q(\IDinst/n10853 ) );
  nnd2s1 \IDinst/U10925  ( .DIN1(\IDinst/n10848 ), .DIN2(n1357), 
        .Q(\IDinst/n10852 ) );
  nnd2s1 \IDinst/U10924  ( .DIN1(\IDinst/n10850 ), .DIN2(\IDinst/n10849 ), 
        .Q(\IDinst/n10851 ) );
  nnd2s1 \IDinst/U10923  ( .DIN1(\IDinst/RegFile[3][21] ), .DIN2(n1202), 
        .Q(\IDinst/n10850 ) );
  nnd2s1 \IDinst/U10922  ( .DIN1(\IDinst/RegFile[2][21] ), .DIN2(n1295), 
        .Q(\IDinst/n10849 ) );
  nnd2s1 \IDinst/U10921  ( .DIN1(\IDinst/n10847 ), .DIN2(\IDinst/n10846 ), 
        .Q(\IDinst/n10848 ) );
  nnd2s1 \IDinst/U10920  ( .DIN1(\IDinst/RegFile[1][21] ), .DIN2(n1202), 
        .Q(\IDinst/n10847 ) );
  nnd2s1 \IDinst/U10919  ( .DIN1(\IDinst/RegFile[0][21] ), .DIN2(n1295), 
        .Q(\IDinst/n10846 ) );
  nnd2s1 \IDinst/U10918  ( .DIN1(\IDinst/n10845 ), .DIN2(n534), 
        .Q(\IDinst/n8932 ) );
  nnd2s1 \IDinst/U10917  ( .DIN1(\IDinst/n10800 ), .DIN2(n634), 
        .Q(\IDinst/n8933 ) );
  nnd2s1 \IDinst/U10916  ( .DIN1(\IDinst/n10844 ), .DIN2(\IDinst/n10843 ), 
        .Q(\IDinst/n10845 ) );
  nnd2s1 \IDinst/U10915  ( .DIN1(\IDinst/n10842 ), .DIN2(n668), 
        .Q(\IDinst/n10844 ) );
  nnd2s1 \IDinst/U10914  ( .DIN1(\IDinst/n10821 ), .DIN2(n680), 
        .Q(\IDinst/n10843 ) );
  nnd2s1 \IDinst/U10913  ( .DIN1(\IDinst/n10841 ), .DIN2(\IDinst/n10840 ), 
        .Q(\IDinst/n10842 ) );
  nnd2s1 \IDinst/U10912  ( .DIN1(\IDinst/n10839 ), .DIN2(\IDinst/N46 ), 
        .Q(\IDinst/n10841 ) );
  nnd2s1 \IDinst/U10911  ( .DIN1(\IDinst/n10830 ), .DIN2(n1370), 
        .Q(\IDinst/n10840 ) );
  nnd2s1 \IDinst/U10910  ( .DIN1(\IDinst/n10838 ), .DIN2(\IDinst/n10837 ), 
        .Q(\IDinst/n10839 ) );
  nnd2s1 \IDinst/U10909  ( .DIN1(\IDinst/n10836 ), .DIN2(n1315), 
        .Q(\IDinst/n10838 ) );
  nnd2s1 \IDinst/U10908  ( .DIN1(\IDinst/n10833 ), .DIN2(n1357), 
        .Q(\IDinst/n10837 ) );
  nnd2s1 \IDinst/U10907  ( .DIN1(\IDinst/n10835 ), .DIN2(\IDinst/n10834 ), 
        .Q(\IDinst/n10836 ) );
  nnd2s1 \IDinst/U10906  ( .DIN1(\IDinst/RegFile[31][20] ), .DIN2(n1202), 
        .Q(\IDinst/n10835 ) );
  nnd2s1 \IDinst/U10905  ( .DIN1(\IDinst/RegFile[30][20] ), .DIN2(n1295), 
        .Q(\IDinst/n10834 ) );
  nnd2s1 \IDinst/U10904  ( .DIN1(\IDinst/n10832 ), .DIN2(\IDinst/n10831 ), 
        .Q(\IDinst/n10833 ) );
  nnd2s1 \IDinst/U10903  ( .DIN1(\IDinst/RegFile[29][20] ), .DIN2(n1202), 
        .Q(\IDinst/n10832 ) );
  nnd2s1 \IDinst/U10902  ( .DIN1(\IDinst/RegFile[28][20] ), .DIN2(n1289), 
        .Q(\IDinst/n10831 ) );
  nnd2s1 \IDinst/U10901  ( .DIN1(\IDinst/n10829 ), .DIN2(\IDinst/n10828 ), 
        .Q(\IDinst/n10830 ) );
  nnd2s1 \IDinst/U10900  ( .DIN1(\IDinst/n10827 ), .DIN2(n1315), 
        .Q(\IDinst/n10829 ) );
  nnd2s1 \IDinst/U10899  ( .DIN1(\IDinst/n10824 ), .DIN2(n1357), 
        .Q(\IDinst/n10828 ) );
  nnd2s1 \IDinst/U10898  ( .DIN1(\IDinst/n10826 ), .DIN2(\IDinst/n10825 ), 
        .Q(\IDinst/n10827 ) );
  nnd2s1 \IDinst/U10897  ( .DIN1(\IDinst/RegFile[27][20] ), .DIN2(n1202), 
        .Q(\IDinst/n10826 ) );
  nnd2s1 \IDinst/U10896  ( .DIN1(\IDinst/RegFile[26][20] ), .DIN2(n1289), 
        .Q(\IDinst/n10825 ) );
  nnd2s1 \IDinst/U10895  ( .DIN1(\IDinst/n10823 ), .DIN2(\IDinst/n10822 ), 
        .Q(\IDinst/n10824 ) );
  nnd2s1 \IDinst/U10894  ( .DIN1(\IDinst/RegFile[25][20] ), .DIN2(n1202), 
        .Q(\IDinst/n10823 ) );
  nnd2s1 \IDinst/U10893  ( .DIN1(\IDinst/RegFile[24][20] ), .DIN2(n1288), 
        .Q(\IDinst/n10822 ) );
  nnd2s1 \IDinst/U10892  ( .DIN1(\IDinst/n10820 ), .DIN2(\IDinst/n10819 ), 
        .Q(\IDinst/n10821 ) );
  nnd2s1 \IDinst/U10891  ( .DIN1(\IDinst/n10818 ), .DIN2(n1380), 
        .Q(\IDinst/n10820 ) );
  nnd2s1 \IDinst/U10890  ( .DIN1(\IDinst/n10809 ), .DIN2(n1370), 
        .Q(\IDinst/n10819 ) );
  nnd2s1 \IDinst/U10889  ( .DIN1(\IDinst/n10817 ), .DIN2(\IDinst/n10816 ), 
        .Q(\IDinst/n10818 ) );
  nnd2s1 \IDinst/U10888  ( .DIN1(\IDinst/n10815 ), .DIN2(n1315), 
        .Q(\IDinst/n10817 ) );
  nnd2s1 \IDinst/U10887  ( .DIN1(\IDinst/n10812 ), .DIN2(n1357), 
        .Q(\IDinst/n10816 ) );
  nnd2s1 \IDinst/U10886  ( .DIN1(\IDinst/n10814 ), .DIN2(\IDinst/n10813 ), 
        .Q(\IDinst/n10815 ) );
  nnd2s1 \IDinst/U10885  ( .DIN1(\IDinst/RegFile[23][20] ), .DIN2(n1202), 
        .Q(\IDinst/n10814 ) );
  nnd2s1 \IDinst/U10884  ( .DIN1(\IDinst/RegFile[22][20] ), .DIN2(n1288), 
        .Q(\IDinst/n10813 ) );
  nnd2s1 \IDinst/U10883  ( .DIN1(\IDinst/n10811 ), .DIN2(\IDinst/n10810 ), 
        .Q(\IDinst/n10812 ) );
  nnd2s1 \IDinst/U10882  ( .DIN1(\IDinst/RegFile[21][20] ), .DIN2(n1202), 
        .Q(\IDinst/n10811 ) );
  nnd2s1 \IDinst/U10881  ( .DIN1(\IDinst/RegFile[20][20] ), .DIN2(n1288), 
        .Q(\IDinst/n10810 ) );
  nnd2s1 \IDinst/U10880  ( .DIN1(\IDinst/n10808 ), .DIN2(\IDinst/n10807 ), 
        .Q(\IDinst/n10809 ) );
  nnd2s1 \IDinst/U10879  ( .DIN1(\IDinst/n10806 ), .DIN2(n1315), 
        .Q(\IDinst/n10808 ) );
  nnd2s1 \IDinst/U10878  ( .DIN1(\IDinst/n10803 ), .DIN2(n1357), 
        .Q(\IDinst/n10807 ) );
  nnd2s1 \IDinst/U10877  ( .DIN1(\IDinst/n10805 ), .DIN2(\IDinst/n10804 ), 
        .Q(\IDinst/n10806 ) );
  nnd2s1 \IDinst/U10876  ( .DIN1(\IDinst/RegFile[19][20] ), .DIN2(n1202), 
        .Q(\IDinst/n10805 ) );
  nnd2s1 \IDinst/U10875  ( .DIN1(\IDinst/RegFile[18][20] ), .DIN2(n1288), 
        .Q(\IDinst/n10804 ) );
  nnd2s1 \IDinst/U10874  ( .DIN1(\IDinst/n10802 ), .DIN2(\IDinst/n10801 ), 
        .Q(\IDinst/n10803 ) );
  nnd2s1 \IDinst/U10873  ( .DIN1(\IDinst/RegFile[17][20] ), .DIN2(n1202), 
        .Q(\IDinst/n10802 ) );
  nnd2s1 \IDinst/U10872  ( .DIN1(\IDinst/RegFile[16][20] ), .DIN2(n1288), 
        .Q(\IDinst/n10801 ) );
  nnd2s1 \IDinst/U10871  ( .DIN1(\IDinst/n10799 ), .DIN2(\IDinst/n10798 ), 
        .Q(\IDinst/n10800 ) );
  nnd2s1 \IDinst/U10870  ( .DIN1(\IDinst/n10797 ), .DIN2(n666), 
        .Q(\IDinst/n10799 ) );
  nnd2s1 \IDinst/U10869  ( .DIN1(\IDinst/n10776 ), .DIN2(n681), 
        .Q(\IDinst/n10798 ) );
  nnd2s1 \IDinst/U10868  ( .DIN1(\IDinst/n10796 ), .DIN2(\IDinst/n10795 ), 
        .Q(\IDinst/n10797 ) );
  nnd2s1 \IDinst/U10867  ( .DIN1(\IDinst/n10794 ), .DIN2(\IDinst/N46 ), 
        .Q(\IDinst/n10796 ) );
  nnd2s1 \IDinst/U10866  ( .DIN1(\IDinst/n10785 ), .DIN2(n1370), 
        .Q(\IDinst/n10795 ) );
  nnd2s1 \IDinst/U10865  ( .DIN1(\IDinst/n10793 ), .DIN2(\IDinst/n10792 ), 
        .Q(\IDinst/n10794 ) );
  nnd2s1 \IDinst/U10864  ( .DIN1(\IDinst/n10791 ), .DIN2(n1315), 
        .Q(\IDinst/n10793 ) );
  nnd2s1 \IDinst/U10863  ( .DIN1(\IDinst/n10788 ), .DIN2(n1357), 
        .Q(\IDinst/n10792 ) );
  nnd2s1 \IDinst/U10862  ( .DIN1(\IDinst/n10790 ), .DIN2(\IDinst/n10789 ), 
        .Q(\IDinst/n10791 ) );
  nnd2s1 \IDinst/U10861  ( .DIN1(\IDinst/RegFile[15][20] ), .DIN2(n1202), 
        .Q(\IDinst/n10790 ) );
  nnd2s1 \IDinst/U10860  ( .DIN1(\IDinst/RegFile[14][20] ), .DIN2(n1288), 
        .Q(\IDinst/n10789 ) );
  nnd2s1 \IDinst/U10859  ( .DIN1(\IDinst/n10787 ), .DIN2(\IDinst/n10786 ), 
        .Q(\IDinst/n10788 ) );
  nnd2s1 \IDinst/U10858  ( .DIN1(\IDinst/RegFile[13][20] ), .DIN2(n1203), 
        .Q(\IDinst/n10787 ) );
  nnd2s1 \IDinst/U10857  ( .DIN1(\IDinst/RegFile[12][20] ), .DIN2(n1288), 
        .Q(\IDinst/n10786 ) );
  nnd2s1 \IDinst/U10856  ( .DIN1(\IDinst/n10784 ), .DIN2(\IDinst/n10783 ), 
        .Q(\IDinst/n10785 ) );
  nnd2s1 \IDinst/U10855  ( .DIN1(\IDinst/n10782 ), .DIN2(n1315), 
        .Q(\IDinst/n10784 ) );
  nnd2s1 \IDinst/U10854  ( .DIN1(\IDinst/n10779 ), .DIN2(n1357), 
        .Q(\IDinst/n10783 ) );
  nnd2s1 \IDinst/U10853  ( .DIN1(\IDinst/n10781 ), .DIN2(\IDinst/n10780 ), 
        .Q(\IDinst/n10782 ) );
  nnd2s1 \IDinst/U10852  ( .DIN1(\IDinst/RegFile[11][20] ), .DIN2(n1203), 
        .Q(\IDinst/n10781 ) );
  nnd2s1 \IDinst/U10851  ( .DIN1(\IDinst/RegFile[10][20] ), .DIN2(n1288), 
        .Q(\IDinst/n10780 ) );
  nnd2s1 \IDinst/U10850  ( .DIN1(\IDinst/n10778 ), .DIN2(\IDinst/n10777 ), 
        .Q(\IDinst/n10779 ) );
  nnd2s1 \IDinst/U10849  ( .DIN1(\IDinst/RegFile[9][20] ), .DIN2(n1203), 
        .Q(\IDinst/n10778 ) );
  nnd2s1 \IDinst/U10848  ( .DIN1(\IDinst/RegFile[8][20] ), .DIN2(n1288), 
        .Q(\IDinst/n10777 ) );
  nnd2s1 \IDinst/U10847  ( .DIN1(\IDinst/n10775 ), .DIN2(\IDinst/n10774 ), 
        .Q(\IDinst/n10776 ) );
  nnd2s1 \IDinst/U10846  ( .DIN1(\IDinst/n10773 ), .DIN2(n1372), 
        .Q(\IDinst/n10775 ) );
  nnd2s1 \IDinst/U10845  ( .DIN1(\IDinst/n10764 ), .DIN2(n1369), 
        .Q(\IDinst/n10774 ) );
  nnd2s1 \IDinst/U10844  ( .DIN1(\IDinst/n10772 ), .DIN2(\IDinst/n10771 ), 
        .Q(\IDinst/n10773 ) );
  nnd2s1 \IDinst/U10843  ( .DIN1(\IDinst/n10770 ), .DIN2(n1315), 
        .Q(\IDinst/n10772 ) );
  nnd2s1 \IDinst/U10842  ( .DIN1(\IDinst/n10767 ), .DIN2(n1357), 
        .Q(\IDinst/n10771 ) );
  nnd2s1 \IDinst/U10841  ( .DIN1(\IDinst/n10769 ), .DIN2(\IDinst/n10768 ), 
        .Q(\IDinst/n10770 ) );
  nnd2s1 \IDinst/U10840  ( .DIN1(\IDinst/RegFile[7][20] ), .DIN2(n1203), 
        .Q(\IDinst/n10769 ) );
  nnd2s1 \IDinst/U10839  ( .DIN1(\IDinst/RegFile[6][20] ), .DIN2(n1287), 
        .Q(\IDinst/n10768 ) );
  nnd2s1 \IDinst/U10838  ( .DIN1(\IDinst/n10766 ), .DIN2(\IDinst/n10765 ), 
        .Q(\IDinst/n10767 ) );
  nnd2s1 \IDinst/U10837  ( .DIN1(\IDinst/RegFile[5][20] ), .DIN2(n1203), 
        .Q(\IDinst/n10766 ) );
  nnd2s1 \IDinst/U10836  ( .DIN1(\IDinst/RegFile[4][20] ), .DIN2(n1287), 
        .Q(\IDinst/n10765 ) );
  nnd2s1 \IDinst/U10835  ( .DIN1(\IDinst/n10763 ), .DIN2(\IDinst/n10762 ), 
        .Q(\IDinst/n10764 ) );
  nnd2s1 \IDinst/U10834  ( .DIN1(\IDinst/n10761 ), .DIN2(n1315), 
        .Q(\IDinst/n10763 ) );
  nnd2s1 \IDinst/U10833  ( .DIN1(\IDinst/n10758 ), .DIN2(n1358), 
        .Q(\IDinst/n10762 ) );
  nnd2s1 \IDinst/U10832  ( .DIN1(\IDinst/n10760 ), .DIN2(\IDinst/n10759 ), 
        .Q(\IDinst/n10761 ) );
  nnd2s1 \IDinst/U10831  ( .DIN1(\IDinst/RegFile[3][20] ), .DIN2(n1203), 
        .Q(\IDinst/n10760 ) );
  nnd2s1 \IDinst/U10830  ( .DIN1(\IDinst/RegFile[2][20] ), .DIN2(n1287), 
        .Q(\IDinst/n10759 ) );
  nnd2s1 \IDinst/U10829  ( .DIN1(\IDinst/n10757 ), .DIN2(\IDinst/n10756 ), 
        .Q(\IDinst/n10758 ) );
  nnd2s1 \IDinst/U10828  ( .DIN1(\IDinst/RegFile[1][20] ), .DIN2(n1203), 
        .Q(\IDinst/n10757 ) );
  nnd2s1 \IDinst/U10827  ( .DIN1(\IDinst/RegFile[0][20] ), .DIN2(n1287), 
        .Q(\IDinst/n10756 ) );
  nnd2s1 \IDinst/U10826  ( .DIN1(\IDinst/n10755 ), .DIN2(\IDinst/N48 ), 
        .Q(\IDinst/n8930 ) );
  nnd2s1 \IDinst/U10825  ( .DIN1(\IDinst/n10710 ), .DIN2(n533), 
        .Q(\IDinst/n8931 ) );
  nnd2s1 \IDinst/U10824  ( .DIN1(\IDinst/n10754 ), .DIN2(\IDinst/n10753 ), 
        .Q(\IDinst/n10755 ) );
  nnd2s1 \IDinst/U10823  ( .DIN1(\IDinst/n10752 ), .DIN2(n667), 
        .Q(\IDinst/n10754 ) );
  nnd2s1 \IDinst/U10822  ( .DIN1(\IDinst/n10731 ), .DIN2(n683), 
        .Q(\IDinst/n10753 ) );
  nnd2s1 \IDinst/U10821  ( .DIN1(\IDinst/n10751 ), .DIN2(\IDinst/n10750 ), 
        .Q(\IDinst/n10752 ) );
  nnd2s1 \IDinst/U10820  ( .DIN1(\IDinst/n10749 ), .DIN2(n1379), 
        .Q(\IDinst/n10751 ) );
  nnd2s1 \IDinst/U10819  ( .DIN1(\IDinst/n10740 ), .DIN2(n1369), 
        .Q(\IDinst/n10750 ) );
  nnd2s1 \IDinst/U10818  ( .DIN1(\IDinst/n10748 ), .DIN2(\IDinst/n10747 ), 
        .Q(\IDinst/n10749 ) );
  nnd2s1 \IDinst/U10817  ( .DIN1(\IDinst/n10746 ), .DIN2(n1315), 
        .Q(\IDinst/n10748 ) );
  nnd2s1 \IDinst/U10816  ( .DIN1(\IDinst/n10743 ), .DIN2(n1358), 
        .Q(\IDinst/n10747 ) );
  nnd2s1 \IDinst/U10815  ( .DIN1(\IDinst/n10745 ), .DIN2(\IDinst/n10744 ), 
        .Q(\IDinst/n10746 ) );
  nnd2s1 \IDinst/U10814  ( .DIN1(\IDinst/RegFile[31][19] ), .DIN2(n1203), 
        .Q(\IDinst/n10745 ) );
  nnd2s1 \IDinst/U10813  ( .DIN1(\IDinst/RegFile[30][19] ), .DIN2(n1287), 
        .Q(\IDinst/n10744 ) );
  nnd2s1 \IDinst/U10812  ( .DIN1(\IDinst/n10742 ), .DIN2(\IDinst/n10741 ), 
        .Q(\IDinst/n10743 ) );
  nnd2s1 \IDinst/U10811  ( .DIN1(\IDinst/RegFile[29][19] ), .DIN2(n1203), 
        .Q(\IDinst/n10742 ) );
  nnd2s1 \IDinst/U10810  ( .DIN1(\IDinst/RegFile[28][19] ), .DIN2(n1287), 
        .Q(\IDinst/n10741 ) );
  nnd2s1 \IDinst/U10809  ( .DIN1(\IDinst/n10739 ), .DIN2(\IDinst/n10738 ), 
        .Q(\IDinst/n10740 ) );
  nnd2s1 \IDinst/U10808  ( .DIN1(\IDinst/n10737 ), .DIN2(n1314), 
        .Q(\IDinst/n10739 ) );
  nnd2s1 \IDinst/U10807  ( .DIN1(\IDinst/n10734 ), .DIN2(n1358), 
        .Q(\IDinst/n10738 ) );
  nnd2s1 \IDinst/U10806  ( .DIN1(\IDinst/n10736 ), .DIN2(\IDinst/n10735 ), 
        .Q(\IDinst/n10737 ) );
  nnd2s1 \IDinst/U10805  ( .DIN1(\IDinst/RegFile[27][19] ), .DIN2(n1203), 
        .Q(\IDinst/n10736 ) );
  nnd2s1 \IDinst/U10804  ( .DIN1(\IDinst/RegFile[26][19] ), .DIN2(n1287), 
        .Q(\IDinst/n10735 ) );
  nnd2s1 \IDinst/U10803  ( .DIN1(\IDinst/n10733 ), .DIN2(\IDinst/n10732 ), 
        .Q(\IDinst/n10734 ) );
  nnd2s1 \IDinst/U10802  ( .DIN1(\IDinst/RegFile[25][19] ), .DIN2(n1203), 
        .Q(\IDinst/n10733 ) );
  nnd2s1 \IDinst/U10801  ( .DIN1(\IDinst/RegFile[24][19] ), .DIN2(n1287), 
        .Q(\IDinst/n10732 ) );
  nnd2s1 \IDinst/U10800  ( .DIN1(\IDinst/n10730 ), .DIN2(\IDinst/n10729 ), 
        .Q(\IDinst/n10731 ) );
  nnd2s1 \IDinst/U10799  ( .DIN1(\IDinst/n10728 ), .DIN2(n1375), 
        .Q(\IDinst/n10730 ) );
  nnd2s1 \IDinst/U10798  ( .DIN1(\IDinst/n10719 ), .DIN2(n1369), 
        .Q(\IDinst/n10729 ) );
  nnd2s1 \IDinst/U10797  ( .DIN1(\IDinst/n10727 ), .DIN2(\IDinst/n10726 ), 
        .Q(\IDinst/n10728 ) );
  nnd2s1 \IDinst/U10796  ( .DIN1(\IDinst/n10725 ), .DIN2(n1314), 
        .Q(\IDinst/n10727 ) );
  nnd2s1 \IDinst/U10795  ( .DIN1(\IDinst/n10722 ), .DIN2(n1358), 
        .Q(\IDinst/n10726 ) );
  nnd2s1 \IDinst/U10794  ( .DIN1(\IDinst/n10724 ), .DIN2(\IDinst/n10723 ), 
        .Q(\IDinst/n10725 ) );
  nnd2s1 \IDinst/U10793  ( .DIN1(\IDinst/RegFile[23][19] ), .DIN2(n1203), 
        .Q(\IDinst/n10724 ) );
  nnd2s1 \IDinst/U10792  ( .DIN1(\IDinst/RegFile[22][19] ), .DIN2(n1287), 
        .Q(\IDinst/n10723 ) );
  nnd2s1 \IDinst/U10791  ( .DIN1(\IDinst/n10721 ), .DIN2(\IDinst/n10720 ), 
        .Q(\IDinst/n10722 ) );
  nnd2s1 \IDinst/U10790  ( .DIN1(\IDinst/RegFile[21][19] ), .DIN2(n1204), 
        .Q(\IDinst/n10721 ) );
  nnd2s1 \IDinst/U10789  ( .DIN1(\IDinst/RegFile[20][19] ), .DIN2(n1286), 
        .Q(\IDinst/n10720 ) );
  nnd2s1 \IDinst/U10788  ( .DIN1(\IDinst/n10718 ), .DIN2(\IDinst/n10717 ), 
        .Q(\IDinst/n10719 ) );
  nnd2s1 \IDinst/U10787  ( .DIN1(\IDinst/n10716 ), .DIN2(n1314), 
        .Q(\IDinst/n10718 ) );
  nnd2s1 \IDinst/U10786  ( .DIN1(\IDinst/n10713 ), .DIN2(n1358), 
        .Q(\IDinst/n10717 ) );
  nnd2s1 \IDinst/U10785  ( .DIN1(\IDinst/n10715 ), .DIN2(\IDinst/n10714 ), 
        .Q(\IDinst/n10716 ) );
  nnd2s1 \IDinst/U10784  ( .DIN1(\IDinst/RegFile[19][19] ), .DIN2(n1204), 
        .Q(\IDinst/n10715 ) );
  nnd2s1 \IDinst/U10783  ( .DIN1(\IDinst/RegFile[18][19] ), .DIN2(n1286), 
        .Q(\IDinst/n10714 ) );
  nnd2s1 \IDinst/U10782  ( .DIN1(\IDinst/n10712 ), .DIN2(\IDinst/n10711 ), 
        .Q(\IDinst/n10713 ) );
  nnd2s1 \IDinst/U10781  ( .DIN1(\IDinst/RegFile[17][19] ), .DIN2(n1204), 
        .Q(\IDinst/n10712 ) );
  nnd2s1 \IDinst/U10780  ( .DIN1(\IDinst/RegFile[16][19] ), .DIN2(n1286), 
        .Q(\IDinst/n10711 ) );
  nnd2s1 \IDinst/U10779  ( .DIN1(\IDinst/n10709 ), .DIN2(\IDinst/n10708 ), 
        .Q(\IDinst/n10710 ) );
  nnd2s1 \IDinst/U10778  ( .DIN1(\IDinst/n10707 ), .DIN2(n665), 
        .Q(\IDinst/n10709 ) );
  nnd2s1 \IDinst/U10777  ( .DIN1(\IDinst/n10686 ), .DIN2(n682), 
        .Q(\IDinst/n10708 ) );
  nnd2s1 \IDinst/U10776  ( .DIN1(\IDinst/n10706 ), .DIN2(\IDinst/n10705 ), 
        .Q(\IDinst/n10707 ) );
  nnd2s1 \IDinst/U10775  ( .DIN1(\IDinst/n10704 ), .DIN2(n1373), 
        .Q(\IDinst/n10706 ) );
  nnd2s1 \IDinst/U10774  ( .DIN1(\IDinst/n10695 ), .DIN2(n1369), 
        .Q(\IDinst/n10705 ) );
  nnd2s1 \IDinst/U10773  ( .DIN1(\IDinst/n10703 ), .DIN2(\IDinst/n10702 ), 
        .Q(\IDinst/n10704 ) );
  nnd2s1 \IDinst/U10772  ( .DIN1(\IDinst/n10701 ), .DIN2(n1314), 
        .Q(\IDinst/n10703 ) );
  nnd2s1 \IDinst/U10771  ( .DIN1(\IDinst/n10698 ), .DIN2(n1358), 
        .Q(\IDinst/n10702 ) );
  nnd2s1 \IDinst/U10770  ( .DIN1(\IDinst/n10700 ), .DIN2(\IDinst/n10699 ), 
        .Q(\IDinst/n10701 ) );
  nnd2s1 \IDinst/U10769  ( .DIN1(\IDinst/RegFile[15][19] ), .DIN2(n1204), 
        .Q(\IDinst/n10700 ) );
  nnd2s1 \IDinst/U10768  ( .DIN1(\IDinst/RegFile[14][19] ), .DIN2(n1286), 
        .Q(\IDinst/n10699 ) );
  nnd2s1 \IDinst/U10767  ( .DIN1(\IDinst/n10697 ), .DIN2(\IDinst/n10696 ), 
        .Q(\IDinst/n10698 ) );
  nnd2s1 \IDinst/U10766  ( .DIN1(\IDinst/RegFile[13][19] ), .DIN2(n1204), 
        .Q(\IDinst/n10697 ) );
  nnd2s1 \IDinst/U10765  ( .DIN1(\IDinst/RegFile[12][19] ), .DIN2(n1286), 
        .Q(\IDinst/n10696 ) );
  nnd2s1 \IDinst/U10764  ( .DIN1(\IDinst/n10694 ), .DIN2(\IDinst/n10693 ), 
        .Q(\IDinst/n10695 ) );
  nnd2s1 \IDinst/U10763  ( .DIN1(\IDinst/n10692 ), .DIN2(n1314), 
        .Q(\IDinst/n10694 ) );
  nnd2s1 \IDinst/U10762  ( .DIN1(\IDinst/n10689 ), .DIN2(n1358), 
        .Q(\IDinst/n10693 ) );
  nnd2s1 \IDinst/U10761  ( .DIN1(\IDinst/n10691 ), .DIN2(\IDinst/n10690 ), 
        .Q(\IDinst/n10692 ) );
  nnd2s1 \IDinst/U10760  ( .DIN1(\IDinst/RegFile[11][19] ), .DIN2(n1204), 
        .Q(\IDinst/n10691 ) );
  nnd2s1 \IDinst/U10759  ( .DIN1(\IDinst/RegFile[10][19] ), .DIN2(n1286), 
        .Q(\IDinst/n10690 ) );
  nnd2s1 \IDinst/U10758  ( .DIN1(\IDinst/n10688 ), .DIN2(\IDinst/n10687 ), 
        .Q(\IDinst/n10689 ) );
  nnd2s1 \IDinst/U10757  ( .DIN1(\IDinst/RegFile[9][19] ), .DIN2(n1204), 
        .Q(\IDinst/n10688 ) );
  nnd2s1 \IDinst/U10756  ( .DIN1(\IDinst/RegFile[8][19] ), .DIN2(n1286), 
        .Q(\IDinst/n10687 ) );
  nnd2s1 \IDinst/U10755  ( .DIN1(\IDinst/n10685 ), .DIN2(\IDinst/n10684 ), 
        .Q(\IDinst/n10686 ) );
  nnd2s1 \IDinst/U10754  ( .DIN1(\IDinst/n10683 ), .DIN2(n1376), 
        .Q(\IDinst/n10685 ) );
  nnd2s1 \IDinst/U10753  ( .DIN1(\IDinst/n10674 ), .DIN2(n1369), 
        .Q(\IDinst/n10684 ) );
  nnd2s1 \IDinst/U10752  ( .DIN1(\IDinst/n10682 ), .DIN2(\IDinst/n10681 ), 
        .Q(\IDinst/n10683 ) );
  nnd2s1 \IDinst/U10751  ( .DIN1(\IDinst/n10680 ), .DIN2(n1314), 
        .Q(\IDinst/n10682 ) );
  nnd2s1 \IDinst/U10750  ( .DIN1(\IDinst/n10677 ), .DIN2(n1358), 
        .Q(\IDinst/n10681 ) );
  nnd2s1 \IDinst/U10749  ( .DIN1(\IDinst/n10679 ), .DIN2(\IDinst/n10678 ), 
        .Q(\IDinst/n10680 ) );
  nnd2s1 \IDinst/U10748  ( .DIN1(\IDinst/RegFile[7][19] ), .DIN2(n1204), 
        .Q(\IDinst/n10679 ) );
  nnd2s1 \IDinst/U10747  ( .DIN1(\IDinst/RegFile[6][19] ), .DIN2(n1286), 
        .Q(\IDinst/n10678 ) );
  nnd2s1 \IDinst/U10746  ( .DIN1(\IDinst/n10676 ), .DIN2(\IDinst/n10675 ), 
        .Q(\IDinst/n10677 ) );
  nnd2s1 \IDinst/U10745  ( .DIN1(\IDinst/RegFile[5][19] ), .DIN2(n1204), 
        .Q(\IDinst/n10676 ) );
  nnd2s1 \IDinst/U10744  ( .DIN1(\IDinst/RegFile[4][19] ), .DIN2(n1286), 
        .Q(\IDinst/n10675 ) );
  nnd2s1 \IDinst/U10743  ( .DIN1(\IDinst/n10673 ), .DIN2(\IDinst/n10672 ), 
        .Q(\IDinst/n10674 ) );
  nnd2s1 \IDinst/U10742  ( .DIN1(\IDinst/n10671 ), .DIN2(n1314), 
        .Q(\IDinst/n10673 ) );
  nnd2s1 \IDinst/U10741  ( .DIN1(\IDinst/n10668 ), .DIN2(n1358), 
        .Q(\IDinst/n10672 ) );
  nnd2s1 \IDinst/U10740  ( .DIN1(\IDinst/n10670 ), .DIN2(\IDinst/n10669 ), 
        .Q(\IDinst/n10671 ) );
  nnd2s1 \IDinst/U10739  ( .DIN1(\IDinst/RegFile[3][19] ), .DIN2(n1204), 
        .Q(\IDinst/n10670 ) );
  nnd2s1 \IDinst/U10738  ( .DIN1(\IDinst/RegFile[2][19] ), .DIN2(n1285), 
        .Q(\IDinst/n10669 ) );
  nnd2s1 \IDinst/U10737  ( .DIN1(\IDinst/n10667 ), .DIN2(\IDinst/n10666 ), 
        .Q(\IDinst/n10668 ) );
  nnd2s1 \IDinst/U10736  ( .DIN1(\IDinst/RegFile[1][19] ), .DIN2(n1204), 
        .Q(\IDinst/n10667 ) );
  nnd2s1 \IDinst/U10735  ( .DIN1(\IDinst/RegFile[0][19] ), .DIN2(n1285), 
        .Q(\IDinst/n10666 ) );
  nnd2s1 \IDinst/U10734  ( .DIN1(\IDinst/n10665 ), .DIN2(n535), 
        .Q(\IDinst/n8928 ) );
  nnd2s1 \IDinst/U10733  ( .DIN1(\IDinst/n10620 ), .DIN2(n634), 
        .Q(\IDinst/n8929 ) );
  nnd2s1 \IDinst/U10732  ( .DIN1(\IDinst/n10664 ), .DIN2(\IDinst/n10663 ), 
        .Q(\IDinst/n10665 ) );
  nnd2s1 \IDinst/U10731  ( .DIN1(\IDinst/n10662 ), .DIN2(n668), 
        .Q(\IDinst/n10664 ) );
  nnd2s1 \IDinst/U10730  ( .DIN1(\IDinst/n10641 ), .DIN2(n680), 
        .Q(\IDinst/n10663 ) );
  nnd2s1 \IDinst/U10729  ( .DIN1(\IDinst/n10661 ), .DIN2(\IDinst/n10660 ), 
        .Q(\IDinst/n10662 ) );
  nnd2s1 \IDinst/U10728  ( .DIN1(\IDinst/n10659 ), .DIN2(n1377), 
        .Q(\IDinst/n10661 ) );
  nnd2s1 \IDinst/U10727  ( .DIN1(\IDinst/n10650 ), .DIN2(n1369), 
        .Q(\IDinst/n10660 ) );
  nnd2s1 \IDinst/U10726  ( .DIN1(\IDinst/n10658 ), .DIN2(\IDinst/n10657 ), 
        .Q(\IDinst/n10659 ) );
  nnd2s1 \IDinst/U10725  ( .DIN1(\IDinst/n10656 ), .DIN2(n1314), 
        .Q(\IDinst/n10658 ) );
  nnd2s1 \IDinst/U10724  ( .DIN1(\IDinst/n10653 ), .DIN2(n1359), 
        .Q(\IDinst/n10657 ) );
  nnd2s1 \IDinst/U10723  ( .DIN1(\IDinst/n10655 ), .DIN2(\IDinst/n10654 ), 
        .Q(\IDinst/n10656 ) );
  nnd2s1 \IDinst/U10722  ( .DIN1(\IDinst/RegFile[31][18] ), .DIN2(n1204), 
        .Q(\IDinst/n10655 ) );
  nnd2s1 \IDinst/U10721  ( .DIN1(\IDinst/RegFile[30][18] ), .DIN2(n1285), 
        .Q(\IDinst/n10654 ) );
  nnd2s1 \IDinst/U10720  ( .DIN1(\IDinst/n10652 ), .DIN2(\IDinst/n10651 ), 
        .Q(\IDinst/n10653 ) );
  nnd2s1 \IDinst/U10719  ( .DIN1(\IDinst/RegFile[29][18] ), .DIN2(n1204), 
        .Q(\IDinst/n10652 ) );
  nnd2s1 \IDinst/U10718  ( .DIN1(\IDinst/RegFile[28][18] ), .DIN2(n1285), 
        .Q(\IDinst/n10651 ) );
  nnd2s1 \IDinst/U10717  ( .DIN1(\IDinst/n10649 ), .DIN2(\IDinst/n10648 ), 
        .Q(\IDinst/n10650 ) );
  nnd2s1 \IDinst/U10716  ( .DIN1(\IDinst/n10647 ), .DIN2(n1314), 
        .Q(\IDinst/n10649 ) );
  nnd2s1 \IDinst/U10715  ( .DIN1(\IDinst/n10644 ), .DIN2(n1359), 
        .Q(\IDinst/n10648 ) );
  nnd2s1 \IDinst/U10714  ( .DIN1(\IDinst/n10646 ), .DIN2(\IDinst/n10645 ), 
        .Q(\IDinst/n10647 ) );
  nnd2s1 \IDinst/U10713  ( .DIN1(\IDinst/RegFile[27][18] ), .DIN2(n1205), 
        .Q(\IDinst/n10646 ) );
  nnd2s1 \IDinst/U10712  ( .DIN1(\IDinst/RegFile[26][18] ), .DIN2(n1285), 
        .Q(\IDinst/n10645 ) );
  nnd2s1 \IDinst/U10711  ( .DIN1(\IDinst/n10643 ), .DIN2(\IDinst/n10642 ), 
        .Q(\IDinst/n10644 ) );
  nnd2s1 \IDinst/U10710  ( .DIN1(\IDinst/RegFile[25][18] ), .DIN2(n1205), 
        .Q(\IDinst/n10643 ) );
  nnd2s1 \IDinst/U10709  ( .DIN1(\IDinst/RegFile[24][18] ), .DIN2(n1285), 
        .Q(\IDinst/n10642 ) );
  nnd2s1 \IDinst/U10708  ( .DIN1(\IDinst/n10640 ), .DIN2(\IDinst/n10639 ), 
        .Q(\IDinst/n10641 ) );
  nnd2s1 \IDinst/U10707  ( .DIN1(\IDinst/n10638 ), .DIN2(n1380), 
        .Q(\IDinst/n10640 ) );
  nnd2s1 \IDinst/U10706  ( .DIN1(\IDinst/n10629 ), .DIN2(n1369), 
        .Q(\IDinst/n10639 ) );
  nnd2s1 \IDinst/U10705  ( .DIN1(\IDinst/n10637 ), .DIN2(\IDinst/n10636 ), 
        .Q(\IDinst/n10638 ) );
  nnd2s1 \IDinst/U10704  ( .DIN1(\IDinst/n10635 ), .DIN2(n1314), 
        .Q(\IDinst/n10637 ) );
  nnd2s1 \IDinst/U10703  ( .DIN1(\IDinst/n10632 ), .DIN2(n1359), 
        .Q(\IDinst/n10636 ) );
  nnd2s1 \IDinst/U10702  ( .DIN1(\IDinst/n10634 ), .DIN2(\IDinst/n10633 ), 
        .Q(\IDinst/n10635 ) );
  nnd2s1 \IDinst/U10701  ( .DIN1(\IDinst/RegFile[23][18] ), .DIN2(n1205), 
        .Q(\IDinst/n10634 ) );
  nnd2s1 \IDinst/U10700  ( .DIN1(\IDinst/RegFile[22][18] ), .DIN2(n1285), 
        .Q(\IDinst/n10633 ) );
  nnd2s1 \IDinst/U10699  ( .DIN1(\IDinst/n10631 ), .DIN2(\IDinst/n10630 ), 
        .Q(\IDinst/n10632 ) );
  nnd2s1 \IDinst/U10698  ( .DIN1(\IDinst/RegFile[21][18] ), .DIN2(n1205), 
        .Q(\IDinst/n10631 ) );
  nnd2s1 \IDinst/U10697  ( .DIN1(\IDinst/RegFile[20][18] ), .DIN2(n1285), 
        .Q(\IDinst/n10630 ) );
  nnd2s1 \IDinst/U10696  ( .DIN1(\IDinst/n10628 ), .DIN2(\IDinst/n10627 ), 
        .Q(\IDinst/n10629 ) );
  nnd2s1 \IDinst/U10695  ( .DIN1(\IDinst/n10626 ), .DIN2(n1314), 
        .Q(\IDinst/n10628 ) );
  nnd2s1 \IDinst/U10694  ( .DIN1(\IDinst/n10623 ), .DIN2(n1359), 
        .Q(\IDinst/n10627 ) );
  nnd2s1 \IDinst/U10693  ( .DIN1(\IDinst/n10625 ), .DIN2(\IDinst/n10624 ), 
        .Q(\IDinst/n10626 ) );
  nnd2s1 \IDinst/U10692  ( .DIN1(\IDinst/RegFile[19][18] ), .DIN2(n1205), 
        .Q(\IDinst/n10625 ) );
  nnd2s1 \IDinst/U10691  ( .DIN1(\IDinst/RegFile[18][18] ), .DIN2(n1285), 
        .Q(\IDinst/n10624 ) );
  nnd2s1 \IDinst/U10690  ( .DIN1(\IDinst/n10622 ), .DIN2(\IDinst/n10621 ), 
        .Q(\IDinst/n10623 ) );
  nnd2s1 \IDinst/U10689  ( .DIN1(\IDinst/RegFile[17][18] ), .DIN2(n1205), 
        .Q(\IDinst/n10622 ) );
  nnd2s1 \IDinst/U10688  ( .DIN1(\IDinst/RegFile[16][18] ), .DIN2(n1284), 
        .Q(\IDinst/n10621 ) );
  nnd2s1 \IDinst/U10687  ( .DIN1(\IDinst/n10619 ), .DIN2(\IDinst/n10618 ), 
        .Q(\IDinst/n10620 ) );
  nnd2s1 \IDinst/U10686  ( .DIN1(\IDinst/n10617 ), .DIN2(n666), 
        .Q(\IDinst/n10619 ) );
  nnd2s1 \IDinst/U10685  ( .DIN1(\IDinst/n10596 ), .DIN2(n681), 
        .Q(\IDinst/n10618 ) );
  nnd2s1 \IDinst/U10684  ( .DIN1(\IDinst/n10616 ), .DIN2(\IDinst/n10615 ), 
        .Q(\IDinst/n10617 ) );
  nnd2s1 \IDinst/U10683  ( .DIN1(\IDinst/n10614 ), .DIN2(n1374), 
        .Q(\IDinst/n10616 ) );
  nnd2s1 \IDinst/U10682  ( .DIN1(\IDinst/n10605 ), .DIN2(n1369), 
        .Q(\IDinst/n10615 ) );
  nnd2s1 \IDinst/U10681  ( .DIN1(\IDinst/n10613 ), .DIN2(\IDinst/n10612 ), 
        .Q(\IDinst/n10614 ) );
  nnd2s1 \IDinst/U10680  ( .DIN1(\IDinst/n10611 ), .DIN2(n1314), 
        .Q(\IDinst/n10613 ) );
  nnd2s1 \IDinst/U10679  ( .DIN1(\IDinst/n10608 ), .DIN2(n1359), 
        .Q(\IDinst/n10612 ) );
  nnd2s1 \IDinst/U10678  ( .DIN1(\IDinst/n10610 ), .DIN2(\IDinst/n10609 ), 
        .Q(\IDinst/n10611 ) );
  nnd2s1 \IDinst/U10677  ( .DIN1(\IDinst/RegFile[15][18] ), .DIN2(n1205), 
        .Q(\IDinst/n10610 ) );
  nnd2s1 \IDinst/U10676  ( .DIN1(\IDinst/RegFile[14][18] ), .DIN2(n1284), 
        .Q(\IDinst/n10609 ) );
  nnd2s1 \IDinst/U10675  ( .DIN1(\IDinst/n10607 ), .DIN2(\IDinst/n10606 ), 
        .Q(\IDinst/n10608 ) );
  nnd2s1 \IDinst/U10674  ( .DIN1(\IDinst/RegFile[13][18] ), .DIN2(n1205), 
        .Q(\IDinst/n10607 ) );
  nnd2s1 \IDinst/U10673  ( .DIN1(\IDinst/RegFile[12][18] ), .DIN2(n1284), 
        .Q(\IDinst/n10606 ) );
  nnd2s1 \IDinst/U10672  ( .DIN1(\IDinst/n10604 ), .DIN2(\IDinst/n10603 ), 
        .Q(\IDinst/n10605 ) );
  nnd2s1 \IDinst/U10671  ( .DIN1(\IDinst/n10602 ), .DIN2(n1314), 
        .Q(\IDinst/n10604 ) );
  nnd2s1 \IDinst/U10670  ( .DIN1(\IDinst/n10599 ), .DIN2(n1359), 
        .Q(\IDinst/n10603 ) );
  nnd2s1 \IDinst/U10669  ( .DIN1(\IDinst/n10601 ), .DIN2(\IDinst/n10600 ), 
        .Q(\IDinst/n10602 ) );
  nnd2s1 \IDinst/U10668  ( .DIN1(\IDinst/RegFile[11][18] ), .DIN2(n1205), 
        .Q(\IDinst/n10601 ) );
  nnd2s1 \IDinst/U10667  ( .DIN1(\IDinst/RegFile[10][18] ), .DIN2(n1284), 
        .Q(\IDinst/n10600 ) );
  nnd2s1 \IDinst/U10666  ( .DIN1(\IDinst/n10598 ), .DIN2(\IDinst/n10597 ), 
        .Q(\IDinst/n10599 ) );
  nnd2s1 \IDinst/U10665  ( .DIN1(\IDinst/RegFile[9][18] ), .DIN2(n1205), 
        .Q(\IDinst/n10598 ) );
  nnd2s1 \IDinst/U10664  ( .DIN1(\IDinst/RegFile[8][18] ), .DIN2(n1284), 
        .Q(\IDinst/n10597 ) );
  nnd2s1 \IDinst/U10663  ( .DIN1(\IDinst/n10595 ), .DIN2(\IDinst/n10594 ), 
        .Q(\IDinst/n10596 ) );
  nnd2s1 \IDinst/U10662  ( .DIN1(\IDinst/n10593 ), .DIN2(n1374), 
        .Q(\IDinst/n10595 ) );
  nnd2s1 \IDinst/U10661  ( .DIN1(\IDinst/n10584 ), .DIN2(n1369), 
        .Q(\IDinst/n10594 ) );
  nnd2s1 \IDinst/U10660  ( .DIN1(\IDinst/n10592 ), .DIN2(\IDinst/n10591 ), 
        .Q(\IDinst/n10593 ) );
  nnd2s1 \IDinst/U10659  ( .DIN1(\IDinst/n10590 ), .DIN2(n1313), 
        .Q(\IDinst/n10592 ) );
  nnd2s1 \IDinst/U10658  ( .DIN1(\IDinst/n10587 ), .DIN2(n1359), 
        .Q(\IDinst/n10591 ) );
  nnd2s1 \IDinst/U10657  ( .DIN1(\IDinst/n10589 ), .DIN2(\IDinst/n10588 ), 
        .Q(\IDinst/n10590 ) );
  nnd2s1 \IDinst/U10656  ( .DIN1(\IDinst/RegFile[7][18] ), .DIN2(n1205), 
        .Q(\IDinst/n10589 ) );
  nnd2s1 \IDinst/U10655  ( .DIN1(\IDinst/RegFile[6][18] ), .DIN2(n1284), 
        .Q(\IDinst/n10588 ) );
  nnd2s1 \IDinst/U10654  ( .DIN1(\IDinst/n10586 ), .DIN2(\IDinst/n10585 ), 
        .Q(\IDinst/n10587 ) );
  nnd2s1 \IDinst/U10653  ( .DIN1(\IDinst/RegFile[5][18] ), .DIN2(n1205), 
        .Q(\IDinst/n10586 ) );
  nnd2s1 \IDinst/U10652  ( .DIN1(\IDinst/RegFile[4][18] ), .DIN2(n1284), 
        .Q(\IDinst/n10585 ) );
  nnd2s1 \IDinst/U10651  ( .DIN1(\IDinst/n10583 ), .DIN2(\IDinst/n10582 ), 
        .Q(\IDinst/n10584 ) );
  nnd2s1 \IDinst/U10650  ( .DIN1(\IDinst/n10581 ), .DIN2(n1313), 
        .Q(\IDinst/n10583 ) );
  nnd2s1 \IDinst/U10649  ( .DIN1(\IDinst/n10578 ), .DIN2(n1359), 
        .Q(\IDinst/n10582 ) );
  nnd2s1 \IDinst/U10648  ( .DIN1(\IDinst/n10580 ), .DIN2(\IDinst/n10579 ), 
        .Q(\IDinst/n10581 ) );
  nnd2s1 \IDinst/U10647  ( .DIN1(\IDinst/RegFile[3][18] ), .DIN2(n1205), 
        .Q(\IDinst/n10580 ) );
  nnd2s1 \IDinst/U10646  ( .DIN1(\IDinst/RegFile[2][18] ), .DIN2(n1284), 
        .Q(\IDinst/n10579 ) );
  nnd2s1 \IDinst/U10645  ( .DIN1(\IDinst/n10577 ), .DIN2(\IDinst/n10576 ), 
        .Q(\IDinst/n10578 ) );
  nnd2s1 \IDinst/U10644  ( .DIN1(\IDinst/RegFile[1][18] ), .DIN2(n1206), 
        .Q(\IDinst/n10577 ) );
  nnd2s1 \IDinst/U10643  ( .DIN1(\IDinst/RegFile[0][18] ), .DIN2(n1284), 
        .Q(\IDinst/n10576 ) );
  nnd2s1 \IDinst/U10642  ( .DIN1(\IDinst/n10575 ), .DIN2(n534), 
        .Q(\IDinst/n8926 ) );
  nnd2s1 \IDinst/U10641  ( .DIN1(\IDinst/n10530 ), .DIN2(n533), 
        .Q(\IDinst/n8927 ) );
  nnd2s1 \IDinst/U10640  ( .DIN1(\IDinst/n10574 ), .DIN2(\IDinst/n10573 ), 
        .Q(\IDinst/n10575 ) );
  nnd2s1 \IDinst/U10639  ( .DIN1(\IDinst/n10572 ), .DIN2(n667), 
        .Q(\IDinst/n10574 ) );
  nnd2s1 \IDinst/U10638  ( .DIN1(\IDinst/n10551 ), .DIN2(n683), 
        .Q(\IDinst/n10573 ) );
  nnd2s1 \IDinst/U10637  ( .DIN1(\IDinst/n10571 ), .DIN2(\IDinst/n10570 ), 
        .Q(\IDinst/n10572 ) );
  nnd2s1 \IDinst/U10636  ( .DIN1(\IDinst/n10569 ), .DIN2(n1374), 
        .Q(\IDinst/n10571 ) );
  nnd2s1 \IDinst/U10635  ( .DIN1(\IDinst/n10560 ), .DIN2(n1369), 
        .Q(\IDinst/n10570 ) );
  nnd2s1 \IDinst/U10634  ( .DIN1(\IDinst/n10568 ), .DIN2(\IDinst/n10567 ), 
        .Q(\IDinst/n10569 ) );
  nnd2s1 \IDinst/U10633  ( .DIN1(\IDinst/n10566 ), .DIN2(n1313), 
        .Q(\IDinst/n10568 ) );
  nnd2s1 \IDinst/U10632  ( .DIN1(\IDinst/n10563 ), .DIN2(n1359), 
        .Q(\IDinst/n10567 ) );
  nnd2s1 \IDinst/U10631  ( .DIN1(\IDinst/n10565 ), .DIN2(\IDinst/n10564 ), 
        .Q(\IDinst/n10566 ) );
  nnd2s1 \IDinst/U10630  ( .DIN1(\IDinst/RegFile[31][17] ), .DIN2(n1206), 
        .Q(\IDinst/n10565 ) );
  nnd2s1 \IDinst/U10629  ( .DIN1(\IDinst/RegFile[30][17] ), .DIN2(n1283), 
        .Q(\IDinst/n10564 ) );
  nnd2s1 \IDinst/U10628  ( .DIN1(\IDinst/n10562 ), .DIN2(\IDinst/n10561 ), 
        .Q(\IDinst/n10563 ) );
  nnd2s1 \IDinst/U10627  ( .DIN1(\IDinst/RegFile[29][17] ), .DIN2(n1206), 
        .Q(\IDinst/n10562 ) );
  nnd2s1 \IDinst/U10626  ( .DIN1(\IDinst/RegFile[28][17] ), .DIN2(n1283), 
        .Q(\IDinst/n10561 ) );
  nnd2s1 \IDinst/U10625  ( .DIN1(\IDinst/n10559 ), .DIN2(\IDinst/n10558 ), 
        .Q(\IDinst/n10560 ) );
  nnd2s1 \IDinst/U10624  ( .DIN1(\IDinst/n10557 ), .DIN2(n1313), 
        .Q(\IDinst/n10559 ) );
  nnd2s1 \IDinst/U10623  ( .DIN1(\IDinst/n10554 ), .DIN2(n1360), 
        .Q(\IDinst/n10558 ) );
  nnd2s1 \IDinst/U10622  ( .DIN1(\IDinst/n10556 ), .DIN2(\IDinst/n10555 ), 
        .Q(\IDinst/n10557 ) );
  nnd2s1 \IDinst/U10621  ( .DIN1(\IDinst/RegFile[27][17] ), .DIN2(n1206), 
        .Q(\IDinst/n10556 ) );
  nnd2s1 \IDinst/U10620  ( .DIN1(\IDinst/RegFile[26][17] ), .DIN2(n1283), 
        .Q(\IDinst/n10555 ) );
  nnd2s1 \IDinst/U10619  ( .DIN1(\IDinst/n10553 ), .DIN2(\IDinst/n10552 ), 
        .Q(\IDinst/n10554 ) );
  nnd2s1 \IDinst/U10618  ( .DIN1(\IDinst/RegFile[25][17] ), .DIN2(n1206), 
        .Q(\IDinst/n10553 ) );
  nnd2s1 \IDinst/U10617  ( .DIN1(\IDinst/RegFile[24][17] ), .DIN2(n1283), 
        .Q(\IDinst/n10552 ) );
  nnd2s1 \IDinst/U10616  ( .DIN1(\IDinst/n10550 ), .DIN2(\IDinst/n10549 ), 
        .Q(\IDinst/n10551 ) );
  nnd2s1 \IDinst/U10615  ( .DIN1(\IDinst/n10548 ), .DIN2(n1374), 
        .Q(\IDinst/n10550 ) );
  nnd2s1 \IDinst/U10614  ( .DIN1(\IDinst/n10539 ), .DIN2(n1369), 
        .Q(\IDinst/n10549 ) );
  nnd2s1 \IDinst/U10613  ( .DIN1(\IDinst/n10547 ), .DIN2(\IDinst/n10546 ), 
        .Q(\IDinst/n10548 ) );
  nnd2s1 \IDinst/U10612  ( .DIN1(\IDinst/n10545 ), .DIN2(n1313), 
        .Q(\IDinst/n10547 ) );
  nnd2s1 \IDinst/U10611  ( .DIN1(\IDinst/n10542 ), .DIN2(n1360), 
        .Q(\IDinst/n10546 ) );
  nnd2s1 \IDinst/U10610  ( .DIN1(\IDinst/n10544 ), .DIN2(\IDinst/n10543 ), 
        .Q(\IDinst/n10545 ) );
  nnd2s1 \IDinst/U10609  ( .DIN1(\IDinst/RegFile[23][17] ), .DIN2(n1206), 
        .Q(\IDinst/n10544 ) );
  nnd2s1 \IDinst/U10608  ( .DIN1(\IDinst/RegFile[22][17] ), .DIN2(n1283), 
        .Q(\IDinst/n10543 ) );
  nnd2s1 \IDinst/U10607  ( .DIN1(\IDinst/n10541 ), .DIN2(\IDinst/n10540 ), 
        .Q(\IDinst/n10542 ) );
  nnd2s1 \IDinst/U10606  ( .DIN1(\IDinst/RegFile[21][17] ), .DIN2(n1206), 
        .Q(\IDinst/n10541 ) );
  nnd2s1 \IDinst/U10605  ( .DIN1(\IDinst/RegFile[20][17] ), .DIN2(n1283), 
        .Q(\IDinst/n10540 ) );
  nnd2s1 \IDinst/U10604  ( .DIN1(\IDinst/n10538 ), .DIN2(\IDinst/n10537 ), 
        .Q(\IDinst/n10539 ) );
  nnd2s1 \IDinst/U10603  ( .DIN1(\IDinst/n10536 ), .DIN2(n1313), 
        .Q(\IDinst/n10538 ) );
  nnd2s1 \IDinst/U10602  ( .DIN1(\IDinst/n10533 ), .DIN2(n1360), 
        .Q(\IDinst/n10537 ) );
  nnd2s1 \IDinst/U10601  ( .DIN1(\IDinst/n10535 ), .DIN2(\IDinst/n10534 ), 
        .Q(\IDinst/n10536 ) );
  nnd2s1 \IDinst/U10600  ( .DIN1(\IDinst/RegFile[19][17] ), .DIN2(n1206), 
        .Q(\IDinst/n10535 ) );
  nnd2s1 \IDinst/U10599  ( .DIN1(\IDinst/RegFile[18][17] ), .DIN2(n1283), 
        .Q(\IDinst/n10534 ) );
  nnd2s1 \IDinst/U10598  ( .DIN1(\IDinst/n10532 ), .DIN2(\IDinst/n10531 ), 
        .Q(\IDinst/n10533 ) );
  nnd2s1 \IDinst/U10597  ( .DIN1(\IDinst/RegFile[17][17] ), .DIN2(n1206), 
        .Q(\IDinst/n10532 ) );
  nnd2s1 \IDinst/U10596  ( .DIN1(\IDinst/RegFile[16][17] ), .DIN2(n1283), 
        .Q(\IDinst/n10531 ) );
  nnd2s1 \IDinst/U10595  ( .DIN1(\IDinst/n10529 ), .DIN2(\IDinst/n10528 ), 
        .Q(\IDinst/n10530 ) );
  nnd2s1 \IDinst/U10594  ( .DIN1(\IDinst/n10527 ), .DIN2(n665), 
        .Q(\IDinst/n10529 ) );
  nnd2s1 \IDinst/U10593  ( .DIN1(\IDinst/n10506 ), .DIN2(n682), 
        .Q(\IDinst/n10528 ) );
  nnd2s1 \IDinst/U10592  ( .DIN1(\IDinst/n10526 ), .DIN2(\IDinst/n10525 ), 
        .Q(\IDinst/n10527 ) );
  nnd2s1 \IDinst/U10591  ( .DIN1(\IDinst/n10524 ), .DIN2(n1374), 
        .Q(\IDinst/n10526 ) );
  nnd2s1 \IDinst/U10590  ( .DIN1(\IDinst/n10515 ), .DIN2(n1369), 
        .Q(\IDinst/n10525 ) );
  nnd2s1 \IDinst/U10589  ( .DIN1(\IDinst/n10523 ), .DIN2(\IDinst/n10522 ), 
        .Q(\IDinst/n10524 ) );
  nnd2s1 \IDinst/U10588  ( .DIN1(\IDinst/n10521 ), .DIN2(n1313), 
        .Q(\IDinst/n10523 ) );
  nnd2s1 \IDinst/U10587  ( .DIN1(\IDinst/n10518 ), .DIN2(n1360), 
        .Q(\IDinst/n10522 ) );
  nnd2s1 \IDinst/U10586  ( .DIN1(\IDinst/n10520 ), .DIN2(\IDinst/n10519 ), 
        .Q(\IDinst/n10521 ) );
  nnd2s1 \IDinst/U10585  ( .DIN1(\IDinst/RegFile[15][17] ), .DIN2(n1206), 
        .Q(\IDinst/n10520 ) );
  nnd2s1 \IDinst/U10584  ( .DIN1(\IDinst/RegFile[14][17] ), .DIN2(n1283), 
        .Q(\IDinst/n10519 ) );
  nnd2s1 \IDinst/U10583  ( .DIN1(\IDinst/n10517 ), .DIN2(\IDinst/n10516 ), 
        .Q(\IDinst/n10518 ) );
  nnd2s1 \IDinst/U10582  ( .DIN1(\IDinst/RegFile[13][17] ), .DIN2(n1206), 
        .Q(\IDinst/n10517 ) );
  nnd2s1 \IDinst/U10581  ( .DIN1(\IDinst/RegFile[12][17] ), .DIN2(n1282), 
        .Q(\IDinst/n10516 ) );
  nnd2s1 \IDinst/U10580  ( .DIN1(\IDinst/n10514 ), .DIN2(\IDinst/n10513 ), 
        .Q(\IDinst/n10515 ) );
  nnd2s1 \IDinst/U10579  ( .DIN1(\IDinst/n10512 ), .DIN2(n1313), 
        .Q(\IDinst/n10514 ) );
  nnd2s1 \IDinst/U10578  ( .DIN1(\IDinst/n10509 ), .DIN2(n1340), 
        .Q(\IDinst/n10513 ) );
  nnd2s1 \IDinst/U10577  ( .DIN1(\IDinst/n10511 ), .DIN2(\IDinst/n10510 ), 
        .Q(\IDinst/n10512 ) );
  nnd2s1 \IDinst/U10576  ( .DIN1(\IDinst/RegFile[11][17] ), .DIN2(n1206), 
        .Q(\IDinst/n10511 ) );
  nnd2s1 \IDinst/U10575  ( .DIN1(\IDinst/RegFile[10][17] ), .DIN2(n1282), 
        .Q(\IDinst/n10510 ) );
  nnd2s1 \IDinst/U10574  ( .DIN1(\IDinst/n10508 ), .DIN2(\IDinst/n10507 ), 
        .Q(\IDinst/n10509 ) );
  nnd2s1 \IDinst/U10573  ( .DIN1(\IDinst/RegFile[9][17] ), .DIN2(n1206), 
        .Q(\IDinst/n10508 ) );
  nnd2s1 \IDinst/U10572  ( .DIN1(\IDinst/RegFile[8][17] ), .DIN2(n1282), 
        .Q(\IDinst/n10507 ) );
  nnd2s1 \IDinst/U10571  ( .DIN1(\IDinst/n10505 ), .DIN2(\IDinst/n10504 ), 
        .Q(\IDinst/n10506 ) );
  nnd2s1 \IDinst/U10570  ( .DIN1(\IDinst/n10503 ), .DIN2(n1374), 
        .Q(\IDinst/n10505 ) );
  nnd2s1 \IDinst/U10569  ( .DIN1(\IDinst/n10494 ), .DIN2(n1369), 
        .Q(\IDinst/n10504 ) );
  nnd2s1 \IDinst/U10568  ( .DIN1(\IDinst/n10502 ), .DIN2(\IDinst/n10501 ), 
        .Q(\IDinst/n10503 ) );
  nnd2s1 \IDinst/U10567  ( .DIN1(\IDinst/n10500 ), .DIN2(n1313), 
        .Q(\IDinst/n10502 ) );
  nnd2s1 \IDinst/U10566  ( .DIN1(\IDinst/n10497 ), .DIN2(n1333), 
        .Q(\IDinst/n10501 ) );
  nnd2s1 \IDinst/U10565  ( .DIN1(\IDinst/n10499 ), .DIN2(\IDinst/n10498 ), 
        .Q(\IDinst/n10500 ) );
  nnd2s1 \IDinst/U10564  ( .DIN1(\IDinst/RegFile[7][17] ), .DIN2(n1207), 
        .Q(\IDinst/n10499 ) );
  nnd2s1 \IDinst/U10563  ( .DIN1(\IDinst/RegFile[6][17] ), .DIN2(n1254), 
        .Q(\IDinst/n10498 ) );
  nnd2s1 \IDinst/U10562  ( .DIN1(\IDinst/n10496 ), .DIN2(\IDinst/n10495 ), 
        .Q(\IDinst/n10497 ) );
  nnd2s1 \IDinst/U10561  ( .DIN1(\IDinst/RegFile[5][17] ), .DIN2(n1207), 
        .Q(\IDinst/n10496 ) );
  nnd2s1 \IDinst/U10560  ( .DIN1(\IDinst/RegFile[4][17] ), .DIN2(n1254), 
        .Q(\IDinst/n10495 ) );
  nnd2s1 \IDinst/U10559  ( .DIN1(\IDinst/n10493 ), .DIN2(\IDinst/n10492 ), 
        .Q(\IDinst/n10494 ) );
  nnd2s1 \IDinst/U10558  ( .DIN1(\IDinst/n10491 ), .DIN2(n1313), 
        .Q(\IDinst/n10493 ) );
  nnd2s1 \IDinst/U10557  ( .DIN1(\IDinst/n10488 ), .DIN2(n1333), 
        .Q(\IDinst/n10492 ) );
  nnd2s1 \IDinst/U10556  ( .DIN1(\IDinst/n10490 ), .DIN2(\IDinst/n10489 ), 
        .Q(\IDinst/n10491 ) );
  nnd2s1 \IDinst/U10555  ( .DIN1(\IDinst/RegFile[3][17] ), .DIN2(n1207), 
        .Q(\IDinst/n10490 ) );
  nnd2s1 \IDinst/U10554  ( .DIN1(\IDinst/RegFile[2][17] ), .DIN2(n1254), 
        .Q(\IDinst/n10489 ) );
  nnd2s1 \IDinst/U10553  ( .DIN1(\IDinst/n10487 ), .DIN2(\IDinst/n10486 ), 
        .Q(\IDinst/n10488 ) );
  nnd2s1 \IDinst/U10552  ( .DIN1(\IDinst/RegFile[1][17] ), .DIN2(n1207), 
        .Q(\IDinst/n10487 ) );
  nnd2s1 \IDinst/U10551  ( .DIN1(\IDinst/RegFile[0][17] ), .DIN2(n1253), 
        .Q(\IDinst/n10486 ) );
  nnd2s1 \IDinst/U10550  ( .DIN1(\IDinst/n10485 ), .DIN2(\IDinst/N48 ), 
        .Q(\IDinst/n8924 ) );
  nnd2s1 \IDinst/U10549  ( .DIN1(\IDinst/n10440 ), .DIN2(n634), 
        .Q(\IDinst/n8925 ) );
  nnd2s1 \IDinst/U10548  ( .DIN1(\IDinst/n10484 ), .DIN2(\IDinst/n10483 ), 
        .Q(\IDinst/n10485 ) );
  nnd2s1 \IDinst/U10547  ( .DIN1(\IDinst/n10482 ), .DIN2(n668), 
        .Q(\IDinst/n10484 ) );
  nnd2s1 \IDinst/U10546  ( .DIN1(\IDinst/n10461 ), .DIN2(n680), 
        .Q(\IDinst/n10483 ) );
  nnd2s1 \IDinst/U10545  ( .DIN1(\IDinst/n10481 ), .DIN2(\IDinst/n10480 ), 
        .Q(\IDinst/n10482 ) );
  nnd2s1 \IDinst/U10544  ( .DIN1(\IDinst/n10479 ), .DIN2(n1374), 
        .Q(\IDinst/n10481 ) );
  nnd2s1 \IDinst/U10543  ( .DIN1(\IDinst/n10470 ), .DIN2(n1368), 
        .Q(\IDinst/n10480 ) );
  nnd2s1 \IDinst/U10542  ( .DIN1(\IDinst/n10478 ), .DIN2(\IDinst/n10477 ), 
        .Q(\IDinst/n10479 ) );
  nnd2s1 \IDinst/U10541  ( .DIN1(\IDinst/n10476 ), .DIN2(n1313), 
        .Q(\IDinst/n10478 ) );
  nnd2s1 \IDinst/U10540  ( .DIN1(\IDinst/n10473 ), .DIN2(n1333), 
        .Q(\IDinst/n10477 ) );
  nnd2s1 \IDinst/U10539  ( .DIN1(\IDinst/n10475 ), .DIN2(\IDinst/n10474 ), 
        .Q(\IDinst/n10476 ) );
  nnd2s1 \IDinst/U10538  ( .DIN1(\IDinst/RegFile[31][16] ), .DIN2(n1207), 
        .Q(\IDinst/n10475 ) );
  nnd2s1 \IDinst/U10537  ( .DIN1(\IDinst/RegFile[30][16] ), .DIN2(n1253), 
        .Q(\IDinst/n10474 ) );
  nnd2s1 \IDinst/U10536  ( .DIN1(\IDinst/n10472 ), .DIN2(\IDinst/n10471 ), 
        .Q(\IDinst/n10473 ) );
  nnd2s1 \IDinst/U10535  ( .DIN1(\IDinst/RegFile[29][16] ), .DIN2(n1207), 
        .Q(\IDinst/n10472 ) );
  nnd2s1 \IDinst/U10534  ( .DIN1(\IDinst/RegFile[28][16] ), .DIN2(n1253), 
        .Q(\IDinst/n10471 ) );
  nnd2s1 \IDinst/U10533  ( .DIN1(\IDinst/n10469 ), .DIN2(\IDinst/n10468 ), 
        .Q(\IDinst/n10470 ) );
  nnd2s1 \IDinst/U10532  ( .DIN1(\IDinst/n10467 ), .DIN2(n1313), 
        .Q(\IDinst/n10469 ) );
  nnd2s1 \IDinst/U10531  ( .DIN1(\IDinst/n10464 ), .DIN2(n1334), 
        .Q(\IDinst/n10468 ) );
  nnd2s1 \IDinst/U10530  ( .DIN1(\IDinst/n10466 ), .DIN2(\IDinst/n10465 ), 
        .Q(\IDinst/n10467 ) );
  nnd2s1 \IDinst/U10529  ( .DIN1(\IDinst/RegFile[27][16] ), .DIN2(n1207), 
        .Q(\IDinst/n10466 ) );
  nnd2s1 \IDinst/U10528  ( .DIN1(\IDinst/RegFile[26][16] ), .DIN2(n1253), 
        .Q(\IDinst/n10465 ) );
  nnd2s1 \IDinst/U10527  ( .DIN1(\IDinst/n10463 ), .DIN2(\IDinst/n10462 ), 
        .Q(\IDinst/n10464 ) );
  nnd2s1 \IDinst/U10526  ( .DIN1(\IDinst/RegFile[25][16] ), .DIN2(n1207), 
        .Q(\IDinst/n10463 ) );
  nnd2s1 \IDinst/U10525  ( .DIN1(\IDinst/RegFile[24][16] ), .DIN2(n1253), 
        .Q(\IDinst/n10462 ) );
  nnd2s1 \IDinst/U10524  ( .DIN1(\IDinst/n10460 ), .DIN2(\IDinst/n10459 ), 
        .Q(\IDinst/n10461 ) );
  nnd2s1 \IDinst/U10523  ( .DIN1(\IDinst/n10458 ), .DIN2(n1374), 
        .Q(\IDinst/n10460 ) );
  nnd2s1 \IDinst/U10522  ( .DIN1(\IDinst/n10449 ), .DIN2(n1368), 
        .Q(\IDinst/n10459 ) );
  nnd2s1 \IDinst/U10521  ( .DIN1(\IDinst/n10457 ), .DIN2(\IDinst/n10456 ), 
        .Q(\IDinst/n10458 ) );
  nnd2s1 \IDinst/U10520  ( .DIN1(\IDinst/n10455 ), .DIN2(n1313), 
        .Q(\IDinst/n10457 ) );
  nnd2s1 \IDinst/U10519  ( .DIN1(\IDinst/n10452 ), .DIN2(n1333), 
        .Q(\IDinst/n10456 ) );
  nnd2s1 \IDinst/U10518  ( .DIN1(\IDinst/n10454 ), .DIN2(\IDinst/n10453 ), 
        .Q(\IDinst/n10455 ) );
  nnd2s1 \IDinst/U10517  ( .DIN1(\IDinst/RegFile[23][16] ), .DIN2(n1207), 
        .Q(\IDinst/n10454 ) );
  nnd2s1 \IDinst/U10516  ( .DIN1(\IDinst/RegFile[22][16] ), .DIN2(n1253), 
        .Q(\IDinst/n10453 ) );
  nnd2s1 \IDinst/U10515  ( .DIN1(\IDinst/n10451 ), .DIN2(\IDinst/n10450 ), 
        .Q(\IDinst/n10452 ) );
  nnd2s1 \IDinst/U10514  ( .DIN1(\IDinst/RegFile[21][16] ), .DIN2(n1207), 
        .Q(\IDinst/n10451 ) );
  nnd2s1 \IDinst/U10513  ( .DIN1(\IDinst/RegFile[20][16] ), .DIN2(n1253), 
        .Q(\IDinst/n10450 ) );
  nnd2s1 \IDinst/U10512  ( .DIN1(\IDinst/n10448 ), .DIN2(\IDinst/n10447 ), 
        .Q(\IDinst/n10449 ) );
  nnd2s1 \IDinst/U10511  ( .DIN1(\IDinst/n10446 ), .DIN2(n1312), 
        .Q(\IDinst/n10448 ) );
  nnd2s1 \IDinst/U10510  ( .DIN1(\IDinst/n10443 ), .DIN2(n1333), 
        .Q(\IDinst/n10447 ) );
  nnd2s1 \IDinst/U10509  ( .DIN1(\IDinst/n10445 ), .DIN2(\IDinst/n10444 ), 
        .Q(\IDinst/n10446 ) );
  nnd2s1 \IDinst/U10508  ( .DIN1(\IDinst/RegFile[19][16] ), .DIN2(n1207), 
        .Q(\IDinst/n10445 ) );
  nnd2s1 \IDinst/U10507  ( .DIN1(\IDinst/RegFile[18][16] ), .DIN2(n1253), 
        .Q(\IDinst/n10444 ) );
  nnd2s1 \IDinst/U10506  ( .DIN1(\IDinst/n10442 ), .DIN2(\IDinst/n10441 ), 
        .Q(\IDinst/n10443 ) );
  nnd2s1 \IDinst/U10505  ( .DIN1(\IDinst/RegFile[17][16] ), .DIN2(n1207), 
        .Q(\IDinst/n10442 ) );
  nnd2s1 \IDinst/U10504  ( .DIN1(\IDinst/RegFile[16][16] ), .DIN2(n1253), 
        .Q(\IDinst/n10441 ) );
  nnd2s1 \IDinst/U10503  ( .DIN1(\IDinst/n10439 ), .DIN2(\IDinst/n10438 ), 
        .Q(\IDinst/n10440 ) );
  nnd2s1 \IDinst/U10502  ( .DIN1(\IDinst/n10437 ), .DIN2(n666), 
        .Q(\IDinst/n10439 ) );
  nnd2s1 \IDinst/U10501  ( .DIN1(\IDinst/n10416 ), .DIN2(n681), 
        .Q(\IDinst/n10438 ) );
  nnd2s1 \IDinst/U10500  ( .DIN1(\IDinst/n10436 ), .DIN2(\IDinst/n10435 ), 
        .Q(\IDinst/n10437 ) );
  nnd2s1 \IDinst/U10499  ( .DIN1(\IDinst/n10434 ), .DIN2(n1374), 
        .Q(\IDinst/n10436 ) );
  nnd2s1 \IDinst/U10498  ( .DIN1(\IDinst/n10425 ), .DIN2(n1368), 
        .Q(\IDinst/n10435 ) );
  nnd2s1 \IDinst/U10497  ( .DIN1(\IDinst/n10433 ), .DIN2(\IDinst/n10432 ), 
        .Q(\IDinst/n10434 ) );
  nnd2s1 \IDinst/U10496  ( .DIN1(\IDinst/n10431 ), .DIN2(n1312), 
        .Q(\IDinst/n10433 ) );
  nnd2s1 \IDinst/U10495  ( .DIN1(\IDinst/n10428 ), .DIN2(n1333), 
        .Q(\IDinst/n10432 ) );
  nnd2s1 \IDinst/U10494  ( .DIN1(\IDinst/n10430 ), .DIN2(\IDinst/n10429 ), 
        .Q(\IDinst/n10431 ) );
  nnd2s1 \IDinst/U10493  ( .DIN1(\IDinst/RegFile[15][16] ), .DIN2(n1207), 
        .Q(\IDinst/n10430 ) );
  nnd2s1 \IDinst/U10492  ( .DIN1(\IDinst/RegFile[14][16] ), .DIN2(n1252), 
        .Q(\IDinst/n10429 ) );
  nnd2s1 \IDinst/U10491  ( .DIN1(\IDinst/n10427 ), .DIN2(\IDinst/n10426 ), 
        .Q(\IDinst/n10428 ) );
  nnd2s1 \IDinst/U10490  ( .DIN1(\IDinst/RegFile[13][16] ), .DIN2(n1208), 
        .Q(\IDinst/n10427 ) );
  nnd2s1 \IDinst/U10489  ( .DIN1(\IDinst/RegFile[12][16] ), .DIN2(n1252), 
        .Q(\IDinst/n10426 ) );
  nnd2s1 \IDinst/U10488  ( .DIN1(\IDinst/n10424 ), .DIN2(\IDinst/n10423 ), 
        .Q(\IDinst/n10425 ) );
  nnd2s1 \IDinst/U10487  ( .DIN1(\IDinst/n10422 ), .DIN2(n1312), 
        .Q(\IDinst/n10424 ) );
  nnd2s1 \IDinst/U10486  ( .DIN1(\IDinst/n10419 ), .DIN2(n1333), 
        .Q(\IDinst/n10423 ) );
  nnd2s1 \IDinst/U10485  ( .DIN1(\IDinst/n10421 ), .DIN2(\IDinst/n10420 ), 
        .Q(\IDinst/n10422 ) );
  nnd2s1 \IDinst/U10484  ( .DIN1(\IDinst/RegFile[11][16] ), .DIN2(n1208), 
        .Q(\IDinst/n10421 ) );
  nnd2s1 \IDinst/U10483  ( .DIN1(\IDinst/RegFile[10][16] ), .DIN2(n1252), 
        .Q(\IDinst/n10420 ) );
  nnd2s1 \IDinst/U10482  ( .DIN1(\IDinst/n10418 ), .DIN2(\IDinst/n10417 ), 
        .Q(\IDinst/n10419 ) );
  nnd2s1 \IDinst/U10481  ( .DIN1(\IDinst/RegFile[9][16] ), .DIN2(n1208), 
        .Q(\IDinst/n10418 ) );
  nnd2s1 \IDinst/U10480  ( .DIN1(\IDinst/RegFile[8][16] ), .DIN2(n1252), 
        .Q(\IDinst/n10417 ) );
  nnd2s1 \IDinst/U10479  ( .DIN1(\IDinst/n10415 ), .DIN2(\IDinst/n10414 ), 
        .Q(\IDinst/n10416 ) );
  nnd2s1 \IDinst/U10478  ( .DIN1(\IDinst/n10413 ), .DIN2(n1374), 
        .Q(\IDinst/n10415 ) );
  nnd2s1 \IDinst/U10477  ( .DIN1(\IDinst/n10404 ), .DIN2(n1368), 
        .Q(\IDinst/n10414 ) );
  nnd2s1 \IDinst/U10476  ( .DIN1(\IDinst/n10412 ), .DIN2(\IDinst/n10411 ), 
        .Q(\IDinst/n10413 ) );
  nnd2s1 \IDinst/U10475  ( .DIN1(\IDinst/n10410 ), .DIN2(n1317), 
        .Q(\IDinst/n10412 ) );
  nnd2s1 \IDinst/U10474  ( .DIN1(\IDinst/n10407 ), .DIN2(n1333), 
        .Q(\IDinst/n10411 ) );
  nnd2s1 \IDinst/U10473  ( .DIN1(\IDinst/n10409 ), .DIN2(\IDinst/n10408 ), 
        .Q(\IDinst/n10410 ) );
  nnd2s1 \IDinst/U10472  ( .DIN1(\IDinst/RegFile[7][16] ), .DIN2(n1208), 
        .Q(\IDinst/n10409 ) );
  nnd2s1 \IDinst/U10471  ( .DIN1(\IDinst/RegFile[6][16] ), .DIN2(n1252), 
        .Q(\IDinst/n10408 ) );
  nnd2s1 \IDinst/U10470  ( .DIN1(\IDinst/n10406 ), .DIN2(\IDinst/n10405 ), 
        .Q(\IDinst/n10407 ) );
  nnd2s1 \IDinst/U10469  ( .DIN1(\IDinst/RegFile[5][16] ), .DIN2(n1208), 
        .Q(\IDinst/n10406 ) );
  nnd2s1 \IDinst/U10468  ( .DIN1(\IDinst/RegFile[4][16] ), .DIN2(n1252), 
        .Q(\IDinst/n10405 ) );
  nnd2s1 \IDinst/U10467  ( .DIN1(\IDinst/n10403 ), .DIN2(\IDinst/n10402 ), 
        .Q(\IDinst/n10404 ) );
  nnd2s1 \IDinst/U10466  ( .DIN1(\IDinst/n10401 ), .DIN2(n1363), 
        .Q(\IDinst/n10403 ) );
  nnd2s1 \IDinst/U10465  ( .DIN1(\IDinst/n10398 ), .DIN2(n1334), 
        .Q(\IDinst/n10402 ) );
  nnd2s1 \IDinst/U10464  ( .DIN1(\IDinst/n10400 ), .DIN2(\IDinst/n10399 ), 
        .Q(\IDinst/n10401 ) );
  nnd2s1 \IDinst/U10463  ( .DIN1(\IDinst/RegFile[3][16] ), .DIN2(n1208), 
        .Q(\IDinst/n10400 ) );
  nnd2s1 \IDinst/U10462  ( .DIN1(\IDinst/RegFile[2][16] ), .DIN2(n1252), 
        .Q(\IDinst/n10399 ) );
  nnd2s1 \IDinst/U10461  ( .DIN1(\IDinst/n10397 ), .DIN2(\IDinst/n10396 ), 
        .Q(\IDinst/n10398 ) );
  nnd2s1 \IDinst/U10460  ( .DIN1(\IDinst/RegFile[1][16] ), .DIN2(n1208), 
        .Q(\IDinst/n10397 ) );
  nnd2s1 \IDinst/U10459  ( .DIN1(\IDinst/RegFile[0][16] ), .DIN2(n1252), 
        .Q(\IDinst/n10396 ) );
  nnd2s1 \IDinst/U10458  ( .DIN1(\IDinst/n10395 ), .DIN2(n535), 
        .Q(\IDinst/n8922 ) );
  nnd2s1 \IDinst/U10457  ( .DIN1(\IDinst/n10350 ), .DIN2(n533), 
        .Q(\IDinst/n8923 ) );
  nnd2s1 \IDinst/U10456  ( .DIN1(\IDinst/n10394 ), .DIN2(\IDinst/n10393 ), 
        .Q(\IDinst/n10395 ) );
  nnd2s1 \IDinst/U10455  ( .DIN1(\IDinst/n10392 ), .DIN2(n667), 
        .Q(\IDinst/n10394 ) );
  nnd2s1 \IDinst/U10454  ( .DIN1(\IDinst/n10371 ), .DIN2(n683), 
        .Q(\IDinst/n10393 ) );
  nnd2s1 \IDinst/U10453  ( .DIN1(\IDinst/n10391 ), .DIN2(\IDinst/n10390 ), 
        .Q(\IDinst/n10392 ) );
  nnd2s1 \IDinst/U10452  ( .DIN1(\IDinst/n10389 ), .DIN2(n1375), 
        .Q(\IDinst/n10391 ) );
  nnd2s1 \IDinst/U10451  ( .DIN1(\IDinst/n10380 ), .DIN2(n1368), 
        .Q(\IDinst/n10390 ) );
  nnd2s1 \IDinst/U10450  ( .DIN1(\IDinst/n10388 ), .DIN2(\IDinst/n10387 ), 
        .Q(\IDinst/n10389 ) );
  nnd2s1 \IDinst/U10449  ( .DIN1(\IDinst/n10386 ), .DIN2(n1362), 
        .Q(\IDinst/n10388 ) );
  nnd2s1 \IDinst/U10448  ( .DIN1(\IDinst/n10383 ), .DIN2(n1334), 
        .Q(\IDinst/n10387 ) );
  nnd2s1 \IDinst/U10447  ( .DIN1(\IDinst/n10385 ), .DIN2(\IDinst/n10384 ), 
        .Q(\IDinst/n10386 ) );
  nnd2s1 \IDinst/U10446  ( .DIN1(\IDinst/RegFile[31][15] ), .DIN2(n1233), 
        .Q(\IDinst/n10385 ) );
  nnd2s1 \IDinst/U10445  ( .DIN1(\IDinst/RegFile[30][15] ), .DIN2(n1252), 
        .Q(\IDinst/n10384 ) );
  nnd2s1 \IDinst/U10444  ( .DIN1(\IDinst/n10382 ), .DIN2(\IDinst/n10381 ), 
        .Q(\IDinst/n10383 ) );
  nnd2s1 \IDinst/U10443  ( .DIN1(\IDinst/RegFile[29][15] ), .DIN2(n1228), 
        .Q(\IDinst/n10382 ) );
  nnd2s1 \IDinst/U10442  ( .DIN1(\IDinst/RegFile[28][15] ), .DIN2(n1251), 
        .Q(\IDinst/n10381 ) );
  nnd2s1 \IDinst/U10441  ( .DIN1(\IDinst/n10379 ), .DIN2(\IDinst/n10378 ), 
        .Q(\IDinst/n10380 ) );
  nnd2s1 \IDinst/U10440  ( .DIN1(\IDinst/n10377 ), .DIN2(\IDinst/N45 ), 
        .Q(\IDinst/n10379 ) );
  nnd2s1 \IDinst/U10439  ( .DIN1(\IDinst/n10374 ), .DIN2(n1334), 
        .Q(\IDinst/n10378 ) );
  nnd2s1 \IDinst/U10438  ( .DIN1(\IDinst/n10376 ), .DIN2(\IDinst/n10375 ), 
        .Q(\IDinst/n10377 ) );
  nnd2s1 \IDinst/U10437  ( .DIN1(\IDinst/RegFile[27][15] ), .DIN2(n1228), 
        .Q(\IDinst/n10376 ) );
  nnd2s1 \IDinst/U10436  ( .DIN1(\IDinst/RegFile[26][15] ), .DIN2(n1251), 
        .Q(\IDinst/n10375 ) );
  nnd2s1 \IDinst/U10435  ( .DIN1(\IDinst/n10373 ), .DIN2(\IDinst/n10372 ), 
        .Q(\IDinst/n10374 ) );
  nnd2s1 \IDinst/U10434  ( .DIN1(\IDinst/RegFile[25][15] ), .DIN2(n1228), 
        .Q(\IDinst/n10373 ) );
  nnd2s1 \IDinst/U10433  ( .DIN1(\IDinst/RegFile[24][15] ), .DIN2(n1251), 
        .Q(\IDinst/n10372 ) );
  nnd2s1 \IDinst/U10432  ( .DIN1(\IDinst/n10370 ), .DIN2(\IDinst/n10369 ), 
        .Q(\IDinst/n10371 ) );
  nnd2s1 \IDinst/U10431  ( .DIN1(\IDinst/n10368 ), .DIN2(n1375), 
        .Q(\IDinst/n10370 ) );
  nnd2s1 \IDinst/U10430  ( .DIN1(\IDinst/n10359 ), .DIN2(n1368), 
        .Q(\IDinst/n10369 ) );
  nnd2s1 \IDinst/U10429  ( .DIN1(\IDinst/n10367 ), .DIN2(\IDinst/n10366 ), 
        .Q(\IDinst/n10368 ) );
  nnd2s1 \IDinst/U10428  ( .DIN1(\IDinst/n10365 ), .DIN2(\IDinst/N45 ), 
        .Q(\IDinst/n10367 ) );
  nnd2s1 \IDinst/U10427  ( .DIN1(\IDinst/n10362 ), .DIN2(n1334), 
        .Q(\IDinst/n10366 ) );
  nnd2s1 \IDinst/U10426  ( .DIN1(\IDinst/n10364 ), .DIN2(\IDinst/n10363 ), 
        .Q(\IDinst/n10365 ) );
  nnd2s1 \IDinst/U10425  ( .DIN1(\IDinst/RegFile[23][15] ), .DIN2(n1228), 
        .Q(\IDinst/n10364 ) );
  nnd2s1 \IDinst/U10424  ( .DIN1(\IDinst/RegFile[22][15] ), .DIN2(n1251), 
        .Q(\IDinst/n10363 ) );
  nnd2s1 \IDinst/U10423  ( .DIN1(\IDinst/n10361 ), .DIN2(\IDinst/n10360 ), 
        .Q(\IDinst/n10362 ) );
  nnd2s1 \IDinst/U10422  ( .DIN1(\IDinst/RegFile[21][15] ), .DIN2(n1228), 
        .Q(\IDinst/n10361 ) );
  nnd2s1 \IDinst/U10421  ( .DIN1(\IDinst/RegFile[20][15] ), .DIN2(n1251), 
        .Q(\IDinst/n10360 ) );
  nnd2s1 \IDinst/U10420  ( .DIN1(\IDinst/n10358 ), .DIN2(\IDinst/n10357 ), 
        .Q(\IDinst/n10359 ) );
  nnd2s1 \IDinst/U10419  ( .DIN1(\IDinst/n10356 ), .DIN2(n1331), 
        .Q(\IDinst/n10358 ) );
  nnd2s1 \IDinst/U10418  ( .DIN1(\IDinst/n10353 ), .DIN2(n1334), 
        .Q(\IDinst/n10357 ) );
  nnd2s1 \IDinst/U10417  ( .DIN1(\IDinst/n10355 ), .DIN2(\IDinst/n10354 ), 
        .Q(\IDinst/n10356 ) );
  nnd2s1 \IDinst/U10416  ( .DIN1(\IDinst/RegFile[19][15] ), .DIN2(n1228), 
        .Q(\IDinst/n10355 ) );
  nnd2s1 \IDinst/U10415  ( .DIN1(\IDinst/RegFile[18][15] ), .DIN2(n1251), 
        .Q(\IDinst/n10354 ) );
  nnd2s1 \IDinst/U10414  ( .DIN1(\IDinst/n10352 ), .DIN2(\IDinst/n10351 ), 
        .Q(\IDinst/n10353 ) );
  nnd2s1 \IDinst/U10413  ( .DIN1(\IDinst/RegFile[17][15] ), .DIN2(n1228), 
        .Q(\IDinst/n10352 ) );
  nnd2s1 \IDinst/U10412  ( .DIN1(\IDinst/RegFile[16][15] ), .DIN2(n1251), 
        .Q(\IDinst/n10351 ) );
  nnd2s1 \IDinst/U10411  ( .DIN1(\IDinst/n10349 ), .DIN2(\IDinst/n10348 ), 
        .Q(\IDinst/n10350 ) );
  nnd2s1 \IDinst/U10410  ( .DIN1(\IDinst/n10347 ), .DIN2(n665), 
        .Q(\IDinst/n10349 ) );
  nnd2s1 \IDinst/U10409  ( .DIN1(\IDinst/n10326 ), .DIN2(n682), 
        .Q(\IDinst/n10348 ) );
  nnd2s1 \IDinst/U10408  ( .DIN1(\IDinst/n10346 ), .DIN2(\IDinst/n10345 ), 
        .Q(\IDinst/n10347 ) );
  nnd2s1 \IDinst/U10407  ( .DIN1(\IDinst/n10344 ), .DIN2(n1375), 
        .Q(\IDinst/n10346 ) );
  nnd2s1 \IDinst/U10406  ( .DIN1(\IDinst/n10335 ), .DIN2(n1368), 
        .Q(\IDinst/n10345 ) );
  nnd2s1 \IDinst/U10405  ( .DIN1(\IDinst/n10343 ), .DIN2(\IDinst/n10342 ), 
        .Q(\IDinst/n10344 ) );
  nnd2s1 \IDinst/U10404  ( .DIN1(\IDinst/n10341 ), .DIN2(n1331), 
        .Q(\IDinst/n10343 ) );
  nnd2s1 \IDinst/U10403  ( .DIN1(\IDinst/n10338 ), .DIN2(n1334), 
        .Q(\IDinst/n10342 ) );
  nnd2s1 \IDinst/U10402  ( .DIN1(\IDinst/n10340 ), .DIN2(\IDinst/n10339 ), 
        .Q(\IDinst/n10341 ) );
  nnd2s1 \IDinst/U10401  ( .DIN1(\IDinst/RegFile[15][15] ), .DIN2(n1228), 
        .Q(\IDinst/n10340 ) );
  nnd2s1 \IDinst/U10400  ( .DIN1(\IDinst/RegFile[14][15] ), .DIN2(n1251), 
        .Q(\IDinst/n10339 ) );
  nnd2s1 \IDinst/U10399  ( .DIN1(\IDinst/n10337 ), .DIN2(\IDinst/n10336 ), 
        .Q(\IDinst/n10338 ) );
  nnd2s1 \IDinst/U10398  ( .DIN1(\IDinst/RegFile[13][15] ), .DIN2(n1228), 
        .Q(\IDinst/n10337 ) );
  nnd2s1 \IDinst/U10397  ( .DIN1(\IDinst/RegFile[12][15] ), .DIN2(n1251), 
        .Q(\IDinst/n10336 ) );
  nnd2s1 \IDinst/U10396  ( .DIN1(\IDinst/n10334 ), .DIN2(\IDinst/n10333 ), 
        .Q(\IDinst/n10335 ) );
  nnd2s1 \IDinst/U10395  ( .DIN1(\IDinst/n10332 ), .DIN2(n1331), 
        .Q(\IDinst/n10334 ) );
  nnd2s1 \IDinst/U10394  ( .DIN1(\IDinst/n10329 ), .DIN2(n1335), 
        .Q(\IDinst/n10333 ) );
  nnd2s1 \IDinst/U10393  ( .DIN1(\IDinst/n10331 ), .DIN2(\IDinst/n10330 ), 
        .Q(\IDinst/n10332 ) );
  nnd2s1 \IDinst/U10392  ( .DIN1(\IDinst/RegFile[11][15] ), .DIN2(n1228), 
        .Q(\IDinst/n10331 ) );
  nnd2s1 \IDinst/U10391  ( .DIN1(\IDinst/RegFile[10][15] ), .DIN2(n1250), 
        .Q(\IDinst/n10330 ) );
  nnd2s1 \IDinst/U10390  ( .DIN1(\IDinst/n10328 ), .DIN2(\IDinst/n10327 ), 
        .Q(\IDinst/n10329 ) );
  nnd2s1 \IDinst/U10389  ( .DIN1(\IDinst/RegFile[9][15] ), .DIN2(n1229), 
        .Q(\IDinst/n10328 ) );
  nnd2s1 \IDinst/U10388  ( .DIN1(\IDinst/RegFile[8][15] ), .DIN2(n1250), 
        .Q(\IDinst/n10327 ) );
  nnd2s1 \IDinst/U10387  ( .DIN1(\IDinst/n10325 ), .DIN2(\IDinst/n10324 ), 
        .Q(\IDinst/n10326 ) );
  nnd2s1 \IDinst/U10386  ( .DIN1(\IDinst/n10323 ), .DIN2(n1375), 
        .Q(\IDinst/n10325 ) );
  nnd2s1 \IDinst/U10385  ( .DIN1(\IDinst/n10314 ), .DIN2(n1368), 
        .Q(\IDinst/n10324 ) );
  nnd2s1 \IDinst/U10384  ( .DIN1(\IDinst/n10322 ), .DIN2(\IDinst/n10321 ), 
        .Q(\IDinst/n10323 ) );
  nnd2s1 \IDinst/U10383  ( .DIN1(\IDinst/n10320 ), .DIN2(n1331), 
        .Q(\IDinst/n10322 ) );
  nnd2s1 \IDinst/U10382  ( .DIN1(\IDinst/n10317 ), .DIN2(n1334), 
        .Q(\IDinst/n10321 ) );
  nnd2s1 \IDinst/U10381  ( .DIN1(\IDinst/n10319 ), .DIN2(\IDinst/n10318 ), 
        .Q(\IDinst/n10320 ) );
  nnd2s1 \IDinst/U10380  ( .DIN1(\IDinst/RegFile[7][15] ), .DIN2(n1229), 
        .Q(\IDinst/n10319 ) );
  nnd2s1 \IDinst/U10379  ( .DIN1(\IDinst/RegFile[6][15] ), .DIN2(n1250), 
        .Q(\IDinst/n10318 ) );
  nnd2s1 \IDinst/U10378  ( .DIN1(\IDinst/n10316 ), .DIN2(\IDinst/n10315 ), 
        .Q(\IDinst/n10317 ) );
  nnd2s1 \IDinst/U10377  ( .DIN1(\IDinst/RegFile[5][15] ), .DIN2(n1229), 
        .Q(\IDinst/n10316 ) );
  nnd2s1 \IDinst/U10376  ( .DIN1(\IDinst/RegFile[4][15] ), .DIN2(n1250), 
        .Q(\IDinst/n10315 ) );
  nnd2s1 \IDinst/U10375  ( .DIN1(\IDinst/n10313 ), .DIN2(\IDinst/n10312 ), 
        .Q(\IDinst/n10314 ) );
  nnd2s1 \IDinst/U10374  ( .DIN1(\IDinst/n10311 ), .DIN2(n1331), 
        .Q(\IDinst/n10313 ) );
  nnd2s1 \IDinst/U10373  ( .DIN1(\IDinst/n10308 ), .DIN2(n1334), 
        .Q(\IDinst/n10312 ) );
  nnd2s1 \IDinst/U10372  ( .DIN1(\IDinst/n10310 ), .DIN2(\IDinst/n10309 ), 
        .Q(\IDinst/n10311 ) );
  nnd2s1 \IDinst/U10371  ( .DIN1(\IDinst/RegFile[3][15] ), .DIN2(n1229), 
        .Q(\IDinst/n10310 ) );
  nnd2s1 \IDinst/U10370  ( .DIN1(\IDinst/RegFile[2][15] ), .DIN2(n1250), 
        .Q(\IDinst/n10309 ) );
  nnd2s1 \IDinst/U10369  ( .DIN1(\IDinst/n10307 ), .DIN2(\IDinst/n10306 ), 
        .Q(\IDinst/n10308 ) );
  nnd2s1 \IDinst/U10368  ( .DIN1(\IDinst/RegFile[1][15] ), .DIN2(n1229), 
        .Q(\IDinst/n10307 ) );
  nnd2s1 \IDinst/U10367  ( .DIN1(\IDinst/RegFile[0][15] ), .DIN2(n1250), 
        .Q(\IDinst/n10306 ) );
  nnd2s1 \IDinst/U10366  ( .DIN1(\IDinst/n10305 ), .DIN2(n534), 
        .Q(\IDinst/n8920 ) );
  nnd2s1 \IDinst/U10365  ( .DIN1(\IDinst/n10260 ), .DIN2(n634), 
        .Q(\IDinst/n8921 ) );
  nnd2s1 \IDinst/U10364  ( .DIN1(\IDinst/n10304 ), .DIN2(\IDinst/n10303 ), 
        .Q(\IDinst/n10305 ) );
  nnd2s1 \IDinst/U10363  ( .DIN1(\IDinst/n10302 ), .DIN2(n668), 
        .Q(\IDinst/n10304 ) );
  nnd2s1 \IDinst/U10362  ( .DIN1(\IDinst/n10281 ), .DIN2(n680), 
        .Q(\IDinst/n10303 ) );
  nnd2s1 \IDinst/U10361  ( .DIN1(\IDinst/n10301 ), .DIN2(\IDinst/n10300 ), 
        .Q(\IDinst/n10302 ) );
  nnd2s1 \IDinst/U10360  ( .DIN1(\IDinst/n10299 ), .DIN2(n1375), 
        .Q(\IDinst/n10301 ) );
  nnd2s1 \IDinst/U10359  ( .DIN1(\IDinst/n10290 ), .DIN2(n1368), 
        .Q(\IDinst/n10300 ) );
  nnd2s1 \IDinst/U10358  ( .DIN1(\IDinst/n10298 ), .DIN2(\IDinst/n10297 ), 
        .Q(\IDinst/n10299 ) );
  nnd2s1 \IDinst/U10357  ( .DIN1(\IDinst/n10296 ), .DIN2(n1331), 
        .Q(\IDinst/n10298 ) );
  nnd2s1 \IDinst/U10356  ( .DIN1(\IDinst/n10293 ), .DIN2(n1335), 
        .Q(\IDinst/n10297 ) );
  nnd2s1 \IDinst/U10355  ( .DIN1(\IDinst/n10295 ), .DIN2(\IDinst/n10294 ), 
        .Q(\IDinst/n10296 ) );
  nnd2s1 \IDinst/U10354  ( .DIN1(\IDinst/RegFile[31][14] ), .DIN2(n1229), 
        .Q(\IDinst/n10295 ) );
  nnd2s1 \IDinst/U10353  ( .DIN1(\IDinst/RegFile[30][14] ), .DIN2(n1250), 
        .Q(\IDinst/n10294 ) );
  nnd2s1 \IDinst/U10352  ( .DIN1(\IDinst/n10292 ), .DIN2(\IDinst/n10291 ), 
        .Q(\IDinst/n10293 ) );
  nnd2s1 \IDinst/U10351  ( .DIN1(\IDinst/RegFile[29][14] ), .DIN2(n1229), 
        .Q(\IDinst/n10292 ) );
  nnd2s1 \IDinst/U10350  ( .DIN1(\IDinst/RegFile[28][14] ), .DIN2(n1250), 
        .Q(\IDinst/n10291 ) );
  nnd2s1 \IDinst/U10349  ( .DIN1(\IDinst/n10289 ), .DIN2(\IDinst/n10288 ), 
        .Q(\IDinst/n10290 ) );
  nnd2s1 \IDinst/U10348  ( .DIN1(\IDinst/n10287 ), .DIN2(n1331), 
        .Q(\IDinst/n10289 ) );
  nnd2s1 \IDinst/U10347  ( .DIN1(\IDinst/n10284 ), .DIN2(n1335), 
        .Q(\IDinst/n10288 ) );
  nnd2s1 \IDinst/U10346  ( .DIN1(\IDinst/n10286 ), .DIN2(\IDinst/n10285 ), 
        .Q(\IDinst/n10287 ) );
  nnd2s1 \IDinst/U10345  ( .DIN1(\IDinst/RegFile[27][14] ), .DIN2(n1229), 
        .Q(\IDinst/n10286 ) );
  nnd2s1 \IDinst/U10344  ( .DIN1(\IDinst/RegFile[26][14] ), .DIN2(n1250), 
        .Q(\IDinst/n10285 ) );
  nnd2s1 \IDinst/U10343  ( .DIN1(\IDinst/n10283 ), .DIN2(\IDinst/n10282 ), 
        .Q(\IDinst/n10284 ) );
  nnd2s1 \IDinst/U10342  ( .DIN1(\IDinst/RegFile[25][14] ), .DIN2(n1229), 
        .Q(\IDinst/n10283 ) );
  nnd2s1 \IDinst/U10341  ( .DIN1(\IDinst/RegFile[24][14] ), .DIN2(n1249), 
        .Q(\IDinst/n10282 ) );
  nnd2s1 \IDinst/U10340  ( .DIN1(\IDinst/n10280 ), .DIN2(\IDinst/n10279 ), 
        .Q(\IDinst/n10281 ) );
  nnd2s1 \IDinst/U10339  ( .DIN1(\IDinst/n10278 ), .DIN2(n1375), 
        .Q(\IDinst/n10280 ) );
  nnd2s1 \IDinst/U10338  ( .DIN1(\IDinst/n10269 ), .DIN2(n1368), 
        .Q(\IDinst/n10279 ) );
  nnd2s1 \IDinst/U10337  ( .DIN1(\IDinst/n10277 ), .DIN2(\IDinst/n10276 ), 
        .Q(\IDinst/n10278 ) );
  nnd2s1 \IDinst/U10336  ( .DIN1(\IDinst/n10275 ), .DIN2(n1331), 
        .Q(\IDinst/n10277 ) );
  nnd2s1 \IDinst/U10335  ( .DIN1(\IDinst/n10272 ), .DIN2(n1335), 
        .Q(\IDinst/n10276 ) );
  nnd2s1 \IDinst/U10334  ( .DIN1(\IDinst/n10274 ), .DIN2(\IDinst/n10273 ), 
        .Q(\IDinst/n10275 ) );
  nnd2s1 \IDinst/U10333  ( .DIN1(\IDinst/RegFile[23][14] ), .DIN2(n1229), 
        .Q(\IDinst/n10274 ) );
  nnd2s1 \IDinst/U10332  ( .DIN1(\IDinst/RegFile[22][14] ), .DIN2(n1249), 
        .Q(\IDinst/n10273 ) );
  nnd2s1 \IDinst/U10331  ( .DIN1(\IDinst/n10271 ), .DIN2(\IDinst/n10270 ), 
        .Q(\IDinst/n10272 ) );
  nnd2s1 \IDinst/U10330  ( .DIN1(\IDinst/RegFile[21][14] ), .DIN2(n1229), 
        .Q(\IDinst/n10271 ) );
  nnd2s1 \IDinst/U10329  ( .DIN1(\IDinst/RegFile[20][14] ), .DIN2(n1249), 
        .Q(\IDinst/n10270 ) );
  nnd2s1 \IDinst/U10328  ( .DIN1(\IDinst/n10268 ), .DIN2(\IDinst/n10267 ), 
        .Q(\IDinst/n10269 ) );
  nnd2s1 \IDinst/U10327  ( .DIN1(\IDinst/n10266 ), .DIN2(n1331), 
        .Q(\IDinst/n10268 ) );
  nnd2s1 \IDinst/U10326  ( .DIN1(\IDinst/n10263 ), .DIN2(n1335), 
        .Q(\IDinst/n10267 ) );
  nnd2s1 \IDinst/U10325  ( .DIN1(\IDinst/n10265 ), .DIN2(\IDinst/n10264 ), 
        .Q(\IDinst/n10266 ) );
  nnd2s1 \IDinst/U10324  ( .DIN1(\IDinst/RegFile[19][14] ), .DIN2(n1229), 
        .Q(\IDinst/n10265 ) );
  nnd2s1 \IDinst/U10323  ( .DIN1(\IDinst/RegFile[18][14] ), .DIN2(n1249), 
        .Q(\IDinst/n10264 ) );
  nnd2s1 \IDinst/U10322  ( .DIN1(\IDinst/n10262 ), .DIN2(\IDinst/n10261 ), 
        .Q(\IDinst/n10263 ) );
  nnd2s1 \IDinst/U10321  ( .DIN1(\IDinst/RegFile[17][14] ), .DIN2(n1229), 
        .Q(\IDinst/n10262 ) );
  nnd2s1 \IDinst/U10320  ( .DIN1(\IDinst/RegFile[16][14] ), .DIN2(n1249), 
        .Q(\IDinst/n10261 ) );
  nnd2s1 \IDinst/U10319  ( .DIN1(\IDinst/n10259 ), .DIN2(\IDinst/n10258 ), 
        .Q(\IDinst/n10260 ) );
  nnd2s1 \IDinst/U10318  ( .DIN1(\IDinst/n10257 ), .DIN2(n666), 
        .Q(\IDinst/n10259 ) );
  nnd2s1 \IDinst/U10317  ( .DIN1(\IDinst/n10236 ), .DIN2(n681), 
        .Q(\IDinst/n10258 ) );
  nnd2s1 \IDinst/U10316  ( .DIN1(\IDinst/n10256 ), .DIN2(\IDinst/n10255 ), 
        .Q(\IDinst/n10257 ) );
  nnd2s1 \IDinst/U10315  ( .DIN1(\IDinst/n10254 ), .DIN2(n1375), 
        .Q(\IDinst/n10256 ) );
  nnd2s1 \IDinst/U10314  ( .DIN1(\IDinst/n10245 ), .DIN2(n1368), 
        .Q(\IDinst/n10255 ) );
  nnd2s1 \IDinst/U10313  ( .DIN1(\IDinst/n10253 ), .DIN2(\IDinst/n10252 ), 
        .Q(\IDinst/n10254 ) );
  nnd2s1 \IDinst/U10312  ( .DIN1(\IDinst/n10251 ), .DIN2(n1331), 
        .Q(\IDinst/n10253 ) );
  nnd2s1 \IDinst/U10311  ( .DIN1(\IDinst/n10248 ), .DIN2(n1335), 
        .Q(\IDinst/n10252 ) );
  nnd2s1 \IDinst/U10310  ( .DIN1(\IDinst/n10250 ), .DIN2(\IDinst/n10249 ), 
        .Q(\IDinst/n10251 ) );
  nnd2s1 \IDinst/U10309  ( .DIN1(\IDinst/RegFile[15][14] ), .DIN2(n1230), 
        .Q(\IDinst/n10250 ) );
  nnd2s1 \IDinst/U10308  ( .DIN1(\IDinst/RegFile[14][14] ), .DIN2(n1249), 
        .Q(\IDinst/n10249 ) );
  nnd2s1 \IDinst/U10307  ( .DIN1(\IDinst/n10247 ), .DIN2(\IDinst/n10246 ), 
        .Q(\IDinst/n10248 ) );
  nnd2s1 \IDinst/U10306  ( .DIN1(\IDinst/RegFile[13][14] ), .DIN2(n1230), 
        .Q(\IDinst/n10247 ) );
  nnd2s1 \IDinst/U10305  ( .DIN1(\IDinst/RegFile[12][14] ), .DIN2(n1249), 
        .Q(\IDinst/n10246 ) );
  nnd2s1 \IDinst/U10304  ( .DIN1(\IDinst/n10244 ), .DIN2(\IDinst/n10243 ), 
        .Q(\IDinst/n10245 ) );
  nnd2s1 \IDinst/U10303  ( .DIN1(\IDinst/n10242 ), .DIN2(n1331), 
        .Q(\IDinst/n10244 ) );
  nnd2s1 \IDinst/U10302  ( .DIN1(\IDinst/n10239 ), .DIN2(n1335), 
        .Q(\IDinst/n10243 ) );
  nnd2s1 \IDinst/U10301  ( .DIN1(\IDinst/n10241 ), .DIN2(\IDinst/n10240 ), 
        .Q(\IDinst/n10242 ) );
  nnd2s1 \IDinst/U10300  ( .DIN1(\IDinst/RegFile[11][14] ), .DIN2(n1230), 
        .Q(\IDinst/n10241 ) );
  nnd2s1 \IDinst/U10299  ( .DIN1(\IDinst/RegFile[10][14] ), .DIN2(n1249), 
        .Q(\IDinst/n10240 ) );
  nnd2s1 \IDinst/U10298  ( .DIN1(\IDinst/n10238 ), .DIN2(\IDinst/n10237 ), 
        .Q(\IDinst/n10239 ) );
  nnd2s1 \IDinst/U10297  ( .DIN1(\IDinst/RegFile[9][14] ), .DIN2(n1230), 
        .Q(\IDinst/n10238 ) );
  nnd2s1 \IDinst/U10296  ( .DIN1(\IDinst/RegFile[8][14] ), .DIN2(n1249), 
        .Q(\IDinst/n10237 ) );
  nnd2s1 \IDinst/U10295  ( .DIN1(\IDinst/n10235 ), .DIN2(\IDinst/n10234 ), 
        .Q(\IDinst/n10236 ) );
  nnd2s1 \IDinst/U10294  ( .DIN1(\IDinst/n10233 ), .DIN2(n1375), 
        .Q(\IDinst/n10235 ) );
  nnd2s1 \IDinst/U10293  ( .DIN1(\IDinst/n10224 ), .DIN2(n1368), 
        .Q(\IDinst/n10234 ) );
  nnd2s1 \IDinst/U10292  ( .DIN1(\IDinst/n10232 ), .DIN2(\IDinst/n10231 ), 
        .Q(\IDinst/n10233 ) );
  nnd2s1 \IDinst/U10291  ( .DIN1(\IDinst/n10230 ), .DIN2(n1331), 
        .Q(\IDinst/n10232 ) );
  nnd2s1 \IDinst/U10290  ( .DIN1(\IDinst/n10227 ), .DIN2(n1335), 
        .Q(\IDinst/n10231 ) );
  nnd2s1 \IDinst/U10289  ( .DIN1(\IDinst/n10229 ), .DIN2(\IDinst/n10228 ), 
        .Q(\IDinst/n10230 ) );
  nnd2s1 \IDinst/U10288  ( .DIN1(\IDinst/RegFile[7][14] ), .DIN2(n1230), 
        .Q(\IDinst/n10229 ) );
  nnd2s1 \IDinst/U10287  ( .DIN1(\IDinst/RegFile[6][14] ), .DIN2(n1248), 
        .Q(\IDinst/n10228 ) );
  nnd2s1 \IDinst/U10286  ( .DIN1(\IDinst/n10226 ), .DIN2(\IDinst/n10225 ), 
        .Q(\IDinst/n10227 ) );
  nnd2s1 \IDinst/U10285  ( .DIN1(\IDinst/RegFile[5][14] ), .DIN2(n1230), 
        .Q(\IDinst/n10226 ) );
  nnd2s1 \IDinst/U10284  ( .DIN1(\IDinst/RegFile[4][14] ), .DIN2(n1248), 
        .Q(\IDinst/n10225 ) );
  nnd2s1 \IDinst/U10283  ( .DIN1(\IDinst/n10223 ), .DIN2(\IDinst/n10222 ), 
        .Q(\IDinst/n10224 ) );
  nnd2s1 \IDinst/U10282  ( .DIN1(\IDinst/n10221 ), .DIN2(n1331), 
        .Q(\IDinst/n10223 ) );
  nnd2s1 \IDinst/U10281  ( .DIN1(\IDinst/n10218 ), .DIN2(n1335), 
        .Q(\IDinst/n10222 ) );
  nnd2s1 \IDinst/U10280  ( .DIN1(\IDinst/n10220 ), .DIN2(\IDinst/n10219 ), 
        .Q(\IDinst/n10221 ) );
  nnd2s1 \IDinst/U10279  ( .DIN1(\IDinst/RegFile[3][14] ), .DIN2(n1230), 
        .Q(\IDinst/n10220 ) );
  nnd2s1 \IDinst/U10278  ( .DIN1(\IDinst/RegFile[2][14] ), .DIN2(n1248), 
        .Q(\IDinst/n10219 ) );
  nnd2s1 \IDinst/U10277  ( .DIN1(\IDinst/n10217 ), .DIN2(\IDinst/n10216 ), 
        .Q(\IDinst/n10218 ) );
  nnd2s1 \IDinst/U10276  ( .DIN1(\IDinst/RegFile[1][14] ), .DIN2(n1230), 
        .Q(\IDinst/n10217 ) );
  nnd2s1 \IDinst/U10275  ( .DIN1(\IDinst/RegFile[0][14] ), .DIN2(n1248), 
        .Q(\IDinst/n10216 ) );
  nnd2s1 \IDinst/U10274  ( .DIN1(\IDinst/n10215 ), .DIN2(\IDinst/N48 ), 
        .Q(\IDinst/n8918 ) );
  nnd2s1 \IDinst/U10273  ( .DIN1(\IDinst/n10170 ), .DIN2(n533), 
        .Q(\IDinst/n8919 ) );
  nnd2s1 \IDinst/U10272  ( .DIN1(\IDinst/n10214 ), .DIN2(\IDinst/n10213 ), 
        .Q(\IDinst/n10215 ) );
  nnd2s1 \IDinst/U10271  ( .DIN1(\IDinst/n10212 ), .DIN2(n667), 
        .Q(\IDinst/n10214 ) );
  nnd2s1 \IDinst/U10270  ( .DIN1(\IDinst/n10191 ), .DIN2(n683), 
        .Q(\IDinst/n10213 ) );
  nnd2s1 \IDinst/U10269  ( .DIN1(\IDinst/n10211 ), .DIN2(\IDinst/n10210 ), 
        .Q(\IDinst/n10212 ) );
  nnd2s1 \IDinst/U10268  ( .DIN1(\IDinst/n10209 ), .DIN2(n1376), 
        .Q(\IDinst/n10211 ) );
  nnd2s1 \IDinst/U10267  ( .DIN1(\IDinst/n10200 ), .DIN2(n1367), 
        .Q(\IDinst/n10210 ) );
  nnd2s1 \IDinst/U10266  ( .DIN1(\IDinst/n10208 ), .DIN2(\IDinst/n10207 ), 
        .Q(\IDinst/n10209 ) );
  nnd2s1 \IDinst/U10265  ( .DIN1(\IDinst/n10206 ), .DIN2(n1330), 
        .Q(\IDinst/n10208 ) );
  nnd2s1 \IDinst/U10264  ( .DIN1(\IDinst/n10203 ), .DIN2(n1336), 
        .Q(\IDinst/n10207 ) );
  nnd2s1 \IDinst/U10263  ( .DIN1(\IDinst/n10205 ), .DIN2(\IDinst/n10204 ), 
        .Q(\IDinst/n10206 ) );
  nnd2s1 \IDinst/U10262  ( .DIN1(\IDinst/RegFile[31][13] ), .DIN2(n1230), 
        .Q(\IDinst/n10205 ) );
  nnd2s1 \IDinst/U10261  ( .DIN1(\IDinst/RegFile[30][13] ), .DIN2(n1248), 
        .Q(\IDinst/n10204 ) );
  nnd2s1 \IDinst/U10260  ( .DIN1(\IDinst/n10202 ), .DIN2(\IDinst/n10201 ), 
        .Q(\IDinst/n10203 ) );
  nnd2s1 \IDinst/U10259  ( .DIN1(\IDinst/RegFile[29][13] ), .DIN2(n1230), 
        .Q(\IDinst/n10202 ) );
  nnd2s1 \IDinst/U10258  ( .DIN1(\IDinst/RegFile[28][13] ), .DIN2(n1248), 
        .Q(\IDinst/n10201 ) );
  nnd2s1 \IDinst/U10257  ( .DIN1(\IDinst/n10199 ), .DIN2(\IDinst/n10198 ), 
        .Q(\IDinst/n10200 ) );
  nnd2s1 \IDinst/U10256  ( .DIN1(\IDinst/n10197 ), .DIN2(n1330), 
        .Q(\IDinst/n10199 ) );
  nnd2s1 \IDinst/U10255  ( .DIN1(\IDinst/n10194 ), .DIN2(n1336), 
        .Q(\IDinst/n10198 ) );
  nnd2s1 \IDinst/U10254  ( .DIN1(\IDinst/n10196 ), .DIN2(\IDinst/n10195 ), 
        .Q(\IDinst/n10197 ) );
  nnd2s1 \IDinst/U10253  ( .DIN1(\IDinst/RegFile[27][13] ), .DIN2(n1230), 
        .Q(\IDinst/n10196 ) );
  nnd2s1 \IDinst/U10252  ( .DIN1(\IDinst/RegFile[26][13] ), .DIN2(n1248), 
        .Q(\IDinst/n10195 ) );
  nnd2s1 \IDinst/U10251  ( .DIN1(\IDinst/n10193 ), .DIN2(\IDinst/n10192 ), 
        .Q(\IDinst/n10194 ) );
  nnd2s1 \IDinst/U10250  ( .DIN1(\IDinst/RegFile[25][13] ), .DIN2(n1230), 
        .Q(\IDinst/n10193 ) );
  nnd2s1 \IDinst/U10249  ( .DIN1(\IDinst/RegFile[24][13] ), .DIN2(n1248), 
        .Q(\IDinst/n10192 ) );
  nnd2s1 \IDinst/U10248  ( .DIN1(\IDinst/n10190 ), .DIN2(\IDinst/n10189 ), 
        .Q(\IDinst/n10191 ) );
  nnd2s1 \IDinst/U10247  ( .DIN1(\IDinst/n10188 ), .DIN2(n1376), 
        .Q(\IDinst/n10190 ) );
  nnd2s1 \IDinst/U10246  ( .DIN1(\IDinst/n10179 ), .DIN2(n1367), 
        .Q(\IDinst/n10189 ) );
  nnd2s1 \IDinst/U10245  ( .DIN1(\IDinst/n10187 ), .DIN2(\IDinst/n10186 ), 
        .Q(\IDinst/n10188 ) );
  nnd2s1 \IDinst/U10244  ( .DIN1(\IDinst/n10185 ), .DIN2(n1330), 
        .Q(\IDinst/n10187 ) );
  nnd2s1 \IDinst/U10243  ( .DIN1(\IDinst/n10182 ), .DIN2(n1336), 
        .Q(\IDinst/n10186 ) );
  nnd2s1 \IDinst/U10242  ( .DIN1(\IDinst/n10184 ), .DIN2(\IDinst/n10183 ), 
        .Q(\IDinst/n10185 ) );
  nnd2s1 \IDinst/U10241  ( .DIN1(\IDinst/RegFile[23][13] ), .DIN2(n1230), 
        .Q(\IDinst/n10184 ) );
  nnd2s1 \IDinst/U10240  ( .DIN1(\IDinst/RegFile[22][13] ), .DIN2(n1248), 
        .Q(\IDinst/n10183 ) );
  nnd2s1 \IDinst/U10239  ( .DIN1(\IDinst/n10181 ), .DIN2(\IDinst/n10180 ), 
        .Q(\IDinst/n10182 ) );
  nnd2s1 \IDinst/U10238  ( .DIN1(\IDinst/RegFile[21][13] ), .DIN2(n1231), 
        .Q(\IDinst/n10181 ) );
  nnd2s1 \IDinst/U10237  ( .DIN1(\IDinst/RegFile[20][13] ), .DIN2(n1247), 
        .Q(\IDinst/n10180 ) );
  nnd2s1 \IDinst/U10236  ( .DIN1(\IDinst/n10178 ), .DIN2(\IDinst/n10177 ), 
        .Q(\IDinst/n10179 ) );
  nnd2s1 \IDinst/U10235  ( .DIN1(\IDinst/n10176 ), .DIN2(n1330), 
        .Q(\IDinst/n10178 ) );
  nnd2s1 \IDinst/U10234  ( .DIN1(\IDinst/n10173 ), .DIN2(n1336), 
        .Q(\IDinst/n10177 ) );
  nnd2s1 \IDinst/U10233  ( .DIN1(\IDinst/n10175 ), .DIN2(\IDinst/n10174 ), 
        .Q(\IDinst/n10176 ) );
  nnd2s1 \IDinst/U10232  ( .DIN1(\IDinst/RegFile[19][13] ), .DIN2(n1231), 
        .Q(\IDinst/n10175 ) );
  nnd2s1 \IDinst/U10231  ( .DIN1(\IDinst/RegFile[18][13] ), .DIN2(n1247), 
        .Q(\IDinst/n10174 ) );
  nnd2s1 \IDinst/U10230  ( .DIN1(\IDinst/n10172 ), .DIN2(\IDinst/n10171 ), 
        .Q(\IDinst/n10173 ) );
  nnd2s1 \IDinst/U10229  ( .DIN1(\IDinst/RegFile[17][13] ), .DIN2(n1231), 
        .Q(\IDinst/n10172 ) );
  nnd2s1 \IDinst/U10228  ( .DIN1(\IDinst/RegFile[16][13] ), .DIN2(n1247), 
        .Q(\IDinst/n10171 ) );
  nnd2s1 \IDinst/U10227  ( .DIN1(\IDinst/n10169 ), .DIN2(\IDinst/n10168 ), 
        .Q(\IDinst/n10170 ) );
  nnd2s1 \IDinst/U10226  ( .DIN1(\IDinst/n10167 ), .DIN2(n665), 
        .Q(\IDinst/n10169 ) );
  nnd2s1 \IDinst/U10225  ( .DIN1(\IDinst/n10146 ), .DIN2(n682), 
        .Q(\IDinst/n10168 ) );
  nnd2s1 \IDinst/U10224  ( .DIN1(\IDinst/n10166 ), .DIN2(\IDinst/n10165 ), 
        .Q(\IDinst/n10167 ) );
  nnd2s1 \IDinst/U10223  ( .DIN1(\IDinst/n10164 ), .DIN2(n1376), 
        .Q(\IDinst/n10166 ) );
  nnd2s1 \IDinst/U10222  ( .DIN1(\IDinst/n10155 ), .DIN2(n1367), 
        .Q(\IDinst/n10165 ) );
  nnd2s1 \IDinst/U10221  ( .DIN1(\IDinst/n10163 ), .DIN2(\IDinst/n10162 ), 
        .Q(\IDinst/n10164 ) );
  nnd2s1 \IDinst/U10220  ( .DIN1(\IDinst/n10161 ), .DIN2(n1330), 
        .Q(\IDinst/n10163 ) );
  nnd2s1 \IDinst/U10219  ( .DIN1(\IDinst/n10158 ), .DIN2(n1336), 
        .Q(\IDinst/n10162 ) );
  nnd2s1 \IDinst/U10218  ( .DIN1(\IDinst/n10160 ), .DIN2(\IDinst/n10159 ), 
        .Q(\IDinst/n10161 ) );
  nnd2s1 \IDinst/U10217  ( .DIN1(\IDinst/RegFile[15][13] ), .DIN2(n1231), 
        .Q(\IDinst/n10160 ) );
  nnd2s1 \IDinst/U10216  ( .DIN1(\IDinst/RegFile[14][13] ), .DIN2(n1247), 
        .Q(\IDinst/n10159 ) );
  nnd2s1 \IDinst/U10215  ( .DIN1(\IDinst/n10157 ), .DIN2(\IDinst/n10156 ), 
        .Q(\IDinst/n10158 ) );
  nnd2s1 \IDinst/U10214  ( .DIN1(\IDinst/RegFile[13][13] ), .DIN2(n1231), 
        .Q(\IDinst/n10157 ) );
  nnd2s1 \IDinst/U10213  ( .DIN1(\IDinst/RegFile[12][13] ), .DIN2(n1247), 
        .Q(\IDinst/n10156 ) );
  nnd2s1 \IDinst/U10212  ( .DIN1(\IDinst/n10154 ), .DIN2(\IDinst/n10153 ), 
        .Q(\IDinst/n10155 ) );
  nnd2s1 \IDinst/U10211  ( .DIN1(\IDinst/n10152 ), .DIN2(n1330), 
        .Q(\IDinst/n10154 ) );
  nnd2s1 \IDinst/U10210  ( .DIN1(\IDinst/n10149 ), .DIN2(n1336), 
        .Q(\IDinst/n10153 ) );
  nnd2s1 \IDinst/U10209  ( .DIN1(\IDinst/n10151 ), .DIN2(\IDinst/n10150 ), 
        .Q(\IDinst/n10152 ) );
  nnd2s1 \IDinst/U10208  ( .DIN1(\IDinst/RegFile[11][13] ), .DIN2(n1231), 
        .Q(\IDinst/n10151 ) );
  nnd2s1 \IDinst/U10207  ( .DIN1(\IDinst/RegFile[10][13] ), .DIN2(n1247), 
        .Q(\IDinst/n10150 ) );
  nnd2s1 \IDinst/U10206  ( .DIN1(\IDinst/n10148 ), .DIN2(\IDinst/n10147 ), 
        .Q(\IDinst/n10149 ) );
  nnd2s1 \IDinst/U10205  ( .DIN1(\IDinst/RegFile[9][13] ), .DIN2(n1231), 
        .Q(\IDinst/n10148 ) );
  nnd2s1 \IDinst/U10204  ( .DIN1(\IDinst/RegFile[8][13] ), .DIN2(n1247), 
        .Q(\IDinst/n10147 ) );
  nnd2s1 \IDinst/U10203  ( .DIN1(\IDinst/n10145 ), .DIN2(\IDinst/n10144 ), 
        .Q(\IDinst/n10146 ) );
  nnd2s1 \IDinst/U10202  ( .DIN1(\IDinst/n10143 ), .DIN2(n1376), 
        .Q(\IDinst/n10145 ) );
  nnd2s1 \IDinst/U10201  ( .DIN1(\IDinst/n10134 ), .DIN2(n1367), 
        .Q(\IDinst/n10144 ) );
  nnd2s1 \IDinst/U10200  ( .DIN1(\IDinst/n10142 ), .DIN2(\IDinst/n10141 ), 
        .Q(\IDinst/n10143 ) );
  nnd2s1 \IDinst/U10199  ( .DIN1(\IDinst/n10140 ), .DIN2(n1330), 
        .Q(\IDinst/n10142 ) );
  nnd2s1 \IDinst/U10198  ( .DIN1(\IDinst/n10137 ), .DIN2(n1336), 
        .Q(\IDinst/n10141 ) );
  nnd2s1 \IDinst/U10197  ( .DIN1(\IDinst/n10139 ), .DIN2(\IDinst/n10138 ), 
        .Q(\IDinst/n10140 ) );
  nnd2s1 \IDinst/U10196  ( .DIN1(\IDinst/RegFile[7][13] ), .DIN2(n1231), 
        .Q(\IDinst/n10139 ) );
  nnd2s1 \IDinst/U10195  ( .DIN1(\IDinst/RegFile[6][13] ), .DIN2(n1247), 
        .Q(\IDinst/n10138 ) );
  nnd2s1 \IDinst/U10194  ( .DIN1(\IDinst/n10136 ), .DIN2(\IDinst/n10135 ), 
        .Q(\IDinst/n10137 ) );
  nnd2s1 \IDinst/U10193  ( .DIN1(\IDinst/RegFile[5][13] ), .DIN2(n1231), 
        .Q(\IDinst/n10136 ) );
  nnd2s1 \IDinst/U10192  ( .DIN1(\IDinst/RegFile[4][13] ), .DIN2(n1247), 
        .Q(\IDinst/n10135 ) );
  nnd2s1 \IDinst/U10191  ( .DIN1(\IDinst/n10133 ), .DIN2(\IDinst/n10132 ), 
        .Q(\IDinst/n10134 ) );
  nnd2s1 \IDinst/U10190  ( .DIN1(\IDinst/n10131 ), .DIN2(n1330), 
        .Q(\IDinst/n10133 ) );
  nnd2s1 \IDinst/U10189  ( .DIN1(\IDinst/n10128 ), .DIN2(n1336), 
        .Q(\IDinst/n10132 ) );
  nnd2s1 \IDinst/U10188  ( .DIN1(\IDinst/n10130 ), .DIN2(\IDinst/n10129 ), 
        .Q(\IDinst/n10131 ) );
  nnd2s1 \IDinst/U10187  ( .DIN1(\IDinst/RegFile[3][13] ), .DIN2(n1231), 
        .Q(\IDinst/n10130 ) );
  nnd2s1 \IDinst/U10186  ( .DIN1(\IDinst/RegFile[2][13] ), .DIN2(n1246), 
        .Q(\IDinst/n10129 ) );
  nnd2s1 \IDinst/U10185  ( .DIN1(\IDinst/n10127 ), .DIN2(\IDinst/n10126 ), 
        .Q(\IDinst/n10128 ) );
  nnd2s1 \IDinst/U10184  ( .DIN1(\IDinst/RegFile[1][13] ), .DIN2(n1231), 
        .Q(\IDinst/n10127 ) );
  nnd2s1 \IDinst/U10183  ( .DIN1(\IDinst/RegFile[0][13] ), .DIN2(n1246), 
        .Q(\IDinst/n10126 ) );
  nnd2s1 \IDinst/U10182  ( .DIN1(\IDinst/n10125 ), .DIN2(n535), 
        .Q(\IDinst/n8916 ) );
  nnd2s1 \IDinst/U10181  ( .DIN1(\IDinst/n10080 ), .DIN2(n634), 
        .Q(\IDinst/n8917 ) );
  nnd2s1 \IDinst/U10180  ( .DIN1(\IDinst/n10124 ), .DIN2(\IDinst/n10123 ), 
        .Q(\IDinst/n10125 ) );
  nnd2s1 \IDinst/U10179  ( .DIN1(\IDinst/n10122 ), .DIN2(n668), 
        .Q(\IDinst/n10124 ) );
  nnd2s1 \IDinst/U10178  ( .DIN1(\IDinst/n10101 ), .DIN2(n680), 
        .Q(\IDinst/n10123 ) );
  nnd2s1 \IDinst/U10177  ( .DIN1(\IDinst/n10121 ), .DIN2(\IDinst/n10120 ), 
        .Q(\IDinst/n10122 ) );
  nnd2s1 \IDinst/U10176  ( .DIN1(\IDinst/n10119 ), .DIN2(n1376), 
        .Q(\IDinst/n10121 ) );
  nnd2s1 \IDinst/U10175  ( .DIN1(\IDinst/n10110 ), .DIN2(n1367), 
        .Q(\IDinst/n10120 ) );
  nnd2s1 \IDinst/U10174  ( .DIN1(\IDinst/n10118 ), .DIN2(\IDinst/n10117 ), 
        .Q(\IDinst/n10119 ) );
  nnd2s1 \IDinst/U10173  ( .DIN1(\IDinst/n10116 ), .DIN2(n1330), 
        .Q(\IDinst/n10118 ) );
  nnd2s1 \IDinst/U10172  ( .DIN1(\IDinst/n10113 ), .DIN2(n1336), 
        .Q(\IDinst/n10117 ) );
  nnd2s1 \IDinst/U10171  ( .DIN1(\IDinst/n10115 ), .DIN2(\IDinst/n10114 ), 
        .Q(\IDinst/n10116 ) );
  nnd2s1 \IDinst/U10170  ( .DIN1(\IDinst/RegFile[31][12] ), .DIN2(n1231), 
        .Q(\IDinst/n10115 ) );
  nnd2s1 \IDinst/U10169  ( .DIN1(\IDinst/RegFile[30][12] ), .DIN2(n1246), 
        .Q(\IDinst/n10114 ) );
  nnd2s1 \IDinst/U10168  ( .DIN1(\IDinst/n10112 ), .DIN2(\IDinst/n10111 ), 
        .Q(\IDinst/n10113 ) );
  nnd2s1 \IDinst/U10167  ( .DIN1(\IDinst/RegFile[29][12] ), .DIN2(n1231), 
        .Q(\IDinst/n10112 ) );
  nnd2s1 \IDinst/U10166  ( .DIN1(\IDinst/RegFile[28][12] ), .DIN2(n1246), 
        .Q(\IDinst/n10111 ) );
  nnd2s1 \IDinst/U10165  ( .DIN1(\IDinst/n10109 ), .DIN2(\IDinst/n10108 ), 
        .Q(\IDinst/n10110 ) );
  nnd2s1 \IDinst/U10164  ( .DIN1(\IDinst/n10107 ), .DIN2(n1330), 
        .Q(\IDinst/n10109 ) );
  nnd2s1 \IDinst/U10163  ( .DIN1(\IDinst/n10104 ), .DIN2(n1337), 
        .Q(\IDinst/n10108 ) );
  nnd2s1 \IDinst/U10162  ( .DIN1(\IDinst/n10106 ), .DIN2(\IDinst/n10105 ), 
        .Q(\IDinst/n10107 ) );
  nnd2s1 \IDinst/U10161  ( .DIN1(\IDinst/RegFile[27][12] ), .DIN2(n1232), 
        .Q(\IDinst/n10106 ) );
  nnd2s1 \IDinst/U10160  ( .DIN1(\IDinst/RegFile[26][12] ), .DIN2(n1246), 
        .Q(\IDinst/n10105 ) );
  nnd2s1 \IDinst/U10159  ( .DIN1(\IDinst/n10103 ), .DIN2(\IDinst/n10102 ), 
        .Q(\IDinst/n10104 ) );
  nnd2s1 \IDinst/U10158  ( .DIN1(\IDinst/RegFile[25][12] ), .DIN2(n1232), 
        .Q(\IDinst/n10103 ) );
  nnd2s1 \IDinst/U10157  ( .DIN1(\IDinst/RegFile[24][12] ), .DIN2(n1246), 
        .Q(\IDinst/n10102 ) );
  nnd2s1 \IDinst/U10156  ( .DIN1(\IDinst/n10100 ), .DIN2(\IDinst/n10099 ), 
        .Q(\IDinst/n10101 ) );
  nnd2s1 \IDinst/U10155  ( .DIN1(\IDinst/n10098 ), .DIN2(n1376), 
        .Q(\IDinst/n10100 ) );
  nnd2s1 \IDinst/U10154  ( .DIN1(\IDinst/n10089 ), .DIN2(n1367), 
        .Q(\IDinst/n10099 ) );
  nnd2s1 \IDinst/U10153  ( .DIN1(\IDinst/n10097 ), .DIN2(\IDinst/n10096 ), 
        .Q(\IDinst/n10098 ) );
  nnd2s1 \IDinst/U10152  ( .DIN1(\IDinst/n10095 ), .DIN2(n1330), 
        .Q(\IDinst/n10097 ) );
  nnd2s1 \IDinst/U10151  ( .DIN1(\IDinst/n10092 ), .DIN2(n1337), 
        .Q(\IDinst/n10096 ) );
  nnd2s1 \IDinst/U10150  ( .DIN1(\IDinst/n10094 ), .DIN2(\IDinst/n10093 ), 
        .Q(\IDinst/n10095 ) );
  nnd2s1 \IDinst/U10149  ( .DIN1(\IDinst/RegFile[23][12] ), .DIN2(n1232), 
        .Q(\IDinst/n10094 ) );
  nnd2s1 \IDinst/U10148  ( .DIN1(\IDinst/RegFile[22][12] ), .DIN2(n1246), 
        .Q(\IDinst/n10093 ) );
  nnd2s1 \IDinst/U10147  ( .DIN1(\IDinst/n10091 ), .DIN2(\IDinst/n10090 ), 
        .Q(\IDinst/n10092 ) );
  nnd2s1 \IDinst/U10146  ( .DIN1(\IDinst/RegFile[21][12] ), .DIN2(n1232), 
        .Q(\IDinst/n10091 ) );
  nnd2s1 \IDinst/U10145  ( .DIN1(\IDinst/RegFile[20][12] ), .DIN2(n1246), 
        .Q(\IDinst/n10090 ) );
  nnd2s1 \IDinst/U10144  ( .DIN1(\IDinst/n10088 ), .DIN2(\IDinst/n10087 ), 
        .Q(\IDinst/n10089 ) );
  nnd2s1 \IDinst/U10143  ( .DIN1(\IDinst/n10086 ), .DIN2(n1330), 
        .Q(\IDinst/n10088 ) );
  nnd2s1 \IDinst/U10142  ( .DIN1(\IDinst/n10083 ), .DIN2(n1337), 
        .Q(\IDinst/n10087 ) );
  nnd2s1 \IDinst/U10141  ( .DIN1(\IDinst/n10085 ), .DIN2(\IDinst/n10084 ), 
        .Q(\IDinst/n10086 ) );
  nnd2s1 \IDinst/U10140  ( .DIN1(\IDinst/RegFile[19][12] ), .DIN2(n1232), 
        .Q(\IDinst/n10085 ) );
  nnd2s1 \IDinst/U10139  ( .DIN1(\IDinst/RegFile[18][12] ), .DIN2(n1245), 
        .Q(\IDinst/n10084 ) );
  nnd2s1 \IDinst/U10138  ( .DIN1(\IDinst/n10082 ), .DIN2(\IDinst/n10081 ), 
        .Q(\IDinst/n10083 ) );
  nnd2s1 \IDinst/U10137  ( .DIN1(\IDinst/RegFile[17][12] ), .DIN2(n1232), 
        .Q(\IDinst/n10082 ) );
  nnd2s1 \IDinst/U10136  ( .DIN1(\IDinst/RegFile[16][12] ), .DIN2(n1245), 
        .Q(\IDinst/n10081 ) );
  nnd2s1 \IDinst/U10135  ( .DIN1(\IDinst/n10079 ), .DIN2(\IDinst/n10078 ), 
        .Q(\IDinst/n10080 ) );
  nnd2s1 \IDinst/U10134  ( .DIN1(\IDinst/n10077 ), .DIN2(n666), 
        .Q(\IDinst/n10079 ) );
  nnd2s1 \IDinst/U10133  ( .DIN1(\IDinst/n10056 ), .DIN2(n681), 
        .Q(\IDinst/n10078 ) );
  nnd2s1 \IDinst/U10132  ( .DIN1(\IDinst/n10076 ), .DIN2(\IDinst/n10075 ), 
        .Q(\IDinst/n10077 ) );
  nnd2s1 \IDinst/U10131  ( .DIN1(\IDinst/n10074 ), .DIN2(n1376), 
        .Q(\IDinst/n10076 ) );
  nnd2s1 \IDinst/U10130  ( .DIN1(\IDinst/n10065 ), .DIN2(n1367), 
        .Q(\IDinst/n10075 ) );
  nnd2s1 \IDinst/U10129  ( .DIN1(\IDinst/n10073 ), .DIN2(\IDinst/n10072 ), 
        .Q(\IDinst/n10074 ) );
  nnd2s1 \IDinst/U10128  ( .DIN1(\IDinst/n10071 ), .DIN2(n1330), 
        .Q(\IDinst/n10073 ) );
  nnd2s1 \IDinst/U10127  ( .DIN1(\IDinst/n10068 ), .DIN2(n1337), 
        .Q(\IDinst/n10072 ) );
  nnd2s1 \IDinst/U10126  ( .DIN1(\IDinst/n10070 ), .DIN2(\IDinst/n10069 ), 
        .Q(\IDinst/n10071 ) );
  nnd2s1 \IDinst/U10125  ( .DIN1(\IDinst/RegFile[15][12] ), .DIN2(n1232), 
        .Q(\IDinst/n10070 ) );
  nnd2s1 \IDinst/U10124  ( .DIN1(\IDinst/RegFile[14][12] ), .DIN2(n1245), 
        .Q(\IDinst/n10069 ) );
  nnd2s1 \IDinst/U10123  ( .DIN1(\IDinst/n10067 ), .DIN2(\IDinst/n10066 ), 
        .Q(\IDinst/n10068 ) );
  nnd2s1 \IDinst/U10122  ( .DIN1(\IDinst/RegFile[13][12] ), .DIN2(n1232), 
        .Q(\IDinst/n10067 ) );
  nnd2s1 \IDinst/U10121  ( .DIN1(\IDinst/RegFile[12][12] ), .DIN2(n1245), 
        .Q(\IDinst/n10066 ) );
  nnd2s1 \IDinst/U10120  ( .DIN1(\IDinst/n10064 ), .DIN2(\IDinst/n10063 ), 
        .Q(\IDinst/n10065 ) );
  nnd2s1 \IDinst/U10119  ( .DIN1(\IDinst/n10062 ), .DIN2(n1329), 
        .Q(\IDinst/n10064 ) );
  nnd2s1 \IDinst/U10118  ( .DIN1(\IDinst/n10059 ), .DIN2(n1337), 
        .Q(\IDinst/n10063 ) );
  nnd2s1 \IDinst/U10117  ( .DIN1(\IDinst/n10061 ), .DIN2(\IDinst/n10060 ), 
        .Q(\IDinst/n10062 ) );
  nnd2s1 \IDinst/U10116  ( .DIN1(\IDinst/RegFile[11][12] ), .DIN2(n1232), 
        .Q(\IDinst/n10061 ) );
  nnd2s1 \IDinst/U10115  ( .DIN1(\IDinst/RegFile[10][12] ), .DIN2(n1245), 
        .Q(\IDinst/n10060 ) );
  nnd2s1 \IDinst/U10114  ( .DIN1(\IDinst/n10058 ), .DIN2(\IDinst/n10057 ), 
        .Q(\IDinst/n10059 ) );
  nnd2s1 \IDinst/U10113  ( .DIN1(\IDinst/RegFile[9][12] ), .DIN2(n1232), 
        .Q(\IDinst/n10058 ) );
  nnd2s1 \IDinst/U10112  ( .DIN1(\IDinst/RegFile[8][12] ), .DIN2(n1245), 
        .Q(\IDinst/n10057 ) );
  nnd2s1 \IDinst/U10111  ( .DIN1(\IDinst/n10055 ), .DIN2(\IDinst/n10054 ), 
        .Q(\IDinst/n10056 ) );
  nnd2s1 \IDinst/U10110  ( .DIN1(\IDinst/n10053 ), .DIN2(n1376), 
        .Q(\IDinst/n10055 ) );
  nnd2s1 \IDinst/U10109  ( .DIN1(\IDinst/n10044 ), .DIN2(n1367), 
        .Q(\IDinst/n10054 ) );
  nnd2s1 \IDinst/U10108  ( .DIN1(\IDinst/n10052 ), .DIN2(\IDinst/n10051 ), 
        .Q(\IDinst/n10053 ) );
  nnd2s1 \IDinst/U10107  ( .DIN1(\IDinst/n10050 ), .DIN2(n1329), 
        .Q(\IDinst/n10052 ) );
  nnd2s1 \IDinst/U10106  ( .DIN1(\IDinst/n10047 ), .DIN2(n1337), 
        .Q(\IDinst/n10051 ) );
  nnd2s1 \IDinst/U10105  ( .DIN1(\IDinst/n10049 ), .DIN2(\IDinst/n10048 ), 
        .Q(\IDinst/n10050 ) );
  nnd2s1 \IDinst/U10104  ( .DIN1(\IDinst/RegFile[7][12] ), .DIN2(n1232), 
        .Q(\IDinst/n10049 ) );
  nnd2s1 \IDinst/U10103  ( .DIN1(\IDinst/RegFile[6][12] ), .DIN2(n1245), 
        .Q(\IDinst/n10048 ) );
  nnd2s1 \IDinst/U10102  ( .DIN1(\IDinst/n10046 ), .DIN2(\IDinst/n10045 ), 
        .Q(\IDinst/n10047 ) );
  nnd2s1 \IDinst/U10101  ( .DIN1(\IDinst/RegFile[5][12] ), .DIN2(n1232), 
        .Q(\IDinst/n10046 ) );
  nnd2s1 \IDinst/U10100  ( .DIN1(\IDinst/RegFile[4][12] ), .DIN2(n1245), 
        .Q(\IDinst/n10045 ) );
  nnd2s1 \IDinst/U10099  ( .DIN1(\IDinst/n10043 ), .DIN2(\IDinst/n10042 ), 
        .Q(\IDinst/n10044 ) );
  nnd2s1 \IDinst/U10098  ( .DIN1(\IDinst/n10041 ), .DIN2(n1329), 
        .Q(\IDinst/n10043 ) );
  nnd2s1 \IDinst/U10097  ( .DIN1(\IDinst/n10038 ), .DIN2(n1337), 
        .Q(\IDinst/n10042 ) );
  nnd2s1 \IDinst/U10096  ( .DIN1(\IDinst/n10040 ), .DIN2(\IDinst/n10039 ), 
        .Q(\IDinst/n10041 ) );
  nnd2s1 \IDinst/U10095  ( .DIN1(\IDinst/RegFile[3][12] ), .DIN2(n1232), 
        .Q(\IDinst/n10040 ) );
  nnd2s1 \IDinst/U10094  ( .DIN1(\IDinst/RegFile[2][12] ), .DIN2(n1245), 
        .Q(\IDinst/n10039 ) );
  nnd2s1 \IDinst/U10093  ( .DIN1(\IDinst/n10037 ), .DIN2(\IDinst/n10036 ), 
        .Q(\IDinst/n10038 ) );
  nnd2s1 \IDinst/U10092  ( .DIN1(\IDinst/RegFile[1][12] ), .DIN2(n1233), 
        .Q(\IDinst/n10037 ) );
  nnd2s1 \IDinst/U10091  ( .DIN1(\IDinst/RegFile[0][12] ), .DIN2(n1244), 
        .Q(\IDinst/n10036 ) );
  nnd2s1 \IDinst/U10090  ( .DIN1(\IDinst/n10035 ), .DIN2(n534), 
        .Q(\IDinst/n8914 ) );
  nnd2s1 \IDinst/U10089  ( .DIN1(\IDinst/n9990 ), .DIN2(n533), 
        .Q(\IDinst/n8915 ) );
  nnd2s1 \IDinst/U10088  ( .DIN1(\IDinst/n10034 ), .DIN2(\IDinst/n10033 ), 
        .Q(\IDinst/n10035 ) );
  nnd2s1 \IDinst/U10087  ( .DIN1(\IDinst/n10032 ), .DIN2(n667), 
        .Q(\IDinst/n10034 ) );
  nnd2s1 \IDinst/U10086  ( .DIN1(\IDinst/n10011 ), .DIN2(n683), 
        .Q(\IDinst/n10033 ) );
  nnd2s1 \IDinst/U10085  ( .DIN1(\IDinst/n10031 ), .DIN2(\IDinst/n10030 ), 
        .Q(\IDinst/n10032 ) );
  nnd2s1 \IDinst/U10084  ( .DIN1(\IDinst/n10029 ), .DIN2(n1376), 
        .Q(\IDinst/n10031 ) );
  nnd2s1 \IDinst/U10083  ( .DIN1(\IDinst/n10020 ), .DIN2(n1367), 
        .Q(\IDinst/n10030 ) );
  nnd2s1 \IDinst/U10082  ( .DIN1(\IDinst/n10028 ), .DIN2(\IDinst/n10027 ), 
        .Q(\IDinst/n10029 ) );
  nnd2s1 \IDinst/U10081  ( .DIN1(\IDinst/n10026 ), .DIN2(n1329), 
        .Q(\IDinst/n10028 ) );
  nnd2s1 \IDinst/U10080  ( .DIN1(\IDinst/n10023 ), .DIN2(n1337), 
        .Q(\IDinst/n10027 ) );
  nnd2s1 \IDinst/U10079  ( .DIN1(\IDinst/n10025 ), .DIN2(\IDinst/n10024 ), 
        .Q(\IDinst/n10026 ) );
  nnd2s1 \IDinst/U10078  ( .DIN1(\IDinst/RegFile[31][11] ), .DIN2(n1233), 
        .Q(\IDinst/n10025 ) );
  nnd2s1 \IDinst/U10077  ( .DIN1(\IDinst/RegFile[30][11] ), .DIN2(n1244), 
        .Q(\IDinst/n10024 ) );
  nnd2s1 \IDinst/U10076  ( .DIN1(\IDinst/n10022 ), .DIN2(\IDinst/n10021 ), 
        .Q(\IDinst/n10023 ) );
  nnd2s1 \IDinst/U10075  ( .DIN1(\IDinst/RegFile[29][11] ), .DIN2(n1233), 
        .Q(\IDinst/n10022 ) );
  nnd2s1 \IDinst/U10074  ( .DIN1(\IDinst/RegFile[28][11] ), .DIN2(n1244), 
        .Q(\IDinst/n10021 ) );
  nnd2s1 \IDinst/U10073  ( .DIN1(\IDinst/n10019 ), .DIN2(\IDinst/n10018 ), 
        .Q(\IDinst/n10020 ) );
  nnd2s1 \IDinst/U10072  ( .DIN1(\IDinst/n10017 ), .DIN2(n1329), 
        .Q(\IDinst/n10019 ) );
  nnd2s1 \IDinst/U10071  ( .DIN1(\IDinst/n10014 ), .DIN2(n1337), 
        .Q(\IDinst/n10018 ) );
  nnd2s1 \IDinst/U10070  ( .DIN1(\IDinst/n10016 ), .DIN2(\IDinst/n10015 ), 
        .Q(\IDinst/n10017 ) );
  nnd2s1 \IDinst/U10069  ( .DIN1(\IDinst/RegFile[27][11] ), .DIN2(n1233), 
        .Q(\IDinst/n10016 ) );
  nnd2s1 \IDinst/U10068  ( .DIN1(\IDinst/RegFile[26][11] ), .DIN2(n1244), 
        .Q(\IDinst/n10015 ) );
  nnd2s1 \IDinst/U10067  ( .DIN1(\IDinst/n10013 ), .DIN2(\IDinst/n10012 ), 
        .Q(\IDinst/n10014 ) );
  nnd2s1 \IDinst/U10066  ( .DIN1(\IDinst/RegFile[25][11] ), .DIN2(n1233), 
        .Q(\IDinst/n10013 ) );
  nnd2s1 \IDinst/U10065  ( .DIN1(\IDinst/RegFile[24][11] ), .DIN2(n1244), 
        .Q(\IDinst/n10012 ) );
  nnd2s1 \IDinst/U10064  ( .DIN1(\IDinst/n10010 ), .DIN2(\IDinst/n10009 ), 
        .Q(\IDinst/n10011 ) );
  nnd2s1 \IDinst/U10063  ( .DIN1(\IDinst/n10008 ), .DIN2(n1377), 
        .Q(\IDinst/n10010 ) );
  nnd2s1 \IDinst/U10062  ( .DIN1(\IDinst/n9999 ), .DIN2(n1367), 
        .Q(\IDinst/n10009 ) );
  nnd2s1 \IDinst/U10061  ( .DIN1(\IDinst/n10007 ), .DIN2(\IDinst/n10006 ), 
        .Q(\IDinst/n10008 ) );
  nnd2s1 \IDinst/U10060  ( .DIN1(\IDinst/n10005 ), .DIN2(n1329), 
        .Q(\IDinst/n10007 ) );
  nnd2s1 \IDinst/U10059  ( .DIN1(\IDinst/n10002 ), .DIN2(n1338), 
        .Q(\IDinst/n10006 ) );
  nnd2s1 \IDinst/U10058  ( .DIN1(\IDinst/n10004 ), .DIN2(\IDinst/n10003 ), 
        .Q(\IDinst/n10005 ) );
  nnd2s1 \IDinst/U10057  ( .DIN1(\IDinst/RegFile[23][11] ), .DIN2(n1233), 
        .Q(\IDinst/n10004 ) );
  nnd2s1 \IDinst/U10056  ( .DIN1(\IDinst/RegFile[22][11] ), .DIN2(n1244), 
        .Q(\IDinst/n10003 ) );
  nnd2s1 \IDinst/U10055  ( .DIN1(\IDinst/n10001 ), .DIN2(\IDinst/n10000 ), 
        .Q(\IDinst/n10002 ) );
  nnd2s1 \IDinst/U10054  ( .DIN1(\IDinst/RegFile[21][11] ), .DIN2(n1233), 
        .Q(\IDinst/n10001 ) );
  nnd2s1 \IDinst/U10053  ( .DIN1(\IDinst/RegFile[20][11] ), .DIN2(n1244), 
        .Q(\IDinst/n10000 ) );
  nnd2s1 \IDinst/U10052  ( .DIN1(\IDinst/n9998 ), .DIN2(\IDinst/n9997 ), 
        .Q(\IDinst/n9999 ) );
  nnd2s1 \IDinst/U10051  ( .DIN1(\IDinst/n9996 ), .DIN2(n1329), 
        .Q(\IDinst/n9998 ) );
  nnd2s1 \IDinst/U10050  ( .DIN1(\IDinst/n9993 ), .DIN2(n1338), 
        .Q(\IDinst/n9997 ) );
  nnd2s1 \IDinst/U10049  ( .DIN1(\IDinst/n9995 ), .DIN2(\IDinst/n9994 ), 
        .Q(\IDinst/n9996 ) );
  nnd2s1 \IDinst/U10048  ( .DIN1(\IDinst/RegFile[19][11] ), .DIN2(n1233), 
        .Q(\IDinst/n9995 ) );
  nnd2s1 \IDinst/U10047  ( .DIN1(\IDinst/RegFile[18][11] ), .DIN2(n1244), 
        .Q(\IDinst/n9994 ) );
  nnd2s1 \IDinst/U10046  ( .DIN1(\IDinst/n9992 ), .DIN2(\IDinst/n9991 ), 
        .Q(\IDinst/n9993 ) );
  nnd2s1 \IDinst/U10045  ( .DIN1(\IDinst/RegFile[17][11] ), .DIN2(n1233), 
        .Q(\IDinst/n9992 ) );
  nnd2s1 \IDinst/U10044  ( .DIN1(\IDinst/RegFile[16][11] ), .DIN2(n1244), 
        .Q(\IDinst/n9991 ) );
  nnd2s1 \IDinst/U10043  ( .DIN1(\IDinst/n9989 ), .DIN2(\IDinst/n9988 ), 
        .Q(\IDinst/n9990 ) );
  nnd2s1 \IDinst/U10042  ( .DIN1(\IDinst/n9987 ), .DIN2(n665), 
        .Q(\IDinst/n9989 ) );
  nnd2s1 \IDinst/U10041  ( .DIN1(\IDinst/n9966 ), .DIN2(n682), 
        .Q(\IDinst/n9988 ) );
  nnd2s1 \IDinst/U10040  ( .DIN1(\IDinst/n9986 ), .DIN2(\IDinst/n9985 ), 
        .Q(\IDinst/n9987 ) );
  nnd2s1 \IDinst/U10039  ( .DIN1(\IDinst/n9984 ), .DIN2(n1377), 
        .Q(\IDinst/n9986 ) );
  nnd2s1 \IDinst/U10038  ( .DIN1(\IDinst/n9975 ), .DIN2(n1367), 
        .Q(\IDinst/n9985 ) );
  nnd2s1 \IDinst/U10037  ( .DIN1(\IDinst/n9983 ), .DIN2(\IDinst/n9982 ), 
        .Q(\IDinst/n9984 ) );
  nnd2s1 \IDinst/U10036  ( .DIN1(\IDinst/n9981 ), .DIN2(n1329), 
        .Q(\IDinst/n9983 ) );
  nnd2s1 \IDinst/U10035  ( .DIN1(\IDinst/n9978 ), .DIN2(n1338), 
        .Q(\IDinst/n9982 ) );
  nnd2s1 \IDinst/U10034  ( .DIN1(\IDinst/n9980 ), .DIN2(\IDinst/n9979 ), 
        .Q(\IDinst/n9981 ) );
  nnd2s1 \IDinst/U10033  ( .DIN1(\IDinst/RegFile[15][11] ), .DIN2(n1233), 
        .Q(\IDinst/n9980 ) );
  nnd2s1 \IDinst/U10032  ( .DIN1(\IDinst/RegFile[14][11] ), .DIN2(n1243), 
        .Q(\IDinst/n9979 ) );
  nnd2s1 \IDinst/U10031  ( .DIN1(\IDinst/n9977 ), .DIN2(\IDinst/n9976 ), 
        .Q(\IDinst/n9978 ) );
  nnd2s1 \IDinst/U10030  ( .DIN1(\IDinst/RegFile[13][11] ), .DIN2(n1233), 
        .Q(\IDinst/n9977 ) );
  nnd2s1 \IDinst/U10029  ( .DIN1(\IDinst/RegFile[12][11] ), .DIN2(n1243), 
        .Q(\IDinst/n9976 ) );
  nnd2s1 \IDinst/U10028  ( .DIN1(\IDinst/n9974 ), .DIN2(\IDinst/n9973 ), 
        .Q(\IDinst/n9975 ) );
  nnd2s1 \IDinst/U10027  ( .DIN1(\IDinst/n9972 ), .DIN2(n1329), 
        .Q(\IDinst/n9974 ) );
  nnd2s1 \IDinst/U10026  ( .DIN1(\IDinst/n9969 ), .DIN2(n1338), 
        .Q(\IDinst/n9973 ) );
  nnd2s1 \IDinst/U10025  ( .DIN1(\IDinst/n9971 ), .DIN2(\IDinst/n9970 ), 
        .Q(\IDinst/n9972 ) );
  nnd2s1 \IDinst/U10024  ( .DIN1(\IDinst/RegFile[11][11] ), .DIN2(n1233), 
        .Q(\IDinst/n9971 ) );
  nnd2s1 \IDinst/U10023  ( .DIN1(\IDinst/RegFile[10][11] ), .DIN2(n1243), 
        .Q(\IDinst/n9970 ) );
  nnd2s1 \IDinst/U10022  ( .DIN1(\IDinst/n9968 ), .DIN2(\IDinst/n9967 ), 
        .Q(\IDinst/n9969 ) );
  nnd2s1 \IDinst/U10021  ( .DIN1(\IDinst/RegFile[9][11] ), .DIN2(n1234), 
        .Q(\IDinst/n9968 ) );
  nnd2s1 \IDinst/U10020  ( .DIN1(\IDinst/RegFile[8][11] ), .DIN2(n1243), 
        .Q(\IDinst/n9967 ) );
  nnd2s1 \IDinst/U10019  ( .DIN1(\IDinst/n9965 ), .DIN2(\IDinst/n9964 ), 
        .Q(\IDinst/n9966 ) );
  nnd2s1 \IDinst/U10018  ( .DIN1(\IDinst/n9963 ), .DIN2(n1377), 
        .Q(\IDinst/n9965 ) );
  nnd2s1 \IDinst/U10017  ( .DIN1(\IDinst/n9954 ), .DIN2(n1367), 
        .Q(\IDinst/n9964 ) );
  nnd2s1 \IDinst/U10016  ( .DIN1(\IDinst/n9962 ), .DIN2(\IDinst/n9961 ), 
        .Q(\IDinst/n9963 ) );
  nnd2s1 \IDinst/U10015  ( .DIN1(\IDinst/n9960 ), .DIN2(n1329), 
        .Q(\IDinst/n9962 ) );
  nnd2s1 \IDinst/U10014  ( .DIN1(\IDinst/n9957 ), .DIN2(n1338), 
        .Q(\IDinst/n9961 ) );
  nnd2s1 \IDinst/U10013  ( .DIN1(\IDinst/n9959 ), .DIN2(\IDinst/n9958 ), 
        .Q(\IDinst/n9960 ) );
  nnd2s1 \IDinst/U10012  ( .DIN1(\IDinst/RegFile[7][11] ), .DIN2(n1234), 
        .Q(\IDinst/n9959 ) );
  nnd2s1 \IDinst/U10011  ( .DIN1(\IDinst/RegFile[6][11] ), .DIN2(n1243), 
        .Q(\IDinst/n9958 ) );
  nnd2s1 \IDinst/U10010  ( .DIN1(\IDinst/n9956 ), .DIN2(\IDinst/n9955 ), 
        .Q(\IDinst/n9957 ) );
  nnd2s1 \IDinst/U10009  ( .DIN1(\IDinst/RegFile[5][11] ), .DIN2(n1234), 
        .Q(\IDinst/n9956 ) );
  nnd2s1 \IDinst/U10008  ( .DIN1(\IDinst/RegFile[4][11] ), .DIN2(n1243), 
        .Q(\IDinst/n9955 ) );
  nnd2s1 \IDinst/U10007  ( .DIN1(\IDinst/n9953 ), .DIN2(\IDinst/n9952 ), 
        .Q(\IDinst/n9954 ) );
  nnd2s1 \IDinst/U10006  ( .DIN1(\IDinst/n9951 ), .DIN2(n1329), 
        .Q(\IDinst/n9953 ) );
  nnd2s1 \IDinst/U10005  ( .DIN1(\IDinst/n9948 ), .DIN2(n1338), 
        .Q(\IDinst/n9952 ) );
  nnd2s1 \IDinst/U10004  ( .DIN1(\IDinst/n9950 ), .DIN2(\IDinst/n9949 ), 
        .Q(\IDinst/n9951 ) );
  nnd2s1 \IDinst/U10003  ( .DIN1(\IDinst/RegFile[3][11] ), .DIN2(n1234), 
        .Q(\IDinst/n9950 ) );
  nnd2s1 \IDinst/U10002  ( .DIN1(\IDinst/RegFile[2][11] ), .DIN2(n1243), 
        .Q(\IDinst/n9949 ) );
  nnd2s1 \IDinst/U10001  ( .DIN1(\IDinst/n9947 ), .DIN2(\IDinst/n9946 ), 
        .Q(\IDinst/n9948 ) );
  nnd2s1 \IDinst/U10000  ( .DIN1(\IDinst/RegFile[1][11] ), .DIN2(n1234), 
        .Q(\IDinst/n9947 ) );
  nnd2s1 \IDinst/U9999  ( .DIN1(\IDinst/RegFile[0][11] ), .DIN2(n1243), 
        .Q(\IDinst/n9946 ) );
  nnd2s1 \IDinst/U9998  ( .DIN1(\IDinst/n9945 ), .DIN2(\IDinst/N48 ), 
        .Q(\IDinst/n8912 ) );
  nnd2s1 \IDinst/U9997  ( .DIN1(\IDinst/n9900 ), .DIN2(n634), 
        .Q(\IDinst/n8913 ) );
  nnd2s1 \IDinst/U9996  ( .DIN1(\IDinst/n9944 ), .DIN2(\IDinst/n9943 ), 
        .Q(\IDinst/n9945 ) );
  nnd2s1 \IDinst/U9995  ( .DIN1(\IDinst/n9942 ), .DIN2(n668), 
        .Q(\IDinst/n9944 ) );
  nnd2s1 \IDinst/U9994  ( .DIN1(\IDinst/n9921 ), .DIN2(n680), 
        .Q(\IDinst/n9943 ) );
  nnd2s1 \IDinst/U9993  ( .DIN1(\IDinst/n9941 ), .DIN2(\IDinst/n9940 ), 
        .Q(\IDinst/n9942 ) );
  nnd2s1 \IDinst/U9992  ( .DIN1(\IDinst/n9939 ), .DIN2(n1377), 
        .Q(\IDinst/n9941 ) );
  nnd2s1 \IDinst/U9991  ( .DIN1(\IDinst/n9930 ), .DIN2(n1367), 
        .Q(\IDinst/n9940 ) );
  nnd2s1 \IDinst/U9990  ( .DIN1(\IDinst/n9938 ), .DIN2(\IDinst/n9937 ), 
        .Q(\IDinst/n9939 ) );
  nnd2s1 \IDinst/U9989  ( .DIN1(\IDinst/n9936 ), .DIN2(n1329), 
        .Q(\IDinst/n9938 ) );
  nnd2s1 \IDinst/U9988  ( .DIN1(\IDinst/n9933 ), .DIN2(n1338), 
        .Q(\IDinst/n9937 ) );
  nnd2s1 \IDinst/U9987  ( .DIN1(\IDinst/n9935 ), .DIN2(\IDinst/n9934 ), 
        .Q(\IDinst/n9936 ) );
  nnd2s1 \IDinst/U9986  ( .DIN1(\IDinst/RegFile[31][10] ), .DIN2(n1234), 
        .Q(\IDinst/n9935 ) );
  nnd2s1 \IDinst/U9985  ( .DIN1(\IDinst/RegFile[30][10] ), .DIN2(n1242), 
        .Q(\IDinst/n9934 ) );
  nnd2s1 \IDinst/U9984  ( .DIN1(\IDinst/n9932 ), .DIN2(\IDinst/n9931 ), 
        .Q(\IDinst/n9933 ) );
  nnd2s1 \IDinst/U9983  ( .DIN1(\IDinst/RegFile[29][10] ), .DIN2(n1234), 
        .Q(\IDinst/n9932 ) );
  nnd2s1 \IDinst/U9982  ( .DIN1(\IDinst/RegFile[28][10] ), .DIN2(n1242), 
        .Q(\IDinst/n9931 ) );
  nnd2s1 \IDinst/U9981  ( .DIN1(\IDinst/n9929 ), .DIN2(\IDinst/n9928 ), 
        .Q(\IDinst/n9930 ) );
  nnd2s1 \IDinst/U9980  ( .DIN1(\IDinst/n9927 ), .DIN2(n1329), 
        .Q(\IDinst/n9929 ) );
  nnd2s1 \IDinst/U9979  ( .DIN1(\IDinst/n9924 ), .DIN2(n1338), 
        .Q(\IDinst/n9928 ) );
  nnd2s1 \IDinst/U9978  ( .DIN1(\IDinst/n9926 ), .DIN2(\IDinst/n9925 ), 
        .Q(\IDinst/n9927 ) );
  nnd2s1 \IDinst/U9977  ( .DIN1(\IDinst/RegFile[27][10] ), .DIN2(n1234), 
        .Q(\IDinst/n9926 ) );
  nnd2s1 \IDinst/U9976  ( .DIN1(\IDinst/RegFile[26][10] ), .DIN2(n1242), 
        .Q(\IDinst/n9925 ) );
  nnd2s1 \IDinst/U9975  ( .DIN1(\IDinst/n9923 ), .DIN2(\IDinst/n9922 ), 
        .Q(\IDinst/n9924 ) );
  nnd2s1 \IDinst/U9974  ( .DIN1(\IDinst/RegFile[25][10] ), .DIN2(n1234), 
        .Q(\IDinst/n9923 ) );
  nnd2s1 \IDinst/U9973  ( .DIN1(\IDinst/RegFile[24][10] ), .DIN2(n1242), 
        .Q(\IDinst/n9922 ) );
  nnd2s1 \IDinst/U9972  ( .DIN1(\IDinst/n9920 ), .DIN2(\IDinst/n9919 ), 
        .Q(\IDinst/n9921 ) );
  nnd2s1 \IDinst/U9971  ( .DIN1(\IDinst/n9918 ), .DIN2(n1377), 
        .Q(\IDinst/n9920 ) );
  nnd2s1 \IDinst/U9970  ( .DIN1(\IDinst/n9909 ), .DIN2(n1366), 
        .Q(\IDinst/n9919 ) );
  nnd2s1 \IDinst/U9969  ( .DIN1(\IDinst/n9917 ), .DIN2(\IDinst/n9916 ), 
        .Q(\IDinst/n9918 ) );
  nnd2s1 \IDinst/U9968  ( .DIN1(\IDinst/n9915 ), .DIN2(n1328), 
        .Q(\IDinst/n9917 ) );
  nnd2s1 \IDinst/U9967  ( .DIN1(\IDinst/n9912 ), .DIN2(n1338), 
        .Q(\IDinst/n9916 ) );
  nnd2s1 \IDinst/U9966  ( .DIN1(\IDinst/n9914 ), .DIN2(\IDinst/n9913 ), 
        .Q(\IDinst/n9915 ) );
  nnd2s1 \IDinst/U9965  ( .DIN1(\IDinst/RegFile[23][10] ), .DIN2(n1234), 
        .Q(\IDinst/n9914 ) );
  nnd2s1 \IDinst/U9964  ( .DIN1(\IDinst/RegFile[22][10] ), .DIN2(n1242), 
        .Q(\IDinst/n9913 ) );
  nnd2s1 \IDinst/U9963  ( .DIN1(\IDinst/n9911 ), .DIN2(\IDinst/n9910 ), 
        .Q(\IDinst/n9912 ) );
  nnd2s1 \IDinst/U9962  ( .DIN1(\IDinst/RegFile[21][10] ), .DIN2(n1234), 
        .Q(\IDinst/n9911 ) );
  nnd2s1 \IDinst/U9961  ( .DIN1(\IDinst/RegFile[20][10] ), .DIN2(n1242), 
        .Q(\IDinst/n9910 ) );
  nnd2s1 \IDinst/U9960  ( .DIN1(\IDinst/n9908 ), .DIN2(\IDinst/n9907 ), 
        .Q(\IDinst/n9909 ) );
  nnd2s1 \IDinst/U9959  ( .DIN1(\IDinst/n9906 ), .DIN2(n1328), 
        .Q(\IDinst/n9908 ) );
  nnd2s1 \IDinst/U9958  ( .DIN1(\IDinst/n9903 ), .DIN2(n1339), 
        .Q(\IDinst/n9907 ) );
  nnd2s1 \IDinst/U9957  ( .DIN1(\IDinst/n9905 ), .DIN2(\IDinst/n9904 ), 
        .Q(\IDinst/n9906 ) );
  nnd2s1 \IDinst/U9956  ( .DIN1(\IDinst/RegFile[19][10] ), .DIN2(n1234), 
        .Q(\IDinst/n9905 ) );
  nnd2s1 \IDinst/U9955  ( .DIN1(\IDinst/RegFile[18][10] ), .DIN2(n1242), 
        .Q(\IDinst/n9904 ) );
  nnd2s1 \IDinst/U9954  ( .DIN1(\IDinst/n9902 ), .DIN2(\IDinst/n9901 ), 
        .Q(\IDinst/n9903 ) );
  nnd2s1 \IDinst/U9953  ( .DIN1(\IDinst/RegFile[17][10] ), .DIN2(n1234), 
        .Q(\IDinst/n9902 ) );
  nnd2s1 \IDinst/U9952  ( .DIN1(\IDinst/RegFile[16][10] ), .DIN2(n1242), 
        .Q(\IDinst/n9901 ) );
  nnd2s1 \IDinst/U9951  ( .DIN1(\IDinst/n9899 ), .DIN2(\IDinst/n9898 ), 
        .Q(\IDinst/n9900 ) );
  nnd2s1 \IDinst/U9950  ( .DIN1(\IDinst/n9897 ), .DIN2(n666), 
        .Q(\IDinst/n9899 ) );
  nnd2s1 \IDinst/U9949  ( .DIN1(\IDinst/n9876 ), .DIN2(n681), 
        .Q(\IDinst/n9898 ) );
  nnd2s1 \IDinst/U9948  ( .DIN1(\IDinst/n9896 ), .DIN2(\IDinst/n9895 ), 
        .Q(\IDinst/n9897 ) );
  nnd2s1 \IDinst/U9947  ( .DIN1(\IDinst/n9894 ), .DIN2(n1377), 
        .Q(\IDinst/n9896 ) );
  nnd2s1 \IDinst/U9946  ( .DIN1(\IDinst/n9885 ), .DIN2(n1366), 
        .Q(\IDinst/n9895 ) );
  nnd2s1 \IDinst/U9945  ( .DIN1(\IDinst/n9893 ), .DIN2(\IDinst/n9892 ), 
        .Q(\IDinst/n9894 ) );
  nnd2s1 \IDinst/U9944  ( .DIN1(\IDinst/n9891 ), .DIN2(n1328), 
        .Q(\IDinst/n9893 ) );
  nnd2s1 \IDinst/U9943  ( .DIN1(\IDinst/n9888 ), .DIN2(n1339), 
        .Q(\IDinst/n9892 ) );
  nnd2s1 \IDinst/U9942  ( .DIN1(\IDinst/n9890 ), .DIN2(\IDinst/n9889 ), 
        .Q(\IDinst/n9891 ) );
  nnd2s1 \IDinst/U9941  ( .DIN1(\IDinst/RegFile[15][10] ), .DIN2(n1235), 
        .Q(\IDinst/n9890 ) );
  nnd2s1 \IDinst/U9940  ( .DIN1(\IDinst/RegFile[14][10] ), .DIN2(n1242), 
        .Q(\IDinst/n9889 ) );
  nnd2s1 \IDinst/U9939  ( .DIN1(\IDinst/n9887 ), .DIN2(\IDinst/n9886 ), 
        .Q(\IDinst/n9888 ) );
  nnd2s1 \IDinst/U9938  ( .DIN1(\IDinst/RegFile[13][10] ), .DIN2(n1235), 
        .Q(\IDinst/n9887 ) );
  nnd2s1 \IDinst/U9937  ( .DIN1(\IDinst/RegFile[12][10] ), .DIN2(n1243), 
        .Q(\IDinst/n9886 ) );
  nnd2s1 \IDinst/U9936  ( .DIN1(\IDinst/n9884 ), .DIN2(\IDinst/n9883 ), 
        .Q(\IDinst/n9885 ) );
  nnd2s1 \IDinst/U9935  ( .DIN1(\IDinst/n9882 ), .DIN2(n1328), 
        .Q(\IDinst/n9884 ) );
  nnd2s1 \IDinst/U9934  ( .DIN1(\IDinst/n9879 ), .DIN2(n1339), 
        .Q(\IDinst/n9883 ) );
  nnd2s1 \IDinst/U9933  ( .DIN1(\IDinst/n9881 ), .DIN2(\IDinst/n9880 ), 
        .Q(\IDinst/n9882 ) );
  nnd2s1 \IDinst/U9932  ( .DIN1(\IDinst/RegFile[11][10] ), .DIN2(n1235), 
        .Q(\IDinst/n9881 ) );
  nnd2s1 \IDinst/U9931  ( .DIN1(\IDinst/RegFile[10][10] ), .DIN2(n1241), 
        .Q(\IDinst/n9880 ) );
  nnd2s1 \IDinst/U9930  ( .DIN1(\IDinst/n9878 ), .DIN2(\IDinst/n9877 ), 
        .Q(\IDinst/n9879 ) );
  nnd2s1 \IDinst/U9929  ( .DIN1(\IDinst/RegFile[9][10] ), .DIN2(n1235), 
        .Q(\IDinst/n9878 ) );
  nnd2s1 \IDinst/U9928  ( .DIN1(\IDinst/RegFile[8][10] ), .DIN2(n1241), 
        .Q(\IDinst/n9877 ) );
  nnd2s1 \IDinst/U9927  ( .DIN1(\IDinst/n9875 ), .DIN2(\IDinst/n9874 ), 
        .Q(\IDinst/n9876 ) );
  nnd2s1 \IDinst/U9926  ( .DIN1(\IDinst/n9873 ), .DIN2(n1377), 
        .Q(\IDinst/n9875 ) );
  nnd2s1 \IDinst/U9925  ( .DIN1(\IDinst/n9864 ), .DIN2(n1366), 
        .Q(\IDinst/n9874 ) );
  nnd2s1 \IDinst/U9924  ( .DIN1(\IDinst/n9872 ), .DIN2(\IDinst/n9871 ), 
        .Q(\IDinst/n9873 ) );
  nnd2s1 \IDinst/U9923  ( .DIN1(\IDinst/n9870 ), .DIN2(n1328), 
        .Q(\IDinst/n9872 ) );
  nnd2s1 \IDinst/U9922  ( .DIN1(\IDinst/n9867 ), .DIN2(n1339), 
        .Q(\IDinst/n9871 ) );
  nnd2s1 \IDinst/U9921  ( .DIN1(\IDinst/n9869 ), .DIN2(\IDinst/n9868 ), 
        .Q(\IDinst/n9870 ) );
  nnd2s1 \IDinst/U9920  ( .DIN1(\IDinst/RegFile[7][10] ), .DIN2(n1235), 
        .Q(\IDinst/n9869 ) );
  nnd2s1 \IDinst/U9919  ( .DIN1(\IDinst/RegFile[6][10] ), .DIN2(n1241), 
        .Q(\IDinst/n9868 ) );
  nnd2s1 \IDinst/U9918  ( .DIN1(\IDinst/n9866 ), .DIN2(\IDinst/n9865 ), 
        .Q(\IDinst/n9867 ) );
  nnd2s1 \IDinst/U9917  ( .DIN1(\IDinst/RegFile[5][10] ), .DIN2(n1235), 
        .Q(\IDinst/n9866 ) );
  nnd2s1 \IDinst/U9916  ( .DIN1(\IDinst/RegFile[4][10] ), .DIN2(n1241), 
        .Q(\IDinst/n9865 ) );
  nnd2s1 \IDinst/U9915  ( .DIN1(\IDinst/n9863 ), .DIN2(\IDinst/n9862 ), 
        .Q(\IDinst/n9864 ) );
  nnd2s1 \IDinst/U9914  ( .DIN1(\IDinst/n9861 ), .DIN2(n1328), 
        .Q(\IDinst/n9863 ) );
  nnd2s1 \IDinst/U9913  ( .DIN1(\IDinst/n9858 ), .DIN2(n1339), 
        .Q(\IDinst/n9862 ) );
  nnd2s1 \IDinst/U9912  ( .DIN1(\IDinst/n9860 ), .DIN2(\IDinst/n9859 ), 
        .Q(\IDinst/n9861 ) );
  nnd2s1 \IDinst/U9911  ( .DIN1(\IDinst/RegFile[3][10] ), .DIN2(n1235), 
        .Q(\IDinst/n9860 ) );
  nnd2s1 \IDinst/U9910  ( .DIN1(\IDinst/RegFile[2][10] ), .DIN2(n1241), 
        .Q(\IDinst/n9859 ) );
  nnd2s1 \IDinst/U9909  ( .DIN1(\IDinst/n9857 ), .DIN2(\IDinst/n9856 ), 
        .Q(\IDinst/n9858 ) );
  nnd2s1 \IDinst/U9908  ( .DIN1(\IDinst/RegFile[1][10] ), .DIN2(n1235), 
        .Q(\IDinst/n9857 ) );
  nnd2s1 \IDinst/U9907  ( .DIN1(\IDinst/RegFile[0][10] ), .DIN2(n1241), 
        .Q(\IDinst/n9856 ) );
  nnd2s1 \IDinst/U9906  ( .DIN1(\IDinst/n9855 ), .DIN2(n535), 
        .Q(\IDinst/n8910 ) );
  nnd2s1 \IDinst/U9905  ( .DIN1(\IDinst/n9810 ), .DIN2(n533), 
        .Q(\IDinst/n8911 ) );
  nnd2s1 \IDinst/U9904  ( .DIN1(\IDinst/n9854 ), .DIN2(\IDinst/n9853 ), 
        .Q(\IDinst/n9855 ) );
  nnd2s1 \IDinst/U9903  ( .DIN1(\IDinst/n9852 ), .DIN2(n667), 
        .Q(\IDinst/n9854 ) );
  nnd2s1 \IDinst/U9902  ( .DIN1(\IDinst/n9831 ), .DIN2(n683), 
        .Q(\IDinst/n9853 ) );
  nnd2s1 \IDinst/U9901  ( .DIN1(\IDinst/n9851 ), .DIN2(\IDinst/n9850 ), 
        .Q(\IDinst/n9852 ) );
  nnd2s1 \IDinst/U9900  ( .DIN1(\IDinst/n9849 ), .DIN2(n1377), 
        .Q(\IDinst/n9851 ) );
  nnd2s1 \IDinst/U9899  ( .DIN1(\IDinst/n9840 ), .DIN2(n1366), 
        .Q(\IDinst/n9850 ) );
  nnd2s1 \IDinst/U9898  ( .DIN1(\IDinst/n9848 ), .DIN2(\IDinst/n9847 ), 
        .Q(\IDinst/n9849 ) );
  nnd2s1 \IDinst/U9897  ( .DIN1(\IDinst/n9846 ), .DIN2(n1328), 
        .Q(\IDinst/n9848 ) );
  nnd2s1 \IDinst/U9896  ( .DIN1(\IDinst/n9843 ), .DIN2(n1339), 
        .Q(\IDinst/n9847 ) );
  nnd2s1 \IDinst/U9895  ( .DIN1(\IDinst/n9845 ), .DIN2(\IDinst/n9844 ), 
        .Q(\IDinst/n9846 ) );
  nnd2s1 \IDinst/U9894  ( .DIN1(\IDinst/RegFile[31][9] ), .DIN2(n1235), 
        .Q(\IDinst/n9845 ) );
  nnd2s1 \IDinst/U9893  ( .DIN1(\IDinst/RegFile[30][9] ), .DIN2(n1241), 
        .Q(\IDinst/n9844 ) );
  nnd2s1 \IDinst/U9892  ( .DIN1(\IDinst/n9842 ), .DIN2(\IDinst/n9841 ), 
        .Q(\IDinst/n9843 ) );
  nnd2s1 \IDinst/U9891  ( .DIN1(\IDinst/RegFile[29][9] ), .DIN2(n1235), 
        .Q(\IDinst/n9842 ) );
  nnd2s1 \IDinst/U9890  ( .DIN1(\IDinst/RegFile[28][9] ), .DIN2(n1241), 
        .Q(\IDinst/n9841 ) );
  nnd2s1 \IDinst/U9889  ( .DIN1(\IDinst/n9839 ), .DIN2(\IDinst/n9838 ), 
        .Q(\IDinst/n9840 ) );
  nnd2s1 \IDinst/U9888  ( .DIN1(\IDinst/n9837 ), .DIN2(n1328), 
        .Q(\IDinst/n9839 ) );
  nnd2s1 \IDinst/U9887  ( .DIN1(\IDinst/n9834 ), .DIN2(n1339), 
        .Q(\IDinst/n9838 ) );
  nnd2s1 \IDinst/U9886  ( .DIN1(\IDinst/n9836 ), .DIN2(\IDinst/n9835 ), 
        .Q(\IDinst/n9837 ) );
  nnd2s1 \IDinst/U9885  ( .DIN1(\IDinst/RegFile[27][9] ), .DIN2(n1235), 
        .Q(\IDinst/n9836 ) );
  nnd2s1 \IDinst/U9884  ( .DIN1(\IDinst/RegFile[26][9] ), .DIN2(n1240), 
        .Q(\IDinst/n9835 ) );
  nnd2s1 \IDinst/U9883  ( .DIN1(\IDinst/n9833 ), .DIN2(\IDinst/n9832 ), 
        .Q(\IDinst/n9834 ) );
  nnd2s1 \IDinst/U9882  ( .DIN1(\IDinst/RegFile[25][9] ), .DIN2(n1235), 
        .Q(\IDinst/n9833 ) );
  nnd2s1 \IDinst/U9881  ( .DIN1(\IDinst/RegFile[24][9] ), .DIN2(n1240), 
        .Q(\IDinst/n9832 ) );
  nnd2s1 \IDinst/U9880  ( .DIN1(\IDinst/n9830 ), .DIN2(\IDinst/n9829 ), 
        .Q(\IDinst/n9831 ) );
  nnd2s1 \IDinst/U9879  ( .DIN1(\IDinst/n9828 ), .DIN2(n1377), 
        .Q(\IDinst/n9830 ) );
  nnd2s1 \IDinst/U9878  ( .DIN1(\IDinst/n9819 ), .DIN2(n1366), 
        .Q(\IDinst/n9829 ) );
  nnd2s1 \IDinst/U9877  ( .DIN1(\IDinst/n9827 ), .DIN2(\IDinst/n9826 ), 
        .Q(\IDinst/n9828 ) );
  nnd2s1 \IDinst/U9876  ( .DIN1(\IDinst/n9825 ), .DIN2(n1328), 
        .Q(\IDinst/n9827 ) );
  nnd2s1 \IDinst/U9875  ( .DIN1(\IDinst/n9822 ), .DIN2(n1339), 
        .Q(\IDinst/n9826 ) );
  nnd2s1 \IDinst/U9874  ( .DIN1(\IDinst/n9824 ), .DIN2(\IDinst/n9823 ), 
        .Q(\IDinst/n9825 ) );
  nnd2s1 \IDinst/U9873  ( .DIN1(\IDinst/RegFile[23][9] ), .DIN2(n1235), 
        .Q(\IDinst/n9824 ) );
  nnd2s1 \IDinst/U9872  ( .DIN1(\IDinst/RegFile[22][9] ), .DIN2(n1240), 
        .Q(\IDinst/n9823 ) );
  nnd2s1 \IDinst/U9871  ( .DIN1(\IDinst/n9821 ), .DIN2(\IDinst/n9820 ), 
        .Q(\IDinst/n9822 ) );
  nnd2s1 \IDinst/U9870  ( .DIN1(\IDinst/RegFile[21][9] ), .DIN2(n1236), 
        .Q(\IDinst/n9821 ) );
  nnd2s1 \IDinst/U9869  ( .DIN1(\IDinst/RegFile[20][9] ), .DIN2(n1240), 
        .Q(\IDinst/n9820 ) );
  nnd2s1 \IDinst/U9868  ( .DIN1(\IDinst/n9818 ), .DIN2(\IDinst/n9817 ), 
        .Q(\IDinst/n9819 ) );
  nnd2s1 \IDinst/U9867  ( .DIN1(\IDinst/n9816 ), .DIN2(n1328), 
        .Q(\IDinst/n9818 ) );
  nnd2s1 \IDinst/U9866  ( .DIN1(\IDinst/n9813 ), .DIN2(n1339), 
        .Q(\IDinst/n9817 ) );
  nnd2s1 \IDinst/U9865  ( .DIN1(\IDinst/n9815 ), .DIN2(\IDinst/n9814 ), 
        .Q(\IDinst/n9816 ) );
  nnd2s1 \IDinst/U9864  ( .DIN1(\IDinst/RegFile[19][9] ), .DIN2(n1236), 
        .Q(\IDinst/n9815 ) );
  nnd2s1 \IDinst/U9863  ( .DIN1(\IDinst/RegFile[18][9] ), .DIN2(n1240), 
        .Q(\IDinst/n9814 ) );
  nnd2s1 \IDinst/U9862  ( .DIN1(\IDinst/n9812 ), .DIN2(\IDinst/n9811 ), 
        .Q(\IDinst/n9813 ) );
  nnd2s1 \IDinst/U9861  ( .DIN1(\IDinst/RegFile[17][9] ), .DIN2(n1236), 
        .Q(\IDinst/n9812 ) );
  nnd2s1 \IDinst/U9860  ( .DIN1(\IDinst/RegFile[16][9] ), .DIN2(n1241), 
        .Q(\IDinst/n9811 ) );
  nnd2s1 \IDinst/U9859  ( .DIN1(\IDinst/n9809 ), .DIN2(\IDinst/n9808 ), 
        .Q(\IDinst/n9810 ) );
  nnd2s1 \IDinst/U9858  ( .DIN1(\IDinst/n9807 ), .DIN2(n665), 
        .Q(\IDinst/n9809 ) );
  nnd2s1 \IDinst/U9857  ( .DIN1(\IDinst/n9786 ), .DIN2(n682), 
        .Q(\IDinst/n9808 ) );
  nnd2s1 \IDinst/U9856  ( .DIN1(\IDinst/n9806 ), .DIN2(\IDinst/n9805 ), 
        .Q(\IDinst/n9807 ) );
  nnd2s1 \IDinst/U9855  ( .DIN1(\IDinst/n9804 ), .DIN2(n1378), 
        .Q(\IDinst/n9806 ) );
  nnd2s1 \IDinst/U9854  ( .DIN1(\IDinst/n9795 ), .DIN2(n1366), 
        .Q(\IDinst/n9805 ) );
  nnd2s1 \IDinst/U9853  ( .DIN1(\IDinst/n9803 ), .DIN2(\IDinst/n9802 ), 
        .Q(\IDinst/n9804 ) );
  nnd2s1 \IDinst/U9852  ( .DIN1(\IDinst/n9801 ), .DIN2(n1328), 
        .Q(\IDinst/n9803 ) );
  nnd2s1 \IDinst/U9851  ( .DIN1(\IDinst/n9798 ), .DIN2(n1340), 
        .Q(\IDinst/n9802 ) );
  nnd2s1 \IDinst/U9850  ( .DIN1(\IDinst/n9800 ), .DIN2(\IDinst/n9799 ), 
        .Q(\IDinst/n9801 ) );
  nnd2s1 \IDinst/U9849  ( .DIN1(\IDinst/RegFile[15][9] ), .DIN2(n1236), 
        .Q(\IDinst/n9800 ) );
  nnd2s1 \IDinst/U9848  ( .DIN1(\IDinst/RegFile[14][9] ), .DIN2(n1240), 
        .Q(\IDinst/n9799 ) );
  nnd2s1 \IDinst/U9847  ( .DIN1(\IDinst/n9797 ), .DIN2(\IDinst/n9796 ), 
        .Q(\IDinst/n9798 ) );
  nnd2s1 \IDinst/U9846  ( .DIN1(\IDinst/RegFile[13][9] ), .DIN2(n1236), 
        .Q(\IDinst/n9797 ) );
  nnd2s1 \IDinst/U9845  ( .DIN1(\IDinst/RegFile[12][9] ), .DIN2(n1240), 
        .Q(\IDinst/n9796 ) );
  nnd2s1 \IDinst/U9844  ( .DIN1(\IDinst/n9794 ), .DIN2(\IDinst/n9793 ), 
        .Q(\IDinst/n9795 ) );
  nnd2s1 \IDinst/U9843  ( .DIN1(\IDinst/n9792 ), .DIN2(n1328), 
        .Q(\IDinst/n9794 ) );
  nnd2s1 \IDinst/U9842  ( .DIN1(\IDinst/n9789 ), .DIN2(n1340), 
        .Q(\IDinst/n9793 ) );
  nnd2s1 \IDinst/U9841  ( .DIN1(\IDinst/n9791 ), .DIN2(\IDinst/n9790 ), 
        .Q(\IDinst/n9792 ) );
  nnd2s1 \IDinst/U9840  ( .DIN1(\IDinst/RegFile[11][9] ), .DIN2(n1236), 
        .Q(\IDinst/n9791 ) );
  nnd2s1 \IDinst/U9839  ( .DIN1(\IDinst/RegFile[10][9] ), .DIN2(n1240), 
        .Q(\IDinst/n9790 ) );
  nnd2s1 \IDinst/U9838  ( .DIN1(\IDinst/n9788 ), .DIN2(\IDinst/n9787 ), 
        .Q(\IDinst/n9789 ) );
  nnd2s1 \IDinst/U9837  ( .DIN1(\IDinst/RegFile[9][9] ), .DIN2(n1236), 
        .Q(\IDinst/n9788 ) );
  nnd2s1 \IDinst/U9836  ( .DIN1(\IDinst/RegFile[8][9] ), .DIN2(n1240), 
        .Q(\IDinst/n9787 ) );
  nnd2s1 \IDinst/U9835  ( .DIN1(\IDinst/n9785 ), .DIN2(\IDinst/n9784 ), 
        .Q(\IDinst/n9786 ) );
  nnd2s1 \IDinst/U9834  ( .DIN1(\IDinst/n9783 ), .DIN2(n1378), 
        .Q(\IDinst/n9785 ) );
  nnd2s1 \IDinst/U9833  ( .DIN1(\IDinst/n9774 ), .DIN2(n1366), 
        .Q(\IDinst/n9784 ) );
  nnd2s1 \IDinst/U9832  ( .DIN1(\IDinst/n9782 ), .DIN2(\IDinst/n9781 ), 
        .Q(\IDinst/n9783 ) );
  nnd2s1 \IDinst/U9831  ( .DIN1(\IDinst/n9780 ), .DIN2(n1328), 
        .Q(\IDinst/n9782 ) );
  nnd2s1 \IDinst/U9830  ( .DIN1(\IDinst/n9777 ), .DIN2(n1340), 
        .Q(\IDinst/n9781 ) );
  nnd2s1 \IDinst/U9829  ( .DIN1(\IDinst/n9779 ), .DIN2(\IDinst/n9778 ), 
        .Q(\IDinst/n9780 ) );
  nnd2s1 \IDinst/U9828  ( .DIN1(\IDinst/RegFile[7][9] ), .DIN2(n1236), 
        .Q(\IDinst/n9779 ) );
  nnd2s1 \IDinst/U9827  ( .DIN1(\IDinst/RegFile[6][9] ), .DIN2(n1239), 
        .Q(\IDinst/n9778 ) );
  nnd2s1 \IDinst/U9826  ( .DIN1(\IDinst/n9776 ), .DIN2(\IDinst/n9775 ), 
        .Q(\IDinst/n9777 ) );
  nnd2s1 \IDinst/U9825  ( .DIN1(\IDinst/RegFile[5][9] ), .DIN2(n1236), 
        .Q(\IDinst/n9776 ) );
  nnd2s1 \IDinst/U9824  ( .DIN1(\IDinst/RegFile[4][9] ), .DIN2(n1239), 
        .Q(\IDinst/n9775 ) );
  nnd2s1 \IDinst/U9823  ( .DIN1(\IDinst/n9773 ), .DIN2(\IDinst/n9772 ), 
        .Q(\IDinst/n9774 ) );
  nnd2s1 \IDinst/U9822  ( .DIN1(\IDinst/n9771 ), .DIN2(n1327), 
        .Q(\IDinst/n9773 ) );
  nnd2s1 \IDinst/U9821  ( .DIN1(\IDinst/n9768 ), .DIN2(n1340), 
        .Q(\IDinst/n9772 ) );
  nnd2s1 \IDinst/U9820  ( .DIN1(\IDinst/n9770 ), .DIN2(\IDinst/n9769 ), 
        .Q(\IDinst/n9771 ) );
  nnd2s1 \IDinst/U9819  ( .DIN1(\IDinst/RegFile[3][9] ), .DIN2(n1236), 
        .Q(\IDinst/n9770 ) );
  nnd2s1 \IDinst/U9818  ( .DIN1(\IDinst/RegFile[2][9] ), .DIN2(n1239), 
        .Q(\IDinst/n9769 ) );
  nnd2s1 \IDinst/U9817  ( .DIN1(\IDinst/n9767 ), .DIN2(\IDinst/n9766 ), 
        .Q(\IDinst/n9768 ) );
  nnd2s1 \IDinst/U9816  ( .DIN1(\IDinst/RegFile[1][9] ), .DIN2(n1236), 
        .Q(\IDinst/n9767 ) );
  nnd2s1 \IDinst/U9815  ( .DIN1(\IDinst/RegFile[0][9] ), .DIN2(n1239), 
        .Q(\IDinst/n9766 ) );
  nnd2s1 \IDinst/U9814  ( .DIN1(\IDinst/n9765 ), .DIN2(n534), 
        .Q(\IDinst/n8908 ) );
  nnd2s1 \IDinst/U9813  ( .DIN1(\IDinst/n9720 ), .DIN2(n634), 
        .Q(\IDinst/n8909 ) );
  nnd2s1 \IDinst/U9812  ( .DIN1(\IDinst/n9764 ), .DIN2(\IDinst/n9763 ), 
        .Q(\IDinst/n9765 ) );
  nnd2s1 \IDinst/U9811  ( .DIN1(\IDinst/n9762 ), .DIN2(n668), 
        .Q(\IDinst/n9764 ) );
  nnd2s1 \IDinst/U9810  ( .DIN1(\IDinst/n9741 ), .DIN2(n680), 
        .Q(\IDinst/n9763 ) );
  nnd2s1 \IDinst/U9809  ( .DIN1(\IDinst/n9761 ), .DIN2(\IDinst/n9760 ), 
        .Q(\IDinst/n9762 ) );
  nnd2s1 \IDinst/U9808  ( .DIN1(\IDinst/n9759 ), .DIN2(n1378), 
        .Q(\IDinst/n9761 ) );
  nnd2s1 \IDinst/U9807  ( .DIN1(\IDinst/n9750 ), .DIN2(n1366), 
        .Q(\IDinst/n9760 ) );
  nnd2s1 \IDinst/U9806  ( .DIN1(\IDinst/n9758 ), .DIN2(\IDinst/n9757 ), 
        .Q(\IDinst/n9759 ) );
  nnd2s1 \IDinst/U9805  ( .DIN1(\IDinst/n9756 ), .DIN2(n1327), 
        .Q(\IDinst/n9758 ) );
  nnd2s1 \IDinst/U9804  ( .DIN1(\IDinst/n9753 ), .DIN2(n1340), 
        .Q(\IDinst/n9757 ) );
  nnd2s1 \IDinst/U9803  ( .DIN1(\IDinst/n9755 ), .DIN2(\IDinst/n9754 ), 
        .Q(\IDinst/n9756 ) );
  nnd2s1 \IDinst/U9802  ( .DIN1(\IDinst/RegFile[31][8] ), .DIN2(n1236), 
        .Q(\IDinst/n9755 ) );
  nnd2s1 \IDinst/U9801  ( .DIN1(\IDinst/RegFile[30][8] ), .DIN2(n1239), 
        .Q(\IDinst/n9754 ) );
  nnd2s1 \IDinst/U9800  ( .DIN1(\IDinst/n9752 ), .DIN2(\IDinst/n9751 ), 
        .Q(\IDinst/n9753 ) );
  nnd2s1 \IDinst/U9799  ( .DIN1(\IDinst/RegFile[29][8] ), .DIN2(n1236), 
        .Q(\IDinst/n9752 ) );
  nnd2s1 \IDinst/U9798  ( .DIN1(\IDinst/RegFile[28][8] ), .DIN2(n1239), 
        .Q(\IDinst/n9751 ) );
  nnd2s1 \IDinst/U9797  ( .DIN1(\IDinst/n9749 ), .DIN2(\IDinst/n9748 ), 
        .Q(\IDinst/n9750 ) );
  nnd2s1 \IDinst/U9796  ( .DIN1(\IDinst/n9747 ), .DIN2(n1327), 
        .Q(\IDinst/n9749 ) );
  nnd2s1 \IDinst/U9795  ( .DIN1(\IDinst/n9744 ), .DIN2(n1340), 
        .Q(\IDinst/n9748 ) );
  nnd2s1 \IDinst/U9794  ( .DIN1(\IDinst/n9746 ), .DIN2(\IDinst/n9745 ), 
        .Q(\IDinst/n9747 ) );
  nnd2s1 \IDinst/U9793  ( .DIN1(\IDinst/RegFile[27][8] ), .DIN2(n1237), 
        .Q(\IDinst/n9746 ) );
  nnd2s1 \IDinst/U9792  ( .DIN1(\IDinst/RegFile[26][8] ), .DIN2(n1239), 
        .Q(\IDinst/n9745 ) );
  nnd2s1 \IDinst/U9791  ( .DIN1(\IDinst/n9743 ), .DIN2(\IDinst/n9742 ), 
        .Q(\IDinst/n9744 ) );
  nnd2s1 \IDinst/U9790  ( .DIN1(\IDinst/RegFile[25][8] ), .DIN2(n1237), 
        .Q(\IDinst/n9743 ) );
  nnd2s1 \IDinst/U9789  ( .DIN1(\IDinst/RegFile[24][8] ), .DIN2(n1239), 
        .Q(\IDinst/n9742 ) );
  nnd2s1 \IDinst/U9788  ( .DIN1(\IDinst/n9740 ), .DIN2(\IDinst/n9739 ), 
        .Q(\IDinst/n9741 ) );
  nnd2s1 \IDinst/U9787  ( .DIN1(\IDinst/n9738 ), .DIN2(n1378), 
        .Q(\IDinst/n9740 ) );
  nnd2s1 \IDinst/U9786  ( .DIN1(\IDinst/n9729 ), .DIN2(n1366), 
        .Q(\IDinst/n9739 ) );
  nnd2s1 \IDinst/U9785  ( .DIN1(\IDinst/n9737 ), .DIN2(\IDinst/n9736 ), 
        .Q(\IDinst/n9738 ) );
  nnd2s1 \IDinst/U9784  ( .DIN1(\IDinst/n9735 ), .DIN2(n1327), 
        .Q(\IDinst/n9737 ) );
  nnd2s1 \IDinst/U9783  ( .DIN1(\IDinst/n9732 ), .DIN2(n1340), 
        .Q(\IDinst/n9736 ) );
  nnd2s1 \IDinst/U9782  ( .DIN1(\IDinst/n9734 ), .DIN2(\IDinst/n9733 ), 
        .Q(\IDinst/n9735 ) );
  nnd2s1 \IDinst/U9781  ( .DIN1(\IDinst/RegFile[23][8] ), .DIN2(n1237), 
        .Q(\IDinst/n9734 ) );
  nnd2s1 \IDinst/U9780  ( .DIN1(\IDinst/RegFile[22][8] ), .DIN2(n1246), 
        .Q(\IDinst/n9733 ) );
  nnd2s1 \IDinst/U9779  ( .DIN1(\IDinst/n9731 ), .DIN2(\IDinst/n9730 ), 
        .Q(\IDinst/n9732 ) );
  nnd2s1 \IDinst/U9778  ( .DIN1(\IDinst/RegFile[21][8] ), .DIN2(n1237), 
        .Q(\IDinst/n9731 ) );
  nnd2s1 \IDinst/U9777  ( .DIN1(\IDinst/RegFile[20][8] ), .DIN2(n1269), 
        .Q(\IDinst/n9730 ) );
  nnd2s1 \IDinst/U9776  ( .DIN1(\IDinst/n9728 ), .DIN2(\IDinst/n9727 ), 
        .Q(\IDinst/n9729 ) );
  nnd2s1 \IDinst/U9775  ( .DIN1(\IDinst/n9726 ), .DIN2(n1327), 
        .Q(\IDinst/n9728 ) );
  nnd2s1 \IDinst/U9774  ( .DIN1(\IDinst/n9723 ), .DIN2(n1340), 
        .Q(\IDinst/n9727 ) );
  nnd2s1 \IDinst/U9773  ( .DIN1(\IDinst/n9725 ), .DIN2(\IDinst/n9724 ), 
        .Q(\IDinst/n9726 ) );
  nnd2s1 \IDinst/U9772  ( .DIN1(\IDinst/RegFile[19][8] ), .DIN2(n1237), 
        .Q(\IDinst/n9725 ) );
  nnd2s1 \IDinst/U9771  ( .DIN1(\IDinst/RegFile[18][8] ), .DIN2(n1269), 
        .Q(\IDinst/n9724 ) );
  nnd2s1 \IDinst/U9770  ( .DIN1(\IDinst/n9722 ), .DIN2(\IDinst/n9721 ), 
        .Q(\IDinst/n9723 ) );
  nnd2s1 \IDinst/U9769  ( .DIN1(\IDinst/RegFile[17][8] ), .DIN2(n1237), 
        .Q(\IDinst/n9722 ) );
  nnd2s1 \IDinst/U9768  ( .DIN1(\IDinst/RegFile[16][8] ), .DIN2(n1269), 
        .Q(\IDinst/n9721 ) );
  nnd2s1 \IDinst/U9767  ( .DIN1(\IDinst/n9719 ), .DIN2(\IDinst/n9718 ), 
        .Q(\IDinst/n9720 ) );
  nnd2s1 \IDinst/U9766  ( .DIN1(\IDinst/n9717 ), .DIN2(n666), 
        .Q(\IDinst/n9719 ) );
  nnd2s1 \IDinst/U9765  ( .DIN1(\IDinst/n9696 ), .DIN2(n681), 
        .Q(\IDinst/n9718 ) );
  nnd2s1 \IDinst/U9764  ( .DIN1(\IDinst/n9716 ), .DIN2(\IDinst/n9715 ), 
        .Q(\IDinst/n9717 ) );
  nnd2s1 \IDinst/U9763  ( .DIN1(\IDinst/n9714 ), .DIN2(n1378), 
        .Q(\IDinst/n9716 ) );
  nnd2s1 \IDinst/U9762  ( .DIN1(\IDinst/n9705 ), .DIN2(n1366), 
        .Q(\IDinst/n9715 ) );
  nnd2s1 \IDinst/U9761  ( .DIN1(\IDinst/n9713 ), .DIN2(\IDinst/n9712 ), 
        .Q(\IDinst/n9714 ) );
  nnd2s1 \IDinst/U9760  ( .DIN1(\IDinst/n9711 ), .DIN2(n1327), 
        .Q(\IDinst/n9713 ) );
  nnd2s1 \IDinst/U9759  ( .DIN1(\IDinst/n9708 ), .DIN2(n1341), 
        .Q(\IDinst/n9712 ) );
  nnd2s1 \IDinst/U9758  ( .DIN1(\IDinst/n9710 ), .DIN2(\IDinst/n9709 ), 
        .Q(\IDinst/n9711 ) );
  nnd2s1 \IDinst/U9757  ( .DIN1(\IDinst/RegFile[15][8] ), .DIN2(n1237), 
        .Q(\IDinst/n9710 ) );
  nnd2s1 \IDinst/U9756  ( .DIN1(\IDinst/RegFile[14][8] ), .DIN2(n1269), 
        .Q(\IDinst/n9709 ) );
  nnd2s1 \IDinst/U9755  ( .DIN1(\IDinst/n9707 ), .DIN2(\IDinst/n9706 ), 
        .Q(\IDinst/n9708 ) );
  nnd2s1 \IDinst/U9754  ( .DIN1(\IDinst/RegFile[13][8] ), .DIN2(n1237), 
        .Q(\IDinst/n9707 ) );
  nnd2s1 \IDinst/U9753  ( .DIN1(\IDinst/RegFile[12][8] ), .DIN2(n1269), 
        .Q(\IDinst/n9706 ) );
  nnd2s1 \IDinst/U9752  ( .DIN1(\IDinst/n9704 ), .DIN2(\IDinst/n9703 ), 
        .Q(\IDinst/n9705 ) );
  nnd2s1 \IDinst/U9751  ( .DIN1(\IDinst/n9702 ), .DIN2(n1327), 
        .Q(\IDinst/n9704 ) );
  nnd2s1 \IDinst/U9750  ( .DIN1(\IDinst/n9699 ), .DIN2(n1341), 
        .Q(\IDinst/n9703 ) );
  nnd2s1 \IDinst/U9749  ( .DIN1(\IDinst/n9701 ), .DIN2(\IDinst/n9700 ), 
        .Q(\IDinst/n9702 ) );
  nnd2s1 \IDinst/U9748  ( .DIN1(\IDinst/RegFile[11][8] ), .DIN2(n1237), 
        .Q(\IDinst/n9701 ) );
  nnd2s1 \IDinst/U9747  ( .DIN1(\IDinst/RegFile[10][8] ), .DIN2(n1268), 
        .Q(\IDinst/n9700 ) );
  nnd2s1 \IDinst/U9746  ( .DIN1(\IDinst/n9698 ), .DIN2(\IDinst/n9697 ), 
        .Q(\IDinst/n9699 ) );
  nnd2s1 \IDinst/U9745  ( .DIN1(\IDinst/RegFile[9][8] ), .DIN2(n1237), 
        .Q(\IDinst/n9698 ) );
  nnd2s1 \IDinst/U9744  ( .DIN1(\IDinst/RegFile[8][8] ), .DIN2(n1268), 
        .Q(\IDinst/n9697 ) );
  nnd2s1 \IDinst/U9743  ( .DIN1(\IDinst/n9695 ), .DIN2(\IDinst/n9694 ), 
        .Q(\IDinst/n9696 ) );
  nnd2s1 \IDinst/U9742  ( .DIN1(\IDinst/n9693 ), .DIN2(n1378), 
        .Q(\IDinst/n9695 ) );
  nnd2s1 \IDinst/U9741  ( .DIN1(\IDinst/n9684 ), .DIN2(n1366), 
        .Q(\IDinst/n9694 ) );
  nnd2s1 \IDinst/U9740  ( .DIN1(\IDinst/n9692 ), .DIN2(\IDinst/n9691 ), 
        .Q(\IDinst/n9693 ) );
  nnd2s1 \IDinst/U9739  ( .DIN1(\IDinst/n9690 ), .DIN2(n1327), 
        .Q(\IDinst/n9692 ) );
  nnd2s1 \IDinst/U9738  ( .DIN1(\IDinst/n9687 ), .DIN2(n1341), 
        .Q(\IDinst/n9691 ) );
  nnd2s1 \IDinst/U9737  ( .DIN1(\IDinst/n9689 ), .DIN2(\IDinst/n9688 ), 
        .Q(\IDinst/n9690 ) );
  nnd2s1 \IDinst/U9736  ( .DIN1(\IDinst/RegFile[7][8] ), .DIN2(n1237), 
        .Q(\IDinst/n9689 ) );
  nnd2s1 \IDinst/U9735  ( .DIN1(\IDinst/RegFile[6][8] ), .DIN2(n1268), 
        .Q(\IDinst/n9688 ) );
  nnd2s1 \IDinst/U9734  ( .DIN1(\IDinst/n9686 ), .DIN2(\IDinst/n9685 ), 
        .Q(\IDinst/n9687 ) );
  nnd2s1 \IDinst/U9733  ( .DIN1(\IDinst/RegFile[5][8] ), .DIN2(n1237), 
        .Q(\IDinst/n9686 ) );
  nnd2s1 \IDinst/U9732  ( .DIN1(\IDinst/RegFile[4][8] ), .DIN2(n1268), 
        .Q(\IDinst/n9685 ) );
  nnd2s1 \IDinst/U9731  ( .DIN1(\IDinst/n9683 ), .DIN2(\IDinst/n9682 ), 
        .Q(\IDinst/n9684 ) );
  nnd2s1 \IDinst/U9730  ( .DIN1(\IDinst/n9681 ), .DIN2(n1327), 
        .Q(\IDinst/n9683 ) );
  nnd2s1 \IDinst/U9729  ( .DIN1(\IDinst/n9678 ), .DIN2(n1341), 
        .Q(\IDinst/n9682 ) );
  nnd2s1 \IDinst/U9728  ( .DIN1(\IDinst/n9680 ), .DIN2(\IDinst/n9679 ), 
        .Q(\IDinst/n9681 ) );
  nnd2s1 \IDinst/U9727  ( .DIN1(\IDinst/RegFile[3][8] ), .DIN2(n1237), 
        .Q(\IDinst/n9680 ) );
  nnd2s1 \IDinst/U9726  ( .DIN1(\IDinst/RegFile[2][8] ), .DIN2(n1268), 
        .Q(\IDinst/n9679 ) );
  nnd2s1 \IDinst/U9725  ( .DIN1(\IDinst/n9677 ), .DIN2(\IDinst/n9676 ), 
        .Q(\IDinst/n9678 ) );
  nnd2s1 \IDinst/U9724  ( .DIN1(\IDinst/RegFile[1][8] ), .DIN2(n1223), 
        .Q(\IDinst/n9677 ) );
  nnd2s1 \IDinst/U9723  ( .DIN1(\IDinst/RegFile[0][8] ), .DIN2(n1268), 
        .Q(\IDinst/n9676 ) );
  nnd2s1 \IDinst/U9722  ( .DIN1(\IDinst/n9675 ), .DIN2(\IDinst/N48 ), 
        .Q(\IDinst/n8906 ) );
  nnd2s1 \IDinst/U9721  ( .DIN1(\IDinst/n9630 ), .DIN2(n533), 
        .Q(\IDinst/n8907 ) );
  nnd2s1 \IDinst/U9720  ( .DIN1(\IDinst/n9674 ), .DIN2(\IDinst/n9673 ), 
        .Q(\IDinst/n9675 ) );
  nnd2s1 \IDinst/U9719  ( .DIN1(\IDinst/n9672 ), .DIN2(n667), 
        .Q(\IDinst/n9674 ) );
  nnd2s1 \IDinst/U9718  ( .DIN1(\IDinst/n9651 ), .DIN2(n683), 
        .Q(\IDinst/n9673 ) );
  nnd2s1 \IDinst/U9717  ( .DIN1(\IDinst/n9671 ), .DIN2(\IDinst/n9670 ), 
        .Q(\IDinst/n9672 ) );
  nnd2s1 \IDinst/U9716  ( .DIN1(\IDinst/n9669 ), .DIN2(n1378), 
        .Q(\IDinst/n9671 ) );
  nnd2s1 \IDinst/U9715  ( .DIN1(\IDinst/n9660 ), .DIN2(n1366), 
        .Q(\IDinst/n9670 ) );
  nnd2s1 \IDinst/U9714  ( .DIN1(\IDinst/n9668 ), .DIN2(\IDinst/n9667 ), 
        .Q(\IDinst/n9669 ) );
  nnd2s1 \IDinst/U9713  ( .DIN1(\IDinst/n9666 ), .DIN2(n1327), 
        .Q(\IDinst/n9668 ) );
  nnd2s1 \IDinst/U9712  ( .DIN1(\IDinst/n9663 ), .DIN2(n1341), 
        .Q(\IDinst/n9667 ) );
  nnd2s1 \IDinst/U9711  ( .DIN1(\IDinst/n9665 ), .DIN2(\IDinst/n9664 ), 
        .Q(\IDinst/n9666 ) );
  nnd2s1 \IDinst/U9710  ( .DIN1(\IDinst/RegFile[31][7] ), .DIN2(n1218), 
        .Q(\IDinst/n9665 ) );
  nnd2s1 \IDinst/U9709  ( .DIN1(\IDinst/RegFile[30][7] ), .DIN2(n1268), 
        .Q(\IDinst/n9664 ) );
  nnd2s1 \IDinst/U9708  ( .DIN1(\IDinst/n9662 ), .DIN2(\IDinst/n9661 ), 
        .Q(\IDinst/n9663 ) );
  nnd2s1 \IDinst/U9707  ( .DIN1(\IDinst/RegFile[29][7] ), .DIN2(n1218), 
        .Q(\IDinst/n9662 ) );
  nnd2s1 \IDinst/U9706  ( .DIN1(\IDinst/RegFile[28][7] ), .DIN2(n1268), 
        .Q(\IDinst/n9661 ) );
  nnd2s1 \IDinst/U9705  ( .DIN1(\IDinst/n9659 ), .DIN2(\IDinst/n9658 ), 
        .Q(\IDinst/n9660 ) );
  nnd2s1 \IDinst/U9704  ( .DIN1(\IDinst/n9657 ), .DIN2(n1327), 
        .Q(\IDinst/n9659 ) );
  nnd2s1 \IDinst/U9703  ( .DIN1(\IDinst/n9654 ), .DIN2(n1341), 
        .Q(\IDinst/n9658 ) );
  nnd2s1 \IDinst/U9702  ( .DIN1(\IDinst/n9656 ), .DIN2(\IDinst/n9655 ), 
        .Q(\IDinst/n9657 ) );
  nnd2s1 \IDinst/U9701  ( .DIN1(\IDinst/RegFile[27][7] ), .DIN2(n1218), 
        .Q(\IDinst/n9656 ) );
  nnd2s1 \IDinst/U9700  ( .DIN1(\IDinst/RegFile[26][7] ), .DIN2(n1268), 
        .Q(\IDinst/n9655 ) );
  nnd2s1 \IDinst/U9699  ( .DIN1(\IDinst/n9653 ), .DIN2(\IDinst/n9652 ), 
        .Q(\IDinst/n9654 ) );
  nnd2s1 \IDinst/U9698  ( .DIN1(\IDinst/RegFile[25][7] ), .DIN2(n1218), 
        .Q(\IDinst/n9653 ) );
  nnd2s1 \IDinst/U9697  ( .DIN1(\IDinst/RegFile[24][7] ), .DIN2(n1267), 
        .Q(\IDinst/n9652 ) );
  nnd2s1 \IDinst/U9696  ( .DIN1(\IDinst/n9650 ), .DIN2(\IDinst/n9649 ), 
        .Q(\IDinst/n9651 ) );
  nnd2s1 \IDinst/U9695  ( .DIN1(\IDinst/n9648 ), .DIN2(n1378), 
        .Q(\IDinst/n9650 ) );
  nnd2s1 \IDinst/U9694  ( .DIN1(\IDinst/n9639 ), .DIN2(n1366), 
        .Q(\IDinst/n9649 ) );
  nnd2s1 \IDinst/U9693  ( .DIN1(\IDinst/n9647 ), .DIN2(\IDinst/n9646 ), 
        .Q(\IDinst/n9648 ) );
  nnd2s1 \IDinst/U9692  ( .DIN1(\IDinst/n9645 ), .DIN2(n1327), 
        .Q(\IDinst/n9647 ) );
  nnd2s1 \IDinst/U9691  ( .DIN1(\IDinst/n9642 ), .DIN2(n1341), 
        .Q(\IDinst/n9646 ) );
  nnd2s1 \IDinst/U9690  ( .DIN1(\IDinst/n9644 ), .DIN2(\IDinst/n9643 ), 
        .Q(\IDinst/n9645 ) );
  nnd2s1 \IDinst/U9689  ( .DIN1(\IDinst/RegFile[23][7] ), .DIN2(n1218), 
        .Q(\IDinst/n9644 ) );
  nnd2s1 \IDinst/U9688  ( .DIN1(\IDinst/RegFile[22][7] ), .DIN2(n1267), 
        .Q(\IDinst/n9643 ) );
  nnd2s1 \IDinst/U9687  ( .DIN1(\IDinst/n9641 ), .DIN2(\IDinst/n9640 ), 
        .Q(\IDinst/n9642 ) );
  nnd2s1 \IDinst/U9686  ( .DIN1(\IDinst/RegFile[21][7] ), .DIN2(n1218), 
        .Q(\IDinst/n9641 ) );
  nnd2s1 \IDinst/U9685  ( .DIN1(\IDinst/RegFile[20][7] ), .DIN2(n1267), 
        .Q(\IDinst/n9640 ) );
  nnd2s1 \IDinst/U9684  ( .DIN1(\IDinst/n9638 ), .DIN2(\IDinst/n9637 ), 
        .Q(\IDinst/n9639 ) );
  nnd2s1 \IDinst/U9683  ( .DIN1(\IDinst/n9636 ), .DIN2(n1326), 
        .Q(\IDinst/n9638 ) );
  nnd2s1 \IDinst/U9682  ( .DIN1(\IDinst/n9633 ), .DIN2(n1341), 
        .Q(\IDinst/n9637 ) );
  nnd2s1 \IDinst/U9681  ( .DIN1(\IDinst/n9635 ), .DIN2(\IDinst/n9634 ), 
        .Q(\IDinst/n9636 ) );
  nnd2s1 \IDinst/U9680  ( .DIN1(\IDinst/RegFile[19][7] ), .DIN2(n1218), 
        .Q(\IDinst/n9635 ) );
  nnd2s1 \IDinst/U9679  ( .DIN1(\IDinst/RegFile[18][7] ), .DIN2(n1267), 
        .Q(\IDinst/n9634 ) );
  nnd2s1 \IDinst/U9678  ( .DIN1(\IDinst/n9632 ), .DIN2(\IDinst/n9631 ), 
        .Q(\IDinst/n9633 ) );
  nnd2s1 \IDinst/U9677  ( .DIN1(\IDinst/RegFile[17][7] ), .DIN2(n1218), 
        .Q(\IDinst/n9632 ) );
  nnd2s1 \IDinst/U9676  ( .DIN1(\IDinst/RegFile[16][7] ), .DIN2(n1267), 
        .Q(\IDinst/n9631 ) );
  nnd2s1 \IDinst/U9675  ( .DIN1(\IDinst/n9629 ), .DIN2(\IDinst/n9628 ), 
        .Q(\IDinst/n9630 ) );
  nnd2s1 \IDinst/U9674  ( .DIN1(\IDinst/n9627 ), .DIN2(n665), 
        .Q(\IDinst/n9629 ) );
  nnd2s1 \IDinst/U9673  ( .DIN1(\IDinst/n9606 ), .DIN2(n682), 
        .Q(\IDinst/n9628 ) );
  nnd2s1 \IDinst/U9672  ( .DIN1(\IDinst/n9626 ), .DIN2(\IDinst/n9625 ), 
        .Q(\IDinst/n9627 ) );
  nnd2s1 \IDinst/U9671  ( .DIN1(\IDinst/n9624 ), .DIN2(n1378), 
        .Q(\IDinst/n9626 ) );
  nnd2s1 \IDinst/U9670  ( .DIN1(\IDinst/n9615 ), .DIN2(n1370), 
        .Q(\IDinst/n9625 ) );
  nnd2s1 \IDinst/U9669  ( .DIN1(\IDinst/n9623 ), .DIN2(\IDinst/n9622 ), 
        .Q(\IDinst/n9624 ) );
  nnd2s1 \IDinst/U9668  ( .DIN1(\IDinst/n9621 ), .DIN2(n1326), 
        .Q(\IDinst/n9623 ) );
  nnd2s1 \IDinst/U9667  ( .DIN1(\IDinst/n9618 ), .DIN2(n1341), 
        .Q(\IDinst/n9622 ) );
  nnd2s1 \IDinst/U9666  ( .DIN1(\IDinst/n9620 ), .DIN2(\IDinst/n9619 ), 
        .Q(\IDinst/n9621 ) );
  nnd2s1 \IDinst/U9665  ( .DIN1(\IDinst/RegFile[15][7] ), .DIN2(n1219), 
        .Q(\IDinst/n9620 ) );
  nnd2s1 \IDinst/U9664  ( .DIN1(\IDinst/RegFile[14][7] ), .DIN2(n1267), 
        .Q(\IDinst/n9619 ) );
  nnd2s1 \IDinst/U9663  ( .DIN1(\IDinst/n9617 ), .DIN2(\IDinst/n9616 ), 
        .Q(\IDinst/n9618 ) );
  nnd2s1 \IDinst/U9662  ( .DIN1(\IDinst/RegFile[13][7] ), .DIN2(n1219), 
        .Q(\IDinst/n9617 ) );
  nnd2s1 \IDinst/U9661  ( .DIN1(\IDinst/RegFile[12][7] ), .DIN2(n1267), 
        .Q(\IDinst/n9616 ) );
  nnd2s1 \IDinst/U9660  ( .DIN1(\IDinst/n9614 ), .DIN2(\IDinst/n9613 ), 
        .Q(\IDinst/n9615 ) );
  nnd2s1 \IDinst/U9659  ( .DIN1(\IDinst/n9612 ), .DIN2(n1326), 
        .Q(\IDinst/n9614 ) );
  nnd2s1 \IDinst/U9658  ( .DIN1(\IDinst/n9609 ), .DIN2(n1342), 
        .Q(\IDinst/n9613 ) );
  nnd2s1 \IDinst/U9657  ( .DIN1(\IDinst/n9611 ), .DIN2(\IDinst/n9610 ), 
        .Q(\IDinst/n9612 ) );
  nnd2s1 \IDinst/U9656  ( .DIN1(\IDinst/RegFile[11][7] ), .DIN2(n1219), 
        .Q(\IDinst/n9611 ) );
  nnd2s1 \IDinst/U9655  ( .DIN1(\IDinst/RegFile[10][7] ), .DIN2(n1267), 
        .Q(\IDinst/n9610 ) );
  nnd2s1 \IDinst/U9654  ( .DIN1(\IDinst/n9608 ), .DIN2(\IDinst/n9607 ), 
        .Q(\IDinst/n9609 ) );
  nnd2s1 \IDinst/U9653  ( .DIN1(\IDinst/RegFile[9][7] ), .DIN2(n1219), 
        .Q(\IDinst/n9608 ) );
  nnd2s1 \IDinst/U9652  ( .DIN1(\IDinst/RegFile[8][7] ), .DIN2(n1267), 
        .Q(\IDinst/n9607 ) );
  nnd2s1 \IDinst/U9651  ( .DIN1(\IDinst/n9605 ), .DIN2(\IDinst/n9604 ), 
        .Q(\IDinst/n9606 ) );
  nnd2s1 \IDinst/U9650  ( .DIN1(\IDinst/n9603 ), .DIN2(n1379), 
        .Q(\IDinst/n9605 ) );
  nnd2s1 \IDinst/U9649  ( .DIN1(\IDinst/n9594 ), .DIN2(n1369), 
        .Q(\IDinst/n9604 ) );
  nnd2s1 \IDinst/U9648  ( .DIN1(\IDinst/n9602 ), .DIN2(\IDinst/n9601 ), 
        .Q(\IDinst/n9603 ) );
  nnd2s1 \IDinst/U9647  ( .DIN1(\IDinst/n9600 ), .DIN2(n1326), 
        .Q(\IDinst/n9602 ) );
  nnd2s1 \IDinst/U9646  ( .DIN1(\IDinst/n9597 ), .DIN2(n1342), 
        .Q(\IDinst/n9601 ) );
  nnd2s1 \IDinst/U9645  ( .DIN1(\IDinst/n9599 ), .DIN2(\IDinst/n9598 ), 
        .Q(\IDinst/n9600 ) );
  nnd2s1 \IDinst/U9644  ( .DIN1(\IDinst/RegFile[7][7] ), .DIN2(n1219), 
        .Q(\IDinst/n9599 ) );
  nnd2s1 \IDinst/U9643  ( .DIN1(\IDinst/RegFile[6][7] ), .DIN2(n1266), 
        .Q(\IDinst/n9598 ) );
  nnd2s1 \IDinst/U9642  ( .DIN1(\IDinst/n9596 ), .DIN2(\IDinst/n9595 ), 
        .Q(\IDinst/n9597 ) );
  nnd2s1 \IDinst/U9641  ( .DIN1(\IDinst/RegFile[5][7] ), .DIN2(n1219), 
        .Q(\IDinst/n9596 ) );
  nnd2s1 \IDinst/U9640  ( .DIN1(\IDinst/RegFile[4][7] ), .DIN2(n1266), 
        .Q(\IDinst/n9595 ) );
  nnd2s1 \IDinst/U9639  ( .DIN1(\IDinst/n9593 ), .DIN2(\IDinst/n9592 ), 
        .Q(\IDinst/n9594 ) );
  nnd2s1 \IDinst/U9638  ( .DIN1(\IDinst/n9591 ), .DIN2(n1326), 
        .Q(\IDinst/n9593 ) );
  nnd2s1 \IDinst/U9637  ( .DIN1(\IDinst/n9588 ), .DIN2(n1342), 
        .Q(\IDinst/n9592 ) );
  nnd2s1 \IDinst/U9636  ( .DIN1(\IDinst/n9590 ), .DIN2(\IDinst/n9589 ), 
        .Q(\IDinst/n9591 ) );
  nnd2s1 \IDinst/U9635  ( .DIN1(\IDinst/RegFile[3][7] ), .DIN2(n1219), 
        .Q(\IDinst/n9590 ) );
  nnd2s1 \IDinst/U9634  ( .DIN1(\IDinst/RegFile[2][7] ), .DIN2(n1266), 
        .Q(\IDinst/n9589 ) );
  nnd2s1 \IDinst/U9633  ( .DIN1(\IDinst/n9587 ), .DIN2(\IDinst/n9586 ), 
        .Q(\IDinst/n9588 ) );
  nnd2s1 \IDinst/U9632  ( .DIN1(\IDinst/RegFile[1][7] ), .DIN2(n1219), 
        .Q(\IDinst/n9587 ) );
  nnd2s1 \IDinst/U9631  ( .DIN1(\IDinst/RegFile[0][7] ), .DIN2(n1266), 
        .Q(\IDinst/n9586 ) );
  nnd2s1 \IDinst/U9630  ( .DIN1(\IDinst/n9585 ), .DIN2(n535), 
        .Q(\IDinst/n8904 ) );
  nnd2s1 \IDinst/U9629  ( .DIN1(\IDinst/n9540 ), .DIN2(n634), 
        .Q(\IDinst/n8905 ) );
  nnd2s1 \IDinst/U9628  ( .DIN1(\IDinst/n9584 ), .DIN2(\IDinst/n9583 ), 
        .Q(\IDinst/n9585 ) );
  nnd2s1 \IDinst/U9627  ( .DIN1(\IDinst/n9582 ), .DIN2(n668), 
        .Q(\IDinst/n9584 ) );
  nnd2s1 \IDinst/U9626  ( .DIN1(\IDinst/n9561 ), .DIN2(n680), 
        .Q(\IDinst/n9583 ) );
  nnd2s1 \IDinst/U9625  ( .DIN1(\IDinst/n9581 ), .DIN2(\IDinst/n9580 ), 
        .Q(\IDinst/n9582 ) );
  nnd2s1 \IDinst/U9624  ( .DIN1(\IDinst/n9579 ), .DIN2(n1379), 
        .Q(\IDinst/n9581 ) );
  nnd2s1 \IDinst/U9623  ( .DIN1(\IDinst/n9570 ), .DIN2(n1368), 
        .Q(\IDinst/n9580 ) );
  nnd2s1 \IDinst/U9622  ( .DIN1(\IDinst/n9578 ), .DIN2(\IDinst/n9577 ), 
        .Q(\IDinst/n9579 ) );
  nnd2s1 \IDinst/U9621  ( .DIN1(\IDinst/n9576 ), .DIN2(n1326), 
        .Q(\IDinst/n9578 ) );
  nnd2s1 \IDinst/U9620  ( .DIN1(\IDinst/n9573 ), .DIN2(n1342), 
        .Q(\IDinst/n9577 ) );
  nnd2s1 \IDinst/U9619  ( .DIN1(\IDinst/n9575 ), .DIN2(\IDinst/n9574 ), 
        .Q(\IDinst/n9576 ) );
  nnd2s1 \IDinst/U9618  ( .DIN1(\IDinst/RegFile[31][6] ), .DIN2(n1219), 
        .Q(\IDinst/n9575 ) );
  nnd2s1 \IDinst/U9617  ( .DIN1(\IDinst/RegFile[30][6] ), .DIN2(n1266), 
        .Q(\IDinst/n9574 ) );
  nnd2s1 \IDinst/U9616  ( .DIN1(\IDinst/n9572 ), .DIN2(\IDinst/n9571 ), 
        .Q(\IDinst/n9573 ) );
  nnd2s1 \IDinst/U9615  ( .DIN1(\IDinst/RegFile[29][6] ), .DIN2(n1219), 
        .Q(\IDinst/n9572 ) );
  nnd2s1 \IDinst/U9614  ( .DIN1(\IDinst/RegFile[28][6] ), .DIN2(n1266), 
        .Q(\IDinst/n9571 ) );
  nnd2s1 \IDinst/U9613  ( .DIN1(\IDinst/n9569 ), .DIN2(\IDinst/n9568 ), 
        .Q(\IDinst/n9570 ) );
  nnd2s1 \IDinst/U9612  ( .DIN1(\IDinst/n9567 ), .DIN2(n1326), 
        .Q(\IDinst/n9569 ) );
  nnd2s1 \IDinst/U9611  ( .DIN1(\IDinst/n9564 ), .DIN2(n1342), 
        .Q(\IDinst/n9568 ) );
  nnd2s1 \IDinst/U9610  ( .DIN1(\IDinst/n9566 ), .DIN2(\IDinst/n9565 ), 
        .Q(\IDinst/n9567 ) );
  nnd2s1 \IDinst/U9609  ( .DIN1(\IDinst/RegFile[27][6] ), .DIN2(n1219), 
        .Q(\IDinst/n9566 ) );
  nnd2s1 \IDinst/U9608  ( .DIN1(\IDinst/RegFile[26][6] ), .DIN2(n1266), 
        .Q(\IDinst/n9565 ) );
  nnd2s1 \IDinst/U9607  ( .DIN1(\IDinst/n9563 ), .DIN2(\IDinst/n9562 ), 
        .Q(\IDinst/n9564 ) );
  nnd2s1 \IDinst/U9606  ( .DIN1(\IDinst/RegFile[25][6] ), .DIN2(n1219), 
        .Q(\IDinst/n9563 ) );
  nnd2s1 \IDinst/U9605  ( .DIN1(\IDinst/RegFile[24][6] ), .DIN2(n1266), 
        .Q(\IDinst/n9562 ) );
  nnd2s1 \IDinst/U9604  ( .DIN1(\IDinst/n9560 ), .DIN2(\IDinst/n9559 ), 
        .Q(\IDinst/n9561 ) );
  nnd2s1 \IDinst/U9603  ( .DIN1(\IDinst/n9558 ), .DIN2(n1379), 
        .Q(\IDinst/n9560 ) );
  nnd2s1 \IDinst/U9602  ( .DIN1(\IDinst/n9549 ), .DIN2(n1367), 
        .Q(\IDinst/n9559 ) );
  nnd2s1 \IDinst/U9601  ( .DIN1(\IDinst/n9557 ), .DIN2(\IDinst/n9556 ), 
        .Q(\IDinst/n9558 ) );
  nnd2s1 \IDinst/U9600  ( .DIN1(\IDinst/n9555 ), .DIN2(n1326), 
        .Q(\IDinst/n9557 ) );
  nnd2s1 \IDinst/U9599  ( .DIN1(\IDinst/n9552 ), .DIN2(n1342), 
        .Q(\IDinst/n9556 ) );
  nnd2s1 \IDinst/U9598  ( .DIN1(\IDinst/n9554 ), .DIN2(\IDinst/n9553 ), 
        .Q(\IDinst/n9555 ) );
  nnd2s1 \IDinst/U9597  ( .DIN1(\IDinst/RegFile[23][6] ), .DIN2(n1219), 
        .Q(\IDinst/n9554 ) );
  nnd2s1 \IDinst/U9596  ( .DIN1(\IDinst/RegFile[22][6] ), .DIN2(n1266), 
        .Q(\IDinst/n9553 ) );
  nnd2s1 \IDinst/U9595  ( .DIN1(\IDinst/n9551 ), .DIN2(\IDinst/n9550 ), 
        .Q(\IDinst/n9552 ) );
  nnd2s1 \IDinst/U9594  ( .DIN1(\IDinst/RegFile[21][6] ), .DIN2(n1220), 
        .Q(\IDinst/n9551 ) );
  nnd2s1 \IDinst/U9593  ( .DIN1(\IDinst/RegFile[20][6] ), .DIN2(n1265), 
        .Q(\IDinst/n9550 ) );
  nnd2s1 \IDinst/U9592  ( .DIN1(\IDinst/n9548 ), .DIN2(\IDinst/n9547 ), 
        .Q(\IDinst/n9549 ) );
  nnd2s1 \IDinst/U9591  ( .DIN1(\IDinst/n9546 ), .DIN2(n1326), 
        .Q(\IDinst/n9548 ) );
  nnd2s1 \IDinst/U9590  ( .DIN1(\IDinst/n9543 ), .DIN2(n1342), 
        .Q(\IDinst/n9547 ) );
  nnd2s1 \IDinst/U9589  ( .DIN1(\IDinst/n9545 ), .DIN2(\IDinst/n9544 ), 
        .Q(\IDinst/n9546 ) );
  nnd2s1 \IDinst/U9588  ( .DIN1(\IDinst/RegFile[19][6] ), .DIN2(n1220), 
        .Q(\IDinst/n9545 ) );
  nnd2s1 \IDinst/U9587  ( .DIN1(\IDinst/RegFile[18][6] ), .DIN2(n1265), 
        .Q(\IDinst/n9544 ) );
  nnd2s1 \IDinst/U9586  ( .DIN1(\IDinst/n9542 ), .DIN2(\IDinst/n9541 ), 
        .Q(\IDinst/n9543 ) );
  nnd2s1 \IDinst/U9585  ( .DIN1(\IDinst/RegFile[17][6] ), .DIN2(n1220), 
        .Q(\IDinst/n9542 ) );
  nnd2s1 \IDinst/U9584  ( .DIN1(\IDinst/RegFile[16][6] ), .DIN2(n1265), 
        .Q(\IDinst/n9541 ) );
  nnd2s1 \IDinst/U9583  ( .DIN1(\IDinst/n9539 ), .DIN2(\IDinst/n9538 ), 
        .Q(\IDinst/n9540 ) );
  nnd2s1 \IDinst/U9582  ( .DIN1(\IDinst/n9537 ), .DIN2(n666), 
        .Q(\IDinst/n9539 ) );
  nnd2s1 \IDinst/U9581  ( .DIN1(\IDinst/n9516 ), .DIN2(n681), 
        .Q(\IDinst/n9538 ) );
  nnd2s1 \IDinst/U9580  ( .DIN1(\IDinst/n9536 ), .DIN2(\IDinst/n9535 ), 
        .Q(\IDinst/n9537 ) );
  nnd2s1 \IDinst/U9579  ( .DIN1(\IDinst/n9534 ), .DIN2(n1379), 
        .Q(\IDinst/n9536 ) );
  nnd2s1 \IDinst/U9578  ( .DIN1(\IDinst/n9525 ), .DIN2(n1366), 
        .Q(\IDinst/n9535 ) );
  nnd2s1 \IDinst/U9577  ( .DIN1(\IDinst/n9533 ), .DIN2(\IDinst/n9532 ), 
        .Q(\IDinst/n9534 ) );
  nnd2s1 \IDinst/U9576  ( .DIN1(\IDinst/n9531 ), .DIN2(n1326), 
        .Q(\IDinst/n9533 ) );
  nnd2s1 \IDinst/U9575  ( .DIN1(\IDinst/n9528 ), .DIN2(n1342), 
        .Q(\IDinst/n9532 ) );
  nnd2s1 \IDinst/U9574  ( .DIN1(\IDinst/n9530 ), .DIN2(\IDinst/n9529 ), 
        .Q(\IDinst/n9531 ) );
  nnd2s1 \IDinst/U9573  ( .DIN1(\IDinst/RegFile[15][6] ), .DIN2(n1220), 
        .Q(\IDinst/n9530 ) );
  nnd2s1 \IDinst/U9572  ( .DIN1(\IDinst/RegFile[14][6] ), .DIN2(n1265), 
        .Q(\IDinst/n9529 ) );
  nnd2s1 \IDinst/U9571  ( .DIN1(\IDinst/n9527 ), .DIN2(\IDinst/n9526 ), 
        .Q(\IDinst/n9528 ) );
  nnd2s1 \IDinst/U9570  ( .DIN1(\IDinst/RegFile[13][6] ), .DIN2(n1220), 
        .Q(\IDinst/n9527 ) );
  nnd2s1 \IDinst/U9569  ( .DIN1(\IDinst/RegFile[12][6] ), .DIN2(n1265), 
        .Q(\IDinst/n9526 ) );
  nnd2s1 \IDinst/U9568  ( .DIN1(\IDinst/n9524 ), .DIN2(\IDinst/n9523 ), 
        .Q(\IDinst/n9525 ) );
  nnd2s1 \IDinst/U9567  ( .DIN1(\IDinst/n9522 ), .DIN2(n1326), 
        .Q(\IDinst/n9524 ) );
  nnd2s1 \IDinst/U9566  ( .DIN1(\IDinst/n9519 ), .DIN2(n1342), 
        .Q(\IDinst/n9523 ) );
  nnd2s1 \IDinst/U9565  ( .DIN1(\IDinst/n9521 ), .DIN2(\IDinst/n9520 ), 
        .Q(\IDinst/n9522 ) );
  nnd2s1 \IDinst/U9564  ( .DIN1(\IDinst/RegFile[11][6] ), .DIN2(n1220), 
        .Q(\IDinst/n9521 ) );
  nnd2s1 \IDinst/U9563  ( .DIN1(\IDinst/RegFile[10][6] ), .DIN2(n1265), 
        .Q(\IDinst/n9520 ) );
  nnd2s1 \IDinst/U9562  ( .DIN1(\IDinst/n9518 ), .DIN2(\IDinst/n9517 ), 
        .Q(\IDinst/n9519 ) );
  nnd2s1 \IDinst/U9561  ( .DIN1(\IDinst/RegFile[9][6] ), .DIN2(n1220), 
        .Q(\IDinst/n9518 ) );
  nnd2s1 \IDinst/U9560  ( .DIN1(\IDinst/RegFile[8][6] ), .DIN2(n1265), 
        .Q(\IDinst/n9517 ) );
  nnd2s1 \IDinst/U9559  ( .DIN1(\IDinst/n9515 ), .DIN2(\IDinst/n9514 ), 
        .Q(\IDinst/n9516 ) );
  nnd2s1 \IDinst/U9558  ( .DIN1(\IDinst/n9513 ), .DIN2(n1379), 
        .Q(\IDinst/n9515 ) );
  nnd2s1 \IDinst/U9557  ( .DIN1(\IDinst/n9504 ), .DIN2(n1365), 
        .Q(\IDinst/n9514 ) );
  nnd2s1 \IDinst/U9556  ( .DIN1(\IDinst/n9512 ), .DIN2(\IDinst/n9511 ), 
        .Q(\IDinst/n9513 ) );
  nnd2s1 \IDinst/U9555  ( .DIN1(\IDinst/n9510 ), .DIN2(n1326), 
        .Q(\IDinst/n9512 ) );
  nnd2s1 \IDinst/U9554  ( .DIN1(\IDinst/n9507 ), .DIN2(n1343), 
        .Q(\IDinst/n9511 ) );
  nnd2s1 \IDinst/U9553  ( .DIN1(\IDinst/n9509 ), .DIN2(\IDinst/n9508 ), 
        .Q(\IDinst/n9510 ) );
  nnd2s1 \IDinst/U9552  ( .DIN1(\IDinst/RegFile[7][6] ), .DIN2(n1220), 
        .Q(\IDinst/n9509 ) );
  nnd2s1 \IDinst/U9551  ( .DIN1(\IDinst/RegFile[6][6] ), .DIN2(n1265), 
        .Q(\IDinst/n9508 ) );
  nnd2s1 \IDinst/U9550  ( .DIN1(\IDinst/n9506 ), .DIN2(\IDinst/n9505 ), 
        .Q(\IDinst/n9507 ) );
  nnd2s1 \IDinst/U9549  ( .DIN1(\IDinst/RegFile[5][6] ), .DIN2(n1220), 
        .Q(\IDinst/n9506 ) );
  nnd2s1 \IDinst/U9548  ( .DIN1(\IDinst/RegFile[4][6] ), .DIN2(n1265), 
        .Q(\IDinst/n9505 ) );
  nnd2s1 \IDinst/U9547  ( .DIN1(\IDinst/n9503 ), .DIN2(\IDinst/n9502 ), 
        .Q(\IDinst/n9504 ) );
  nnd2s1 \IDinst/U9546  ( .DIN1(\IDinst/n9501 ), .DIN2(n1326), 
        .Q(\IDinst/n9503 ) );
  nnd2s1 \IDinst/U9545  ( .DIN1(\IDinst/n9498 ), .DIN2(n1343), 
        .Q(\IDinst/n9502 ) );
  nnd2s1 \IDinst/U9544  ( .DIN1(\IDinst/n9500 ), .DIN2(\IDinst/n9499 ), 
        .Q(\IDinst/n9501 ) );
  nnd2s1 \IDinst/U9543  ( .DIN1(\IDinst/RegFile[3][6] ), .DIN2(n1220), 
        .Q(\IDinst/n9500 ) );
  nnd2s1 \IDinst/U9542  ( .DIN1(\IDinst/RegFile[2][6] ), .DIN2(n1264), 
        .Q(\IDinst/n9499 ) );
  nnd2s1 \IDinst/U9541  ( .DIN1(\IDinst/n9497 ), .DIN2(\IDinst/n9496 ), 
        .Q(\IDinst/n9498 ) );
  nnd2s1 \IDinst/U9540  ( .DIN1(\IDinst/RegFile[1][6] ), .DIN2(n1220), 
        .Q(\IDinst/n9497 ) );
  nnd2s1 \IDinst/U9539  ( .DIN1(\IDinst/RegFile[0][6] ), .DIN2(n1264), 
        .Q(\IDinst/n9496 ) );
  nnd2s1 \IDinst/U9538  ( .DIN1(\IDinst/n9495 ), .DIN2(n534), 
        .Q(\IDinst/n8902 ) );
  nnd2s1 \IDinst/U9537  ( .DIN1(\IDinst/n9450 ), .DIN2(n533), 
        .Q(\IDinst/n8903 ) );
  nnd2s1 \IDinst/U9536  ( .DIN1(\IDinst/n9494 ), .DIN2(\IDinst/n9493 ), 
        .Q(\IDinst/n9495 ) );
  nnd2s1 \IDinst/U9535  ( .DIN1(\IDinst/n9492 ), .DIN2(n667), 
        .Q(\IDinst/n9494 ) );
  nnd2s1 \IDinst/U9534  ( .DIN1(\IDinst/n9471 ), .DIN2(n683), 
        .Q(\IDinst/n9493 ) );
  nnd2s1 \IDinst/U9533  ( .DIN1(\IDinst/n9491 ), .DIN2(\IDinst/n9490 ), 
        .Q(\IDinst/n9492 ) );
  nnd2s1 \IDinst/U9532  ( .DIN1(\IDinst/n9489 ), .DIN2(n1379), 
        .Q(\IDinst/n9491 ) );
  nnd2s1 \IDinst/U9531  ( .DIN1(\IDinst/n9480 ), .DIN2(n1371), 
        .Q(\IDinst/n9490 ) );
  nnd2s1 \IDinst/U9530  ( .DIN1(\IDinst/n9488 ), .DIN2(\IDinst/n9487 ), 
        .Q(\IDinst/n9489 ) );
  nnd2s1 \IDinst/U9529  ( .DIN1(\IDinst/n9486 ), .DIN2(n1325), 
        .Q(\IDinst/n9488 ) );
  nnd2s1 \IDinst/U9528  ( .DIN1(\IDinst/n9483 ), .DIN2(n1343), 
        .Q(\IDinst/n9487 ) );
  nnd2s1 \IDinst/U9527  ( .DIN1(\IDinst/n9485 ), .DIN2(\IDinst/n9484 ), 
        .Q(\IDinst/n9486 ) );
  nnd2s1 \IDinst/U9526  ( .DIN1(\IDinst/RegFile[31][5] ), .DIN2(n1220), 
        .Q(\IDinst/n9485 ) );
  nnd2s1 \IDinst/U9525  ( .DIN1(\IDinst/RegFile[30][5] ), .DIN2(n1264), 
        .Q(\IDinst/n9484 ) );
  nnd2s1 \IDinst/U9524  ( .DIN1(\IDinst/n9482 ), .DIN2(\IDinst/n9481 ), 
        .Q(\IDinst/n9483 ) );
  nnd2s1 \IDinst/U9523  ( .DIN1(\IDinst/RegFile[29][5] ), .DIN2(n1220), 
        .Q(\IDinst/n9482 ) );
  nnd2s1 \IDinst/U9522  ( .DIN1(\IDinst/RegFile[28][5] ), .DIN2(n1264), 
        .Q(\IDinst/n9481 ) );
  nnd2s1 \IDinst/U9521  ( .DIN1(\IDinst/n9479 ), .DIN2(\IDinst/n9478 ), 
        .Q(\IDinst/n9480 ) );
  nnd2s1 \IDinst/U9520  ( .DIN1(\IDinst/n9477 ), .DIN2(n1325), 
        .Q(\IDinst/n9479 ) );
  nnd2s1 \IDinst/U9519  ( .DIN1(\IDinst/n9474 ), .DIN2(n1343), 
        .Q(\IDinst/n9478 ) );
  nnd2s1 \IDinst/U9518  ( .DIN1(\IDinst/n9476 ), .DIN2(\IDinst/n9475 ), 
        .Q(\IDinst/n9477 ) );
  nnd2s1 \IDinst/U9517  ( .DIN1(\IDinst/RegFile[27][5] ), .DIN2(n1221), 
        .Q(\IDinst/n9476 ) );
  nnd2s1 \IDinst/U9516  ( .DIN1(\IDinst/RegFile[26][5] ), .DIN2(n1264), 
        .Q(\IDinst/n9475 ) );
  nnd2s1 \IDinst/U9515  ( .DIN1(\IDinst/n9473 ), .DIN2(\IDinst/n9472 ), 
        .Q(\IDinst/n9474 ) );
  nnd2s1 \IDinst/U9514  ( .DIN1(\IDinst/RegFile[25][5] ), .DIN2(n1221), 
        .Q(\IDinst/n9473 ) );
  nnd2s1 \IDinst/U9513  ( .DIN1(\IDinst/RegFile[24][5] ), .DIN2(n1264), 
        .Q(\IDinst/n9472 ) );
  nnd2s1 \IDinst/U9512  ( .DIN1(\IDinst/n9470 ), .DIN2(\IDinst/n9469 ), 
        .Q(\IDinst/n9471 ) );
  nnd2s1 \IDinst/U9511  ( .DIN1(\IDinst/n9468 ), .DIN2(n1379), 
        .Q(\IDinst/n9470 ) );
  nnd2s1 \IDinst/U9510  ( .DIN1(\IDinst/n9459 ), .DIN2(n1370), 
        .Q(\IDinst/n9469 ) );
  nnd2s1 \IDinst/U9509  ( .DIN1(\IDinst/n9467 ), .DIN2(\IDinst/n9466 ), 
        .Q(\IDinst/n9468 ) );
  nnd2s1 \IDinst/U9508  ( .DIN1(\IDinst/n9465 ), .DIN2(n1325), 
        .Q(\IDinst/n9467 ) );
  nnd2s1 \IDinst/U9507  ( .DIN1(\IDinst/n9462 ), .DIN2(n1343), 
        .Q(\IDinst/n9466 ) );
  nnd2s1 \IDinst/U9506  ( .DIN1(\IDinst/n9464 ), .DIN2(\IDinst/n9463 ), 
        .Q(\IDinst/n9465 ) );
  nnd2s1 \IDinst/U9505  ( .DIN1(\IDinst/RegFile[23][5] ), .DIN2(n1221), 
        .Q(\IDinst/n9464 ) );
  nnd2s1 \IDinst/U9504  ( .DIN1(\IDinst/RegFile[22][5] ), .DIN2(n1264), 
        .Q(\IDinst/n9463 ) );
  nnd2s1 \IDinst/U9503  ( .DIN1(\IDinst/n9461 ), .DIN2(\IDinst/n9460 ), 
        .Q(\IDinst/n9462 ) );
  nnd2s1 \IDinst/U9502  ( .DIN1(\IDinst/RegFile[21][5] ), .DIN2(n1221), 
        .Q(\IDinst/n9461 ) );
  nnd2s1 \IDinst/U9501  ( .DIN1(\IDinst/RegFile[20][5] ), .DIN2(n1264), 
        .Q(\IDinst/n9460 ) );
  nnd2s1 \IDinst/U9500  ( .DIN1(\IDinst/n9458 ), .DIN2(\IDinst/n9457 ), 
        .Q(\IDinst/n9459 ) );
  nnd2s1 \IDinst/U9499  ( .DIN1(\IDinst/n9456 ), .DIN2(n1325), 
        .Q(\IDinst/n9458 ) );
  nnd2s1 \IDinst/U9498  ( .DIN1(\IDinst/n9453 ), .DIN2(n1343), 
        .Q(\IDinst/n9457 ) );
  nnd2s1 \IDinst/U9497  ( .DIN1(\IDinst/n9455 ), .DIN2(\IDinst/n9454 ), 
        .Q(\IDinst/n9456 ) );
  nnd2s1 \IDinst/U9496  ( .DIN1(\IDinst/RegFile[19][5] ), .DIN2(n1221), 
        .Q(\IDinst/n9455 ) );
  nnd2s1 \IDinst/U9495  ( .DIN1(\IDinst/RegFile[18][5] ), .DIN2(n1264), 
        .Q(\IDinst/n9454 ) );
  nnd2s1 \IDinst/U9494  ( .DIN1(\IDinst/n9452 ), .DIN2(\IDinst/n9451 ), 
        .Q(\IDinst/n9453 ) );
  nnd2s1 \IDinst/U9493  ( .DIN1(\IDinst/RegFile[17][5] ), .DIN2(n1221), 
        .Q(\IDinst/n9452 ) );
  nnd2s1 \IDinst/U9492  ( .DIN1(\IDinst/RegFile[16][5] ), .DIN2(n1263), 
        .Q(\IDinst/n9451 ) );
  nnd2s1 \IDinst/U9491  ( .DIN1(\IDinst/n9449 ), .DIN2(\IDinst/n9448 ), 
        .Q(\IDinst/n9450 ) );
  nnd2s1 \IDinst/U9490  ( .DIN1(\IDinst/n9447 ), .DIN2(n665), 
        .Q(\IDinst/n9449 ) );
  nnd2s1 \IDinst/U9489  ( .DIN1(\IDinst/n9426 ), .DIN2(n682), 
        .Q(\IDinst/n9448 ) );
  nnd2s1 \IDinst/U9488  ( .DIN1(\IDinst/n9446 ), .DIN2(\IDinst/n9445 ), 
        .Q(\IDinst/n9447 ) );
  nnd2s1 \IDinst/U9487  ( .DIN1(\IDinst/n9444 ), .DIN2(n1379), 
        .Q(\IDinst/n9446 ) );
  nnd2s1 \IDinst/U9486  ( .DIN1(\IDinst/n9435 ), .DIN2(n1369), 
        .Q(\IDinst/n9445 ) );
  nnd2s1 \IDinst/U9485  ( .DIN1(\IDinst/n9443 ), .DIN2(\IDinst/n9442 ), 
        .Q(\IDinst/n9444 ) );
  nnd2s1 \IDinst/U9484  ( .DIN1(\IDinst/n9441 ), .DIN2(n1325), 
        .Q(\IDinst/n9443 ) );
  nnd2s1 \IDinst/U9483  ( .DIN1(\IDinst/n9438 ), .DIN2(n1343), 
        .Q(\IDinst/n9442 ) );
  nnd2s1 \IDinst/U9482  ( .DIN1(\IDinst/n9440 ), .DIN2(\IDinst/n9439 ), 
        .Q(\IDinst/n9441 ) );
  nnd2s1 \IDinst/U9481  ( .DIN1(\IDinst/RegFile[15][5] ), .DIN2(n1221), 
        .Q(\IDinst/n9440 ) );
  nnd2s1 \IDinst/U9480  ( .DIN1(\IDinst/RegFile[14][5] ), .DIN2(n1263), 
        .Q(\IDinst/n9439 ) );
  nnd2s1 \IDinst/U9479  ( .DIN1(\IDinst/n9437 ), .DIN2(\IDinst/n9436 ), 
        .Q(\IDinst/n9438 ) );
  nnd2s1 \IDinst/U9478  ( .DIN1(\IDinst/RegFile[13][5] ), .DIN2(n1221), 
        .Q(\IDinst/n9437 ) );
  nnd2s1 \IDinst/U9477  ( .DIN1(\IDinst/RegFile[12][5] ), .DIN2(n1263), 
        .Q(\IDinst/n9436 ) );
  nnd2s1 \IDinst/U9476  ( .DIN1(\IDinst/n9434 ), .DIN2(\IDinst/n9433 ), 
        .Q(\IDinst/n9435 ) );
  nnd2s1 \IDinst/U9475  ( .DIN1(\IDinst/n9432 ), .DIN2(n1325), 
        .Q(\IDinst/n9434 ) );
  nnd2s1 \IDinst/U9474  ( .DIN1(\IDinst/n9429 ), .DIN2(n1343), 
        .Q(\IDinst/n9433 ) );
  nnd2s1 \IDinst/U9473  ( .DIN1(\IDinst/n9431 ), .DIN2(\IDinst/n9430 ), 
        .Q(\IDinst/n9432 ) );
  nnd2s1 \IDinst/U9472  ( .DIN1(\IDinst/RegFile[11][5] ), .DIN2(n1221), 
        .Q(\IDinst/n9431 ) );
  nnd2s1 \IDinst/U9471  ( .DIN1(\IDinst/RegFile[10][5] ), .DIN2(n1263), 
        .Q(\IDinst/n9430 ) );
  nnd2s1 \IDinst/U9470  ( .DIN1(\IDinst/n9428 ), .DIN2(\IDinst/n9427 ), 
        .Q(\IDinst/n9429 ) );
  nnd2s1 \IDinst/U9469  ( .DIN1(\IDinst/RegFile[9][5] ), .DIN2(n1221), 
        .Q(\IDinst/n9428 ) );
  nnd2s1 \IDinst/U9468  ( .DIN1(\IDinst/RegFile[8][5] ), .DIN2(n1263), 
        .Q(\IDinst/n9427 ) );
  nnd2s1 \IDinst/U9467  ( .DIN1(\IDinst/n9425 ), .DIN2(\IDinst/n9424 ), 
        .Q(\IDinst/n9426 ) );
  nnd2s1 \IDinst/U9466  ( .DIN1(\IDinst/n9423 ), .DIN2(n1379), 
        .Q(\IDinst/n9425 ) );
  nnd2s1 \IDinst/U9465  ( .DIN1(\IDinst/n9414 ), .DIN2(n1368), 
        .Q(\IDinst/n9424 ) );
  nnd2s1 \IDinst/U9464  ( .DIN1(\IDinst/n9422 ), .DIN2(\IDinst/n9421 ), 
        .Q(\IDinst/n9423 ) );
  nnd2s1 \IDinst/U9463  ( .DIN1(\IDinst/n9420 ), .DIN2(n1325), 
        .Q(\IDinst/n9422 ) );
  nnd2s1 \IDinst/U9462  ( .DIN1(\IDinst/n9417 ), .DIN2(n1343), 
        .Q(\IDinst/n9421 ) );
  nnd2s1 \IDinst/U9461  ( .DIN1(\IDinst/n9419 ), .DIN2(\IDinst/n9418 ), 
        .Q(\IDinst/n9420 ) );
  nnd2s1 \IDinst/U9460  ( .DIN1(\IDinst/RegFile[7][5] ), .DIN2(n1221), 
        .Q(\IDinst/n9419 ) );
  nnd2s1 \IDinst/U9459  ( .DIN1(\IDinst/RegFile[6][5] ), .DIN2(n1263), 
        .Q(\IDinst/n9418 ) );
  nnd2s1 \IDinst/U9458  ( .DIN1(\IDinst/n9416 ), .DIN2(\IDinst/n9415 ), 
        .Q(\IDinst/n9417 ) );
  nnd2s1 \IDinst/U9457  ( .DIN1(\IDinst/RegFile[5][5] ), .DIN2(n1221), 
        .Q(\IDinst/n9416 ) );
  nnd2s1 \IDinst/U9456  ( .DIN1(\IDinst/RegFile[4][5] ), .DIN2(n1263), 
        .Q(\IDinst/n9415 ) );
  nnd2s1 \IDinst/U9455  ( .DIN1(\IDinst/n9413 ), .DIN2(\IDinst/n9412 ), 
        .Q(\IDinst/n9414 ) );
  nnd2s1 \IDinst/U9454  ( .DIN1(\IDinst/n9411 ), .DIN2(n1325), 
        .Q(\IDinst/n9413 ) );
  nnd2s1 \IDinst/U9453  ( .DIN1(\IDinst/n9408 ), .DIN2(n1344), 
        .Q(\IDinst/n9412 ) );
  nnd2s1 \IDinst/U9452  ( .DIN1(\IDinst/n9410 ), .DIN2(\IDinst/n9409 ), 
        .Q(\IDinst/n9411 ) );
  nnd2s1 \IDinst/U9451  ( .DIN1(\IDinst/RegFile[3][5] ), .DIN2(n1221), 
        .Q(\IDinst/n9410 ) );
  nnd2s1 \IDinst/U9450  ( .DIN1(\IDinst/RegFile[2][5] ), .DIN2(n1263), 
        .Q(\IDinst/n9409 ) );
  nnd2s1 \IDinst/U9449  ( .DIN1(\IDinst/n9407 ), .DIN2(\IDinst/n9406 ), 
        .Q(\IDinst/n9408 ) );
  nnd2s1 \IDinst/U9448  ( .DIN1(\IDinst/RegFile[1][5] ), .DIN2(n1222), 
        .Q(\IDinst/n9407 ) );
  nnd2s1 \IDinst/U9447  ( .DIN1(\IDinst/RegFile[0][5] ), .DIN2(n1263), 
        .Q(\IDinst/n9406 ) );
  nnd2s1 \IDinst/U9446  ( .DIN1(\IDinst/n9405 ), .DIN2(\IDinst/N48 ), 
        .Q(\IDinst/n8900 ) );
  nnd2s1 \IDinst/U9445  ( .DIN1(\IDinst/n9360 ), .DIN2(n634), 
        .Q(\IDinst/n8901 ) );
  nnd2s1 \IDinst/U9444  ( .DIN1(\IDinst/n9404 ), .DIN2(\IDinst/n9403 ), 
        .Q(\IDinst/n9405 ) );
  nnd2s1 \IDinst/U9443  ( .DIN1(\IDinst/n9402 ), .DIN2(n668), 
        .Q(\IDinst/n9404 ) );
  nnd2s1 \IDinst/U9442  ( .DIN1(\IDinst/n9381 ), .DIN2(n680), 
        .Q(\IDinst/n9403 ) );
  nnd2s1 \IDinst/U9441  ( .DIN1(\IDinst/n9401 ), .DIN2(\IDinst/n9400 ), 
        .Q(\IDinst/n9402 ) );
  nnd2s1 \IDinst/U9440  ( .DIN1(\IDinst/n9399 ), .DIN2(n1378), 
        .Q(\IDinst/n9401 ) );
  nnd2s1 \IDinst/U9439  ( .DIN1(\IDinst/n9390 ), .DIN2(n1367), 
        .Q(\IDinst/n9400 ) );
  nnd2s1 \IDinst/U9438  ( .DIN1(\IDinst/n9398 ), .DIN2(\IDinst/n9397 ), 
        .Q(\IDinst/n9399 ) );
  nnd2s1 \IDinst/U9437  ( .DIN1(\IDinst/n9396 ), .DIN2(n1325), 
        .Q(\IDinst/n9398 ) );
  nnd2s1 \IDinst/U9436  ( .DIN1(\IDinst/n9393 ), .DIN2(n1344), 
        .Q(\IDinst/n9397 ) );
  nnd2s1 \IDinst/U9435  ( .DIN1(\IDinst/n9395 ), .DIN2(\IDinst/n9394 ), 
        .Q(\IDinst/n9396 ) );
  nnd2s1 \IDinst/U9434  ( .DIN1(\IDinst/RegFile[31][4] ), .DIN2(n1222), 
        .Q(\IDinst/n9395 ) );
  nnd2s1 \IDinst/U9433  ( .DIN1(\IDinst/RegFile[30][4] ), .DIN2(n1262), 
        .Q(\IDinst/n9394 ) );
  nnd2s1 \IDinst/U9432  ( .DIN1(\IDinst/n9392 ), .DIN2(\IDinst/n9391 ), 
        .Q(\IDinst/n9393 ) );
  nnd2s1 \IDinst/U9431  ( .DIN1(\IDinst/RegFile[29][4] ), .DIN2(n1222), 
        .Q(\IDinst/n9392 ) );
  nnd2s1 \IDinst/U9430  ( .DIN1(\IDinst/RegFile[28][4] ), .DIN2(n1262), 
        .Q(\IDinst/n9391 ) );
  nnd2s1 \IDinst/U9429  ( .DIN1(\IDinst/n9389 ), .DIN2(\IDinst/n9388 ), 
        .Q(\IDinst/n9390 ) );
  nnd2s1 \IDinst/U9428  ( .DIN1(\IDinst/n9387 ), .DIN2(n1325), 
        .Q(\IDinst/n9389 ) );
  nnd2s1 \IDinst/U9427  ( .DIN1(\IDinst/n9384 ), .DIN2(n1344), 
        .Q(\IDinst/n9388 ) );
  nnd2s1 \IDinst/U9426  ( .DIN1(\IDinst/n9386 ), .DIN2(\IDinst/n9385 ), 
        .Q(\IDinst/n9387 ) );
  nnd2s1 \IDinst/U9425  ( .DIN1(\IDinst/RegFile[27][4] ), .DIN2(n1222), 
        .Q(\IDinst/n9386 ) );
  nnd2s1 \IDinst/U9424  ( .DIN1(\IDinst/RegFile[26][4] ), .DIN2(n1262), 
        .Q(\IDinst/n9385 ) );
  nnd2s1 \IDinst/U9423  ( .DIN1(\IDinst/n9383 ), .DIN2(\IDinst/n9382 ), 
        .Q(\IDinst/n9384 ) );
  nnd2s1 \IDinst/U9422  ( .DIN1(\IDinst/RegFile[25][4] ), .DIN2(n1222), 
        .Q(\IDinst/n9383 ) );
  nnd2s1 \IDinst/U9421  ( .DIN1(\IDinst/RegFile[24][4] ), .DIN2(n1262), 
        .Q(\IDinst/n9382 ) );
  nnd2s1 \IDinst/U9420  ( .DIN1(\IDinst/n9380 ), .DIN2(\IDinst/n9379 ), 
        .Q(\IDinst/n9381 ) );
  nnd2s1 \IDinst/U9419  ( .DIN1(\IDinst/n9378 ), .DIN2(n1377), 
        .Q(\IDinst/n9380 ) );
  nnd2s1 \IDinst/U9418  ( .DIN1(\IDinst/n9369 ), .DIN2(n1366), 
        .Q(\IDinst/n9379 ) );
  nnd2s1 \IDinst/U9417  ( .DIN1(\IDinst/n9377 ), .DIN2(\IDinst/n9376 ), 
        .Q(\IDinst/n9378 ) );
  nnd2s1 \IDinst/U9416  ( .DIN1(\IDinst/n9375 ), .DIN2(n1325), 
        .Q(\IDinst/n9377 ) );
  nnd2s1 \IDinst/U9415  ( .DIN1(\IDinst/n9372 ), .DIN2(n1344), 
        .Q(\IDinst/n9376 ) );
  nnd2s1 \IDinst/U9414  ( .DIN1(\IDinst/n9374 ), .DIN2(\IDinst/n9373 ), 
        .Q(\IDinst/n9375 ) );
  nnd2s1 \IDinst/U9413  ( .DIN1(\IDinst/RegFile[23][4] ), .DIN2(n1222), 
        .Q(\IDinst/n9374 ) );
  nnd2s1 \IDinst/U9412  ( .DIN1(\IDinst/RegFile[22][4] ), .DIN2(n1262), 
        .Q(\IDinst/n9373 ) );
  nnd2s1 \IDinst/U9411  ( .DIN1(\IDinst/n9371 ), .DIN2(\IDinst/n9370 ), 
        .Q(\IDinst/n9372 ) );
  nnd2s1 \IDinst/U9410  ( .DIN1(\IDinst/RegFile[21][4] ), .DIN2(n1222), 
        .Q(\IDinst/n9371 ) );
  nnd2s1 \IDinst/U9409  ( .DIN1(\IDinst/RegFile[20][4] ), .DIN2(n1262), 
        .Q(\IDinst/n9370 ) );
  nnd2s1 \IDinst/U9408  ( .DIN1(\IDinst/n9368 ), .DIN2(\IDinst/n9367 ), 
        .Q(\IDinst/n9369 ) );
  nnd2s1 \IDinst/U9407  ( .DIN1(\IDinst/n9366 ), .DIN2(n1325), 
        .Q(\IDinst/n9368 ) );
  nnd2s1 \IDinst/U9406  ( .DIN1(\IDinst/n9363 ), .DIN2(n1344), 
        .Q(\IDinst/n9367 ) );
  nnd2s1 \IDinst/U9405  ( .DIN1(\IDinst/n9365 ), .DIN2(\IDinst/n9364 ), 
        .Q(\IDinst/n9366 ) );
  nnd2s1 \IDinst/U9404  ( .DIN1(\IDinst/RegFile[19][4] ), .DIN2(n1222), 
        .Q(\IDinst/n9365 ) );
  nnd2s1 \IDinst/U9403  ( .DIN1(\IDinst/RegFile[18][4] ), .DIN2(n1262), 
        .Q(\IDinst/n9364 ) );
  nnd2s1 \IDinst/U9402  ( .DIN1(\IDinst/n9362 ), .DIN2(\IDinst/n9361 ), 
        .Q(\IDinst/n9363 ) );
  nnd2s1 \IDinst/U9401  ( .DIN1(\IDinst/RegFile[17][4] ), .DIN2(n1222), 
        .Q(\IDinst/n9362 ) );
  nnd2s1 \IDinst/U9400  ( .DIN1(\IDinst/RegFile[16][4] ), .DIN2(n1262), 
        .Q(\IDinst/n9361 ) );
  nnd2s1 \IDinst/U9399  ( .DIN1(\IDinst/n9359 ), .DIN2(\IDinst/n9358 ), 
        .Q(\IDinst/n9360 ) );
  nnd2s1 \IDinst/U9398  ( .DIN1(\IDinst/n9357 ), .DIN2(n667), 
        .Q(\IDinst/n9359 ) );
  nnd2s1 \IDinst/U9397  ( .DIN1(\IDinst/n9336 ), .DIN2(n681), 
        .Q(\IDinst/n9358 ) );
  nnd2s1 \IDinst/U9396  ( .DIN1(\IDinst/n9356 ), .DIN2(\IDinst/n9355 ), 
        .Q(\IDinst/n9357 ) );
  nnd2s1 \IDinst/U9395  ( .DIN1(\IDinst/n9354 ), .DIN2(n1374), 
        .Q(\IDinst/n9356 ) );
  nnd2s1 \IDinst/U9394  ( .DIN1(\IDinst/n9345 ), .DIN2(n1365), 
        .Q(\IDinst/n9355 ) );
  nnd2s1 \IDinst/U9393  ( .DIN1(\IDinst/n9353 ), .DIN2(\IDinst/n9352 ), 
        .Q(\IDinst/n9354 ) );
  nnd2s1 \IDinst/U9392  ( .DIN1(\IDinst/n9351 ), .DIN2(n1325), 
        .Q(\IDinst/n9353 ) );
  nnd2s1 \IDinst/U9391  ( .DIN1(\IDinst/n9348 ), .DIN2(n1344), 
        .Q(\IDinst/n9352 ) );
  nnd2s1 \IDinst/U9390  ( .DIN1(\IDinst/n9350 ), .DIN2(\IDinst/n9349 ), 
        .Q(\IDinst/n9351 ) );
  nnd2s1 \IDinst/U9389  ( .DIN1(\IDinst/RegFile[15][4] ), .DIN2(n1222), 
        .Q(\IDinst/n9350 ) );
  nnd2s1 \IDinst/U9388  ( .DIN1(\IDinst/RegFile[14][4] ), .DIN2(n1262), 
        .Q(\IDinst/n9349 ) );
  nnd2s1 \IDinst/U9387  ( .DIN1(\IDinst/n9347 ), .DIN2(\IDinst/n9346 ), 
        .Q(\IDinst/n9348 ) );
  nnd2s1 \IDinst/U9386  ( .DIN1(\IDinst/RegFile[13][4] ), .DIN2(n1222), 
        .Q(\IDinst/n9347 ) );
  nnd2s1 \IDinst/U9385  ( .DIN1(\IDinst/RegFile[12][4] ), .DIN2(n1261), 
        .Q(\IDinst/n9346 ) );
  nnd2s1 \IDinst/U9384  ( .DIN1(\IDinst/n9344 ), .DIN2(\IDinst/n9343 ), 
        .Q(\IDinst/n9345 ) );
  nnd2s1 \IDinst/U9383  ( .DIN1(\IDinst/n9342 ), .DIN2(n1324), 
        .Q(\IDinst/n9344 ) );
  nnd2s1 \IDinst/U9382  ( .DIN1(\IDinst/n9339 ), .DIN2(n1344), 
        .Q(\IDinst/n9343 ) );
  nnd2s1 \IDinst/U9381  ( .DIN1(\IDinst/n9341 ), .DIN2(\IDinst/n9340 ), 
        .Q(\IDinst/n9342 ) );
  nnd2s1 \IDinst/U9380  ( .DIN1(\IDinst/RegFile[11][4] ), .DIN2(n1222), 
        .Q(\IDinst/n9341 ) );
  nnd2s1 \IDinst/U9379  ( .DIN1(\IDinst/RegFile[10][4] ), .DIN2(n1261), 
        .Q(\IDinst/n9340 ) );
  nnd2s1 \IDinst/U9378  ( .DIN1(\IDinst/n9338 ), .DIN2(\IDinst/n9337 ), 
        .Q(\IDinst/n9339 ) );
  nnd2s1 \IDinst/U9377  ( .DIN1(\IDinst/RegFile[9][4] ), .DIN2(n1222), 
        .Q(\IDinst/n9338 ) );
  nnd2s1 \IDinst/U9376  ( .DIN1(\IDinst/RegFile[8][4] ), .DIN2(n1261), 
        .Q(\IDinst/n9337 ) );
  nnd2s1 \IDinst/U9375  ( .DIN1(\IDinst/n9335 ), .DIN2(\IDinst/n9334 ), 
        .Q(\IDinst/n9336 ) );
  nnd2s1 \IDinst/U9374  ( .DIN1(\IDinst/n9333 ), .DIN2(n1372), 
        .Q(\IDinst/n9335 ) );
  nnd2s1 \IDinst/U9373  ( .DIN1(\IDinst/n9324 ), .DIN2(n1365), 
        .Q(\IDinst/n9334 ) );
  nnd2s1 \IDinst/U9372  ( .DIN1(\IDinst/n9332 ), .DIN2(\IDinst/n9331 ), 
        .Q(\IDinst/n9333 ) );
  nnd2s1 \IDinst/U9371  ( .DIN1(\IDinst/n9330 ), .DIN2(n1324), 
        .Q(\IDinst/n9332 ) );
  nnd2s1 \IDinst/U9370  ( .DIN1(\IDinst/n9327 ), .DIN2(n1344), 
        .Q(\IDinst/n9331 ) );
  nnd2s1 \IDinst/U9369  ( .DIN1(\IDinst/n9329 ), .DIN2(\IDinst/n9328 ), 
        .Q(\IDinst/n9330 ) );
  nnd2s1 \IDinst/U9368  ( .DIN1(\IDinst/RegFile[7][4] ), .DIN2(n1223), 
        .Q(\IDinst/n9329 ) );
  nnd2s1 \IDinst/U9367  ( .DIN1(\IDinst/RegFile[6][4] ), .DIN2(n1261), 
        .Q(\IDinst/n9328 ) );
  nnd2s1 \IDinst/U9366  ( .DIN1(\IDinst/n9326 ), .DIN2(\IDinst/n9325 ), 
        .Q(\IDinst/n9327 ) );
  nnd2s1 \IDinst/U9365  ( .DIN1(\IDinst/RegFile[5][4] ), .DIN2(n1223), 
        .Q(\IDinst/n9326 ) );
  nnd2s1 \IDinst/U9364  ( .DIN1(\IDinst/RegFile[4][4] ), .DIN2(n1261), 
        .Q(\IDinst/n9325 ) );
  nnd2s1 \IDinst/U9363  ( .DIN1(\IDinst/n9323 ), .DIN2(\IDinst/n9322 ), 
        .Q(\IDinst/n9324 ) );
  nnd2s1 \IDinst/U9362  ( .DIN1(\IDinst/n9321 ), .DIN2(n1324), 
        .Q(\IDinst/n9323 ) );
  nnd2s1 \IDinst/U9361  ( .DIN1(\IDinst/n9318 ), .DIN2(n1344), 
        .Q(\IDinst/n9322 ) );
  nnd2s1 \IDinst/U9360  ( .DIN1(\IDinst/n9320 ), .DIN2(\IDinst/n9319 ), 
        .Q(\IDinst/n9321 ) );
  nnd2s1 \IDinst/U9359  ( .DIN1(\IDinst/RegFile[3][4] ), .DIN2(n1223), 
        .Q(\IDinst/n9320 ) );
  nnd2s1 \IDinst/U9358  ( .DIN1(\IDinst/RegFile[2][4] ), .DIN2(n1261), 
        .Q(\IDinst/n9319 ) );
  nnd2s1 \IDinst/U9357  ( .DIN1(\IDinst/n9317 ), .DIN2(\IDinst/n9316 ), 
        .Q(\IDinst/n9318 ) );
  nnd2s1 \IDinst/U9356  ( .DIN1(\IDinst/RegFile[1][4] ), .DIN2(n1223), 
        .Q(\IDinst/n9317 ) );
  nnd2s1 \IDinst/U9355  ( .DIN1(\IDinst/RegFile[0][4] ), .DIN2(n1261), 
        .Q(\IDinst/n9316 ) );
  nnd2s1 \IDinst/U9354  ( .DIN1(\IDinst/n9315 ), .DIN2(n535), 
        .Q(\IDinst/n8898 ) );
  nnd2s1 \IDinst/U9353  ( .DIN1(\IDinst/n9270 ), .DIN2(n533), 
        .Q(\IDinst/n8899 ) );
  nnd2s1 \IDinst/U9352  ( .DIN1(\IDinst/n9314 ), .DIN2(\IDinst/n9313 ), 
        .Q(\IDinst/n9315 ) );
  nnd2s1 \IDinst/U9351  ( .DIN1(\IDinst/n9312 ), .DIN2(n665), 
        .Q(\IDinst/n9314 ) );
  nnd2s1 \IDinst/U9350  ( .DIN1(\IDinst/n9291 ), .DIN2(n683), 
        .Q(\IDinst/n9313 ) );
  nnd2s1 \IDinst/U9349  ( .DIN1(\IDinst/n9311 ), .DIN2(\IDinst/n9310 ), 
        .Q(\IDinst/n9312 ) );
  nnd2s1 \IDinst/U9348  ( .DIN1(\IDinst/n9309 ), .DIN2(\IDinst/N46 ), 
        .Q(\IDinst/n9311 ) );
  nnd2s1 \IDinst/U9347  ( .DIN1(\IDinst/n9300 ), .DIN2(n1365), 
        .Q(\IDinst/n9310 ) );
  nnd2s1 \IDinst/U9346  ( .DIN1(\IDinst/n9308 ), .DIN2(\IDinst/n9307 ), 
        .Q(\IDinst/n9309 ) );
  nnd2s1 \IDinst/U9345  ( .DIN1(\IDinst/n9306 ), .DIN2(n1324), 
        .Q(\IDinst/n9308 ) );
  nnd2s1 \IDinst/U9344  ( .DIN1(\IDinst/n9303 ), .DIN2(n1345), 
        .Q(\IDinst/n9307 ) );
  nnd2s1 \IDinst/U9343  ( .DIN1(\IDinst/n9305 ), .DIN2(\IDinst/n9304 ), 
        .Q(\IDinst/n9306 ) );
  nnd2s1 \IDinst/U9342  ( .DIN1(\IDinst/RegFile[31][3] ), .DIN2(n1223), 
        .Q(\IDinst/n9305 ) );
  nnd2s1 \IDinst/U9341  ( .DIN1(\IDinst/RegFile[30][3] ), .DIN2(n1261), 
        .Q(\IDinst/n9304 ) );
  nnd2s1 \IDinst/U9340  ( .DIN1(\IDinst/n9302 ), .DIN2(\IDinst/n9301 ), 
        .Q(\IDinst/n9303 ) );
  nnd2s1 \IDinst/U9339  ( .DIN1(\IDinst/RegFile[29][3] ), .DIN2(n1223), 
        .Q(\IDinst/n9302 ) );
  nnd2s1 \IDinst/U9338  ( .DIN1(\IDinst/RegFile[28][3] ), .DIN2(n1260), 
        .Q(\IDinst/n9301 ) );
  nnd2s1 \IDinst/U9337  ( .DIN1(\IDinst/n9299 ), .DIN2(\IDinst/n9298 ), 
        .Q(\IDinst/n9300 ) );
  nnd2s1 \IDinst/U9336  ( .DIN1(\IDinst/n9297 ), .DIN2(n1324), 
        .Q(\IDinst/n9299 ) );
  nnd2s1 \IDinst/U9335  ( .DIN1(\IDinst/n9294 ), .DIN2(n1345), 
        .Q(\IDinst/n9298 ) );
  nnd2s1 \IDinst/U9334  ( .DIN1(\IDinst/n9296 ), .DIN2(\IDinst/n9295 ), 
        .Q(\IDinst/n9297 ) );
  nnd2s1 \IDinst/U9333  ( .DIN1(\IDinst/RegFile[27][3] ), .DIN2(n1223), 
        .Q(\IDinst/n9296 ) );
  nnd2s1 \IDinst/U9332  ( .DIN1(\IDinst/RegFile[26][3] ), .DIN2(n1260), 
        .Q(\IDinst/n9295 ) );
  nnd2s1 \IDinst/U9331  ( .DIN1(\IDinst/n9293 ), .DIN2(\IDinst/n9292 ), 
        .Q(\IDinst/n9294 ) );
  nnd2s1 \IDinst/U9330  ( .DIN1(\IDinst/RegFile[25][3] ), .DIN2(n1223), 
        .Q(\IDinst/n9293 ) );
  nnd2s1 \IDinst/U9329  ( .DIN1(\IDinst/RegFile[24][3] ), .DIN2(n1260), 
        .Q(\IDinst/n9292 ) );
  nnd2s1 \IDinst/U9328  ( .DIN1(\IDinst/n9290 ), .DIN2(\IDinst/n9289 ), 
        .Q(\IDinst/n9291 ) );
  nnd2s1 \IDinst/U9327  ( .DIN1(\IDinst/n9288 ), .DIN2(n1380), 
        .Q(\IDinst/n9290 ) );
  nnd2s1 \IDinst/U9326  ( .DIN1(\IDinst/n9279 ), .DIN2(n1365), 
        .Q(\IDinst/n9289 ) );
  nnd2s1 \IDinst/U9325  ( .DIN1(\IDinst/n9287 ), .DIN2(\IDinst/n9286 ), 
        .Q(\IDinst/n9288 ) );
  nnd2s1 \IDinst/U9324  ( .DIN1(\IDinst/n9285 ), .DIN2(n1324), 
        .Q(\IDinst/n9287 ) );
  nnd2s1 \IDinst/U9323  ( .DIN1(\IDinst/n9282 ), .DIN2(n1345), 
        .Q(\IDinst/n9286 ) );
  nnd2s1 \IDinst/U9322  ( .DIN1(\IDinst/n9284 ), .DIN2(\IDinst/n9283 ), 
        .Q(\IDinst/n9285 ) );
  nnd2s1 \IDinst/U9321  ( .DIN1(\IDinst/RegFile[23][3] ), .DIN2(n1223), 
        .Q(\IDinst/n9284 ) );
  nnd2s1 \IDinst/U9320  ( .DIN1(\IDinst/RegFile[22][3] ), .DIN2(n1260), 
        .Q(\IDinst/n9283 ) );
  nnd2s1 \IDinst/U9319  ( .DIN1(\IDinst/n9281 ), .DIN2(\IDinst/n9280 ), 
        .Q(\IDinst/n9282 ) );
  nnd2s1 \IDinst/U9318  ( .DIN1(\IDinst/RegFile[21][3] ), .DIN2(n1223), 
        .Q(\IDinst/n9281 ) );
  nnd2s1 \IDinst/U9317  ( .DIN1(\IDinst/RegFile[20][3] ), .DIN2(n1260), 
        .Q(\IDinst/n9280 ) );
  nnd2s1 \IDinst/U9316  ( .DIN1(\IDinst/n9278 ), .DIN2(\IDinst/n9277 ), 
        .Q(\IDinst/n9279 ) );
  nnd2s1 \IDinst/U9315  ( .DIN1(\IDinst/n9276 ), .DIN2(n1324), 
        .Q(\IDinst/n9278 ) );
  nnd2s1 \IDinst/U9314  ( .DIN1(\IDinst/n9273 ), .DIN2(n1345), 
        .Q(\IDinst/n9277 ) );
  nnd2s1 \IDinst/U9313  ( .DIN1(\IDinst/n9275 ), .DIN2(\IDinst/n9274 ), 
        .Q(\IDinst/n9276 ) );
  nnd2s1 \IDinst/U9312  ( .DIN1(\IDinst/RegFile[19][3] ), .DIN2(n1223), 
        .Q(\IDinst/n9275 ) );
  nnd2s1 \IDinst/U9311  ( .DIN1(\IDinst/RegFile[18][3] ), .DIN2(n1260), 
        .Q(\IDinst/n9274 ) );
  nnd2s1 \IDinst/U9310  ( .DIN1(\IDinst/n9272 ), .DIN2(\IDinst/n9271 ), 
        .Q(\IDinst/n9273 ) );
  nnd2s1 \IDinst/U9309  ( .DIN1(\IDinst/RegFile[17][3] ), .DIN2(n1223), 
        .Q(\IDinst/n9272 ) );
  nnd2s1 \IDinst/U9308  ( .DIN1(\IDinst/RegFile[16][3] ), .DIN2(n1260), 
        .Q(\IDinst/n9271 ) );
  nnd2s1 \IDinst/U9307  ( .DIN1(\IDinst/n9269 ), .DIN2(\IDinst/n9268 ), 
        .Q(\IDinst/n9270 ) );
  nnd2s1 \IDinst/U9306  ( .DIN1(\IDinst/n9267 ), .DIN2(n668), 
        .Q(\IDinst/n9269 ) );
  nnd2s1 \IDinst/U9305  ( .DIN1(\IDinst/n9246 ), .DIN2(n682), 
        .Q(\IDinst/n9268 ) );
  nnd2s1 \IDinst/U9304  ( .DIN1(\IDinst/n9266 ), .DIN2(\IDinst/n9265 ), 
        .Q(\IDinst/n9267 ) );
  nnd2s1 \IDinst/U9303  ( .DIN1(\IDinst/n9264 ), .DIN2(n1379), 
        .Q(\IDinst/n9266 ) );
  nnd2s1 \IDinst/U9302  ( .DIN1(\IDinst/n9255 ), .DIN2(n1365), 
        .Q(\IDinst/n9265 ) );
  nnd2s1 \IDinst/U9301  ( .DIN1(\IDinst/n9263 ), .DIN2(\IDinst/n9262 ), 
        .Q(\IDinst/n9264 ) );
  nnd2s1 \IDinst/U9300  ( .DIN1(\IDinst/n9261 ), .DIN2(n1324), 
        .Q(\IDinst/n9263 ) );
  nnd2s1 \IDinst/U9299  ( .DIN1(\IDinst/n9258 ), .DIN2(n1345), 
        .Q(\IDinst/n9262 ) );
  nnd2s1 \IDinst/U9298  ( .DIN1(\IDinst/n9260 ), .DIN2(\IDinst/n9259 ), 
        .Q(\IDinst/n9261 ) );
  nnd2s1 \IDinst/U9297  ( .DIN1(\IDinst/RegFile[15][3] ), .DIN2(n1224), 
        .Q(\IDinst/n9260 ) );
  nnd2s1 \IDinst/U9296  ( .DIN1(\IDinst/RegFile[14][3] ), .DIN2(n1260), 
        .Q(\IDinst/n9259 ) );
  nnd2s1 \IDinst/U9295  ( .DIN1(\IDinst/n9257 ), .DIN2(\IDinst/n9256 ), 
        .Q(\IDinst/n9258 ) );
  nnd2s1 \IDinst/U9294  ( .DIN1(\IDinst/RegFile[13][3] ), .DIN2(n1224), 
        .Q(\IDinst/n9257 ) );
  nnd2s1 \IDinst/U9293  ( .DIN1(\IDinst/RegFile[12][3] ), .DIN2(n1260), 
        .Q(\IDinst/n9256 ) );
  nnd2s1 \IDinst/U9292  ( .DIN1(\IDinst/n9254 ), .DIN2(\IDinst/n9253 ), 
        .Q(\IDinst/n9255 ) );
  nnd2s1 \IDinst/U9291  ( .DIN1(\IDinst/n9252 ), .DIN2(n1324), 
        .Q(\IDinst/n9254 ) );
  nnd2s1 \IDinst/U9290  ( .DIN1(\IDinst/n9249 ), .DIN2(n1345), 
        .Q(\IDinst/n9253 ) );
  nnd2s1 \IDinst/U9289  ( .DIN1(\IDinst/n9251 ), .DIN2(\IDinst/n9250 ), 
        .Q(\IDinst/n9252 ) );
  nnd2s1 \IDinst/U9288  ( .DIN1(\IDinst/RegFile[11][3] ), .DIN2(n1224), 
        .Q(\IDinst/n9251 ) );
  nnd2s1 \IDinst/U9287  ( .DIN1(\IDinst/RegFile[10][3] ), .DIN2(n1259), 
        .Q(\IDinst/n9250 ) );
  nnd2s1 \IDinst/U9286  ( .DIN1(\IDinst/n9248 ), .DIN2(\IDinst/n9247 ), 
        .Q(\IDinst/n9249 ) );
  nnd2s1 \IDinst/U9285  ( .DIN1(\IDinst/RegFile[9][3] ), .DIN2(n1224), 
        .Q(\IDinst/n9248 ) );
  nnd2s1 \IDinst/U9284  ( .DIN1(\IDinst/RegFile[8][3] ), .DIN2(n1259), 
        .Q(\IDinst/n9247 ) );
  nnd2s1 \IDinst/U9283  ( .DIN1(\IDinst/n9245 ), .DIN2(\IDinst/n9244 ), 
        .Q(\IDinst/n9246 ) );
  nnd2s1 \IDinst/U9282  ( .DIN1(\IDinst/n9243 ), .DIN2(n1375), 
        .Q(\IDinst/n9245 ) );
  nnd2s1 \IDinst/U9281  ( .DIN1(\IDinst/n9234 ), .DIN2(n1365), 
        .Q(\IDinst/n9244 ) );
  nnd2s1 \IDinst/U9280  ( .DIN1(\IDinst/n9242 ), .DIN2(\IDinst/n9241 ), 
        .Q(\IDinst/n9243 ) );
  nnd2s1 \IDinst/U9279  ( .DIN1(\IDinst/n9240 ), .DIN2(n1324), 
        .Q(\IDinst/n9242 ) );
  nnd2s1 \IDinst/U9278  ( .DIN1(\IDinst/n9237 ), .DIN2(n1345), 
        .Q(\IDinst/n9241 ) );
  nnd2s1 \IDinst/U9277  ( .DIN1(\IDinst/n9239 ), .DIN2(\IDinst/n9238 ), 
        .Q(\IDinst/n9240 ) );
  nnd2s1 \IDinst/U9276  ( .DIN1(\IDinst/RegFile[7][3] ), .DIN2(n1224), 
        .Q(\IDinst/n9239 ) );
  nnd2s1 \IDinst/U9275  ( .DIN1(\IDinst/RegFile[6][3] ), .DIN2(n1259), 
        .Q(\IDinst/n9238 ) );
  nnd2s1 \IDinst/U9274  ( .DIN1(\IDinst/n9236 ), .DIN2(\IDinst/n9235 ), 
        .Q(\IDinst/n9237 ) );
  nnd2s1 \IDinst/U9273  ( .DIN1(\IDinst/RegFile[5][3] ), .DIN2(n1224), 
        .Q(\IDinst/n9236 ) );
  nnd2s1 \IDinst/U9272  ( .DIN1(\IDinst/RegFile[4][3] ), .DIN2(n1259), 
        .Q(\IDinst/n9235 ) );
  nnd2s1 \IDinst/U9271  ( .DIN1(\IDinst/n9233 ), .DIN2(\IDinst/n9232 ), 
        .Q(\IDinst/n9234 ) );
  nnd2s1 \IDinst/U9270  ( .DIN1(\IDinst/n9231 ), .DIN2(n1324), 
        .Q(\IDinst/n9233 ) );
  nnd2s1 \IDinst/U9269  ( .DIN1(\IDinst/n9228 ), .DIN2(n1345), 
        .Q(\IDinst/n9232 ) );
  nnd2s1 \IDinst/U9268  ( .DIN1(\IDinst/n9230 ), .DIN2(\IDinst/n9229 ), 
        .Q(\IDinst/n9231 ) );
  nnd2s1 \IDinst/U9267  ( .DIN1(\IDinst/RegFile[3][3] ), .DIN2(n1224), 
        .Q(\IDinst/n9230 ) );
  nnd2s1 \IDinst/U9266  ( .DIN1(\IDinst/RegFile[2][3] ), .DIN2(n1259), 
        .Q(\IDinst/n9229 ) );
  nnd2s1 \IDinst/U9265  ( .DIN1(\IDinst/n9227 ), .DIN2(\IDinst/n9226 ), 
        .Q(\IDinst/n9228 ) );
  nnd2s1 \IDinst/U9264  ( .DIN1(\IDinst/RegFile[1][3] ), .DIN2(n1224), 
        .Q(\IDinst/n9227 ) );
  nnd2s1 \IDinst/U9263  ( .DIN1(\IDinst/RegFile[0][3] ), .DIN2(n1259), 
        .Q(\IDinst/n9226 ) );
  nnd2s1 \IDinst/U9262  ( .DIN1(\IDinst/n9225 ), .DIN2(n534), 
        .Q(\IDinst/n8896 ) );
  nnd2s1 \IDinst/U9261  ( .DIN1(\IDinst/n9180 ), .DIN2(n634), 
        .Q(\IDinst/n8897 ) );
  nnd2s1 \IDinst/U9260  ( .DIN1(\IDinst/n9224 ), .DIN2(\IDinst/n9223 ), 
        .Q(\IDinst/n9225 ) );
  nnd2s1 \IDinst/U9259  ( .DIN1(\IDinst/n9222 ), .DIN2(n667), 
        .Q(\IDinst/n9224 ) );
  nnd2s1 \IDinst/U9258  ( .DIN1(\IDinst/n9201 ), .DIN2(n680), 
        .Q(\IDinst/n9223 ) );
  nnd2s1 \IDinst/U9257  ( .DIN1(\IDinst/n9221 ), .DIN2(\IDinst/n9220 ), 
        .Q(\IDinst/n9222 ) );
  nnd2s1 \IDinst/U9256  ( .DIN1(\IDinst/n9219 ), .DIN2(n1373), 
        .Q(\IDinst/n9221 ) );
  nnd2s1 \IDinst/U9255  ( .DIN1(\IDinst/n9210 ), .DIN2(n1365), 
        .Q(\IDinst/n9220 ) );
  nnd2s1 \IDinst/U9254  ( .DIN1(\IDinst/n9218 ), .DIN2(\IDinst/n9217 ), 
        .Q(\IDinst/n9219 ) );
  nnd2s1 \IDinst/U9253  ( .DIN1(\IDinst/n9216 ), .DIN2(n1324), 
        .Q(\IDinst/n9218 ) );
  nnd2s1 \IDinst/U9252  ( .DIN1(\IDinst/n9213 ), .DIN2(n1345), 
        .Q(\IDinst/n9217 ) );
  nnd2s1 \IDinst/U9251  ( .DIN1(\IDinst/n9215 ), .DIN2(\IDinst/n9214 ), 
        .Q(\IDinst/n9216 ) );
  nnd2s1 \IDinst/U9250  ( .DIN1(\IDinst/RegFile[31][2] ), .DIN2(n1224), 
        .Q(\IDinst/n9215 ) );
  nnd2s1 \IDinst/U9249  ( .DIN1(\IDinst/RegFile[30][2] ), .DIN2(n1259), 
        .Q(\IDinst/n9214 ) );
  nnd2s1 \IDinst/U9248  ( .DIN1(\IDinst/n9212 ), .DIN2(\IDinst/n9211 ), 
        .Q(\IDinst/n9213 ) );
  nnd2s1 \IDinst/U9247  ( .DIN1(\IDinst/RegFile[29][2] ), .DIN2(n1224), 
        .Q(\IDinst/n9212 ) );
  nnd2s1 \IDinst/U9246  ( .DIN1(\IDinst/RegFile[28][2] ), .DIN2(n1259), 
        .Q(\IDinst/n9211 ) );
  nnd2s1 \IDinst/U9245  ( .DIN1(\IDinst/n9209 ), .DIN2(\IDinst/n9208 ), 
        .Q(\IDinst/n9210 ) );
  nnd2s1 \IDinst/U9244  ( .DIN1(\IDinst/n9207 ), .DIN2(n1324), 
        .Q(\IDinst/n9209 ) );
  nnd2s1 \IDinst/U9243  ( .DIN1(\IDinst/n9204 ), .DIN2(n1346), 
        .Q(\IDinst/n9208 ) );
  nnd2s1 \IDinst/U9242  ( .DIN1(\IDinst/n9206 ), .DIN2(\IDinst/n9205 ), 
        .Q(\IDinst/n9207 ) );
  nnd2s1 \IDinst/U9241  ( .DIN1(\IDinst/RegFile[27][2] ), .DIN2(n1224), 
        .Q(\IDinst/n9206 ) );
  nnd2s1 \IDinst/U9240  ( .DIN1(\IDinst/RegFile[26][2] ), .DIN2(n1259), 
        .Q(\IDinst/n9205 ) );
  nnd2s1 \IDinst/U9239  ( .DIN1(\IDinst/n9203 ), .DIN2(\IDinst/n9202 ), 
        .Q(\IDinst/n9204 ) );
  nnd2s1 \IDinst/U9238  ( .DIN1(\IDinst/RegFile[25][2] ), .DIN2(n1224), 
        .Q(\IDinst/n9203 ) );
  nnd2s1 \IDinst/U9237  ( .DIN1(\IDinst/RegFile[24][2] ), .DIN2(n1258), 
        .Q(\IDinst/n9202 ) );
  nnd2s1 \IDinst/U9236  ( .DIN1(\IDinst/n9200 ), .DIN2(\IDinst/n9199 ), 
        .Q(\IDinst/n9201 ) );
  nnd2s1 \IDinst/U9235  ( .DIN1(\IDinst/n9198 ), .DIN2(n1380), 
        .Q(\IDinst/n9200 ) );
  nnd2s1 \IDinst/U9234  ( .DIN1(\IDinst/n9189 ), .DIN2(n1365), 
        .Q(\IDinst/n9199 ) );
  nnd2s1 \IDinst/U9233  ( .DIN1(\IDinst/n9197 ), .DIN2(\IDinst/n9196 ), 
        .Q(\IDinst/n9198 ) );
  nnd2s1 \IDinst/U9232  ( .DIN1(\IDinst/n9195 ), .DIN2(n1323), 
        .Q(\IDinst/n9197 ) );
  nnd2s1 \IDinst/U9231  ( .DIN1(\IDinst/n9192 ), .DIN2(n1346), 
        .Q(\IDinst/n9196 ) );
  nnd2s1 \IDinst/U9230  ( .DIN1(\IDinst/n9194 ), .DIN2(\IDinst/n9193 ), 
        .Q(\IDinst/n9195 ) );
  nnd2s1 \IDinst/U9229  ( .DIN1(\IDinst/RegFile[23][2] ), .DIN2(n1224), 
        .Q(\IDinst/n9194 ) );
  nnd2s1 \IDinst/U9228  ( .DIN1(\IDinst/RegFile[22][2] ), .DIN2(n1258), 
        .Q(\IDinst/n9193 ) );
  nnd2s1 \IDinst/U9227  ( .DIN1(\IDinst/n9191 ), .DIN2(\IDinst/n9190 ), 
        .Q(\IDinst/n9192 ) );
  nnd2s1 \IDinst/U9226  ( .DIN1(\IDinst/RegFile[21][2] ), .DIN2(n1225), 
        .Q(\IDinst/n9191 ) );
  nnd2s1 \IDinst/U9225  ( .DIN1(\IDinst/RegFile[20][2] ), .DIN2(n1258), 
        .Q(\IDinst/n9190 ) );
  nnd2s1 \IDinst/U9224  ( .DIN1(\IDinst/n9188 ), .DIN2(\IDinst/n9187 ), 
        .Q(\IDinst/n9189 ) );
  nnd2s1 \IDinst/U9223  ( .DIN1(\IDinst/n9186 ), .DIN2(n1323), 
        .Q(\IDinst/n9188 ) );
  nnd2s1 \IDinst/U9222  ( .DIN1(\IDinst/n9183 ), .DIN2(n1346), 
        .Q(\IDinst/n9187 ) );
  nnd2s1 \IDinst/U9221  ( .DIN1(\IDinst/n9185 ), .DIN2(\IDinst/n9184 ), 
        .Q(\IDinst/n9186 ) );
  nnd2s1 \IDinst/U9220  ( .DIN1(\IDinst/RegFile[19][2] ), .DIN2(n1225), 
        .Q(\IDinst/n9185 ) );
  nnd2s1 \IDinst/U9219  ( .DIN1(\IDinst/RegFile[18][2] ), .DIN2(n1258), 
        .Q(\IDinst/n9184 ) );
  nnd2s1 \IDinst/U9218  ( .DIN1(\IDinst/n9182 ), .DIN2(\IDinst/n9181 ), 
        .Q(\IDinst/n9183 ) );
  nnd2s1 \IDinst/U9217  ( .DIN1(\IDinst/RegFile[17][2] ), .DIN2(n1225), 
        .Q(\IDinst/n9182 ) );
  nnd2s1 \IDinst/U9216  ( .DIN1(\IDinst/RegFile[16][2] ), .DIN2(n1258), 
        .Q(\IDinst/n9181 ) );
  nnd2s1 \IDinst/U9215  ( .DIN1(\IDinst/n9179 ), .DIN2(\IDinst/n9178 ), 
        .Q(\IDinst/n9180 ) );
  nnd2s1 \IDinst/U9214  ( .DIN1(\IDinst/n9177 ), .DIN2(n665), 
        .Q(\IDinst/n9179 ) );
  nnd2s1 \IDinst/U9213  ( .DIN1(\IDinst/n9156 ), .DIN2(n681), 
        .Q(\IDinst/n9178 ) );
  nnd2s1 \IDinst/U9212  ( .DIN1(\IDinst/n9176 ), .DIN2(\IDinst/n9175 ), 
        .Q(\IDinst/n9177 ) );
  nnd2s1 \IDinst/U9211  ( .DIN1(\IDinst/n9174 ), .DIN2(n1380), 
        .Q(\IDinst/n9176 ) );
  nnd2s1 \IDinst/U9210  ( .DIN1(\IDinst/n9165 ), .DIN2(n1365), 
        .Q(\IDinst/n9175 ) );
  nnd2s1 \IDinst/U9209  ( .DIN1(\IDinst/n9173 ), .DIN2(\IDinst/n9172 ), 
        .Q(\IDinst/n9174 ) );
  nnd2s1 \IDinst/U9208  ( .DIN1(\IDinst/n9171 ), .DIN2(n1323), 
        .Q(\IDinst/n9173 ) );
  nnd2s1 \IDinst/U9207  ( .DIN1(\IDinst/n9168 ), .DIN2(n1346), 
        .Q(\IDinst/n9172 ) );
  nnd2s1 \IDinst/U9206  ( .DIN1(\IDinst/n9170 ), .DIN2(\IDinst/n9169 ), 
        .Q(\IDinst/n9171 ) );
  nnd2s1 \IDinst/U9205  ( .DIN1(\IDinst/RegFile[15][2] ), .DIN2(n1225), 
        .Q(\IDinst/n9170 ) );
  nnd2s1 \IDinst/U9204  ( .DIN1(\IDinst/RegFile[14][2] ), .DIN2(n1258), 
        .Q(\IDinst/n9169 ) );
  nnd2s1 \IDinst/U9203  ( .DIN1(\IDinst/n9167 ), .DIN2(\IDinst/n9166 ), 
        .Q(\IDinst/n9168 ) );
  nnd2s1 \IDinst/U9202  ( .DIN1(\IDinst/RegFile[13][2] ), .DIN2(n1225), 
        .Q(\IDinst/n9167 ) );
  nnd2s1 \IDinst/U9201  ( .DIN1(\IDinst/RegFile[12][2] ), .DIN2(n1258), 
        .Q(\IDinst/n9166 ) );
  nnd2s1 \IDinst/U9200  ( .DIN1(\IDinst/n9164 ), .DIN2(\IDinst/n9163 ), 
        .Q(\IDinst/n9165 ) );
  nnd2s1 \IDinst/U9199  ( .DIN1(\IDinst/n9162 ), .DIN2(n1323), 
        .Q(\IDinst/n9164 ) );
  nnd2s1 \IDinst/U9198  ( .DIN1(\IDinst/n9159 ), .DIN2(n1346), 
        .Q(\IDinst/n9163 ) );
  nnd2s1 \IDinst/U9197  ( .DIN1(\IDinst/n9161 ), .DIN2(\IDinst/n9160 ), 
        .Q(\IDinst/n9162 ) );
  nnd2s1 \IDinst/U9196  ( .DIN1(\IDinst/RegFile[11][2] ), .DIN2(n1225), 
        .Q(\IDinst/n9161 ) );
  nnd2s1 \IDinst/U9195  ( .DIN1(\IDinst/RegFile[10][2] ), .DIN2(n1258), 
        .Q(\IDinst/n9160 ) );
  nnd2s1 \IDinst/U9194  ( .DIN1(\IDinst/n9158 ), .DIN2(\IDinst/n9157 ), 
        .Q(\IDinst/n9159 ) );
  nnd2s1 \IDinst/U9193  ( .DIN1(\IDinst/RegFile[9][2] ), .DIN2(n1225), 
        .Q(\IDinst/n9158 ) );
  nnd2s1 \IDinst/U9192  ( .DIN1(\IDinst/RegFile[8][2] ), .DIN2(n1258), 
        .Q(\IDinst/n9157 ) );
  nnd2s1 \IDinst/U9191  ( .DIN1(\IDinst/n9155 ), .DIN2(\IDinst/n9154 ), 
        .Q(\IDinst/n9156 ) );
  nnd2s1 \IDinst/U9190  ( .DIN1(\IDinst/n9153 ), .DIN2(n1380), 
        .Q(\IDinst/n9155 ) );
  nnd2s1 \IDinst/U9189  ( .DIN1(\IDinst/n9144 ), .DIN2(n1365), 
        .Q(\IDinst/n9154 ) );
  nnd2s1 \IDinst/U9188  ( .DIN1(\IDinst/n9152 ), .DIN2(\IDinst/n9151 ), 
        .Q(\IDinst/n9153 ) );
  nnd2s1 \IDinst/U9187  ( .DIN1(\IDinst/n9150 ), .DIN2(n1323), 
        .Q(\IDinst/n9152 ) );
  nnd2s1 \IDinst/U9186  ( .DIN1(\IDinst/n9147 ), .DIN2(n1346), 
        .Q(\IDinst/n9151 ) );
  nnd2s1 \IDinst/U9185  ( .DIN1(\IDinst/n9149 ), .DIN2(\IDinst/n9148 ), 
        .Q(\IDinst/n9150 ) );
  nnd2s1 \IDinst/U9184  ( .DIN1(\IDinst/RegFile[7][2] ), .DIN2(n1225), 
        .Q(\IDinst/n9149 ) );
  nnd2s1 \IDinst/U9183  ( .DIN1(\IDinst/RegFile[6][2] ), .DIN2(n1257), 
        .Q(\IDinst/n9148 ) );
  nnd2s1 \IDinst/U9182  ( .DIN1(\IDinst/n9146 ), .DIN2(\IDinst/n9145 ), 
        .Q(\IDinst/n9147 ) );
  nnd2s1 \IDinst/U9181  ( .DIN1(\IDinst/RegFile[5][2] ), .DIN2(n1225), 
        .Q(\IDinst/n9146 ) );
  nnd2s1 \IDinst/U9180  ( .DIN1(\IDinst/RegFile[4][2] ), .DIN2(n1257), 
        .Q(\IDinst/n9145 ) );
  nnd2s1 \IDinst/U9179  ( .DIN1(\IDinst/n9143 ), .DIN2(\IDinst/n9142 ), 
        .Q(\IDinst/n9144 ) );
  nnd2s1 \IDinst/U9178  ( .DIN1(\IDinst/n9141 ), .DIN2(n1323), 
        .Q(\IDinst/n9143 ) );
  nnd2s1 \IDinst/U9177  ( .DIN1(\IDinst/n9138 ), .DIN2(n1346), 
        .Q(\IDinst/n9142 ) );
  nnd2s1 \IDinst/U9176  ( .DIN1(\IDinst/n9140 ), .DIN2(\IDinst/n9139 ), 
        .Q(\IDinst/n9141 ) );
  nnd2s1 \IDinst/U9175  ( .DIN1(\IDinst/RegFile[3][2] ), .DIN2(n1225), 
        .Q(\IDinst/n9140 ) );
  nnd2s1 \IDinst/U9174  ( .DIN1(\IDinst/RegFile[2][2] ), .DIN2(n1257), 
        .Q(\IDinst/n9139 ) );
  nnd2s1 \IDinst/U9173  ( .DIN1(\IDinst/n9137 ), .DIN2(\IDinst/n9136 ), 
        .Q(\IDinst/n9138 ) );
  nnd2s1 \IDinst/U9172  ( .DIN1(\IDinst/RegFile[1][2] ), .DIN2(n1225), 
        .Q(\IDinst/n9137 ) );
  nnd2s1 \IDinst/U9171  ( .DIN1(\IDinst/RegFile[0][2] ), .DIN2(n1257), 
        .Q(\IDinst/n9136 ) );
  nnd2s1 \IDinst/U9170  ( .DIN1(\IDinst/n9135 ), .DIN2(\IDinst/N48 ), 
        .Q(\IDinst/n8894 ) );
  nnd2s1 \IDinst/U9169  ( .DIN1(\IDinst/n9090 ), .DIN2(n533), 
        .Q(\IDinst/n8895 ) );
  nnd2s1 \IDinst/U9168  ( .DIN1(\IDinst/n9134 ), .DIN2(\IDinst/n9133 ), 
        .Q(\IDinst/n9135 ) );
  nnd2s1 \IDinst/U9167  ( .DIN1(\IDinst/n9132 ), .DIN2(n668), 
        .Q(\IDinst/n9134 ) );
  nnd2s1 \IDinst/U9166  ( .DIN1(\IDinst/n9111 ), .DIN2(n683), 
        .Q(\IDinst/n9133 ) );
  nnd2s1 \IDinst/U9165  ( .DIN1(\IDinst/n9131 ), .DIN2(\IDinst/n9130 ), 
        .Q(\IDinst/n9132 ) );
  nnd2s1 \IDinst/U9164  ( .DIN1(\IDinst/n9129 ), .DIN2(n1380), 
        .Q(\IDinst/n9131 ) );
  nnd2s1 \IDinst/U9163  ( .DIN1(\IDinst/n9120 ), .DIN2(n1365), 
        .Q(\IDinst/n9130 ) );
  nnd2s1 \IDinst/U9162  ( .DIN1(\IDinst/n9128 ), .DIN2(\IDinst/n9127 ), 
        .Q(\IDinst/n9129 ) );
  nnd2s1 \IDinst/U9161  ( .DIN1(\IDinst/n9126 ), .DIN2(n1323), 
        .Q(\IDinst/n9128 ) );
  nnd2s1 \IDinst/U9160  ( .DIN1(\IDinst/n9123 ), .DIN2(n1346), 
        .Q(\IDinst/n9127 ) );
  nnd2s1 \IDinst/U9159  ( .DIN1(\IDinst/n9125 ), .DIN2(\IDinst/n9124 ), 
        .Q(\IDinst/n9126 ) );
  nnd2s1 \IDinst/U9158  ( .DIN1(\IDinst/RegFile[31][1] ), .DIN2(n1225), 
        .Q(\IDinst/n9125 ) );
  nnd2s1 \IDinst/U9157  ( .DIN1(\IDinst/RegFile[30][1] ), .DIN2(n1257), 
        .Q(\IDinst/n9124 ) );
  nnd2s1 \IDinst/U9156  ( .DIN1(\IDinst/n9122 ), .DIN2(\IDinst/n9121 ), 
        .Q(\IDinst/n9123 ) );
  nnd2s1 \IDinst/U9155  ( .DIN1(\IDinst/RegFile[29][1] ), .DIN2(n1225), 
        .Q(\IDinst/n9122 ) );
  nnd2s1 \IDinst/U9154  ( .DIN1(\IDinst/RegFile[28][1] ), .DIN2(n1257), 
        .Q(\IDinst/n9121 ) );
  nnd2s1 \IDinst/U9153  ( .DIN1(\IDinst/n9119 ), .DIN2(\IDinst/n9118 ), 
        .Q(\IDinst/n9120 ) );
  nnd2s1 \IDinst/U9152  ( .DIN1(\IDinst/n9117 ), .DIN2(n1323), 
        .Q(\IDinst/n9119 ) );
  nnd2s1 \IDinst/U9151  ( .DIN1(\IDinst/n9114 ), .DIN2(n1346), 
        .Q(\IDinst/n9118 ) );
  nnd2s1 \IDinst/U9150  ( .DIN1(\IDinst/n9116 ), .DIN2(\IDinst/n9115 ), 
        .Q(\IDinst/n9117 ) );
  nnd2s1 \IDinst/U9149  ( .DIN1(\IDinst/RegFile[27][1] ), .DIN2(n1226), 
        .Q(\IDinst/n9116 ) );
  nnd2s1 \IDinst/U9148  ( .DIN1(\IDinst/RegFile[26][1] ), .DIN2(n1257), 
        .Q(\IDinst/n9115 ) );
  nnd2s1 \IDinst/U9147  ( .DIN1(\IDinst/n9113 ), .DIN2(\IDinst/n9112 ), 
        .Q(\IDinst/n9114 ) );
  nnd2s1 \IDinst/U9146  ( .DIN1(\IDinst/RegFile[25][1] ), .DIN2(n1226), 
        .Q(\IDinst/n9113 ) );
  nnd2s1 \IDinst/U9145  ( .DIN1(\IDinst/RegFile[24][1] ), .DIN2(n1257), 
        .Q(\IDinst/n9112 ) );
  nnd2s1 \IDinst/U9144  ( .DIN1(\IDinst/n9110 ), .DIN2(\IDinst/n9109 ), 
        .Q(\IDinst/n9111 ) );
  nnd2s1 \IDinst/U9143  ( .DIN1(\IDinst/n9108 ), .DIN2(n1380), 
        .Q(\IDinst/n9110 ) );
  nnd2s1 \IDinst/U9142  ( .DIN1(\IDinst/n9099 ), .DIN2(n1365), 
        .Q(\IDinst/n9109 ) );
  nnd2s1 \IDinst/U9141  ( .DIN1(\IDinst/n9107 ), .DIN2(\IDinst/n9106 ), 
        .Q(\IDinst/n9108 ) );
  nnd2s1 \IDinst/U9140  ( .DIN1(\IDinst/n9105 ), .DIN2(n1323), 
        .Q(\IDinst/n9107 ) );
  nnd2s1 \IDinst/U9139  ( .DIN1(\IDinst/n9102 ), .DIN2(n1347), 
        .Q(\IDinst/n9106 ) );
  nnd2s1 \IDinst/U9138  ( .DIN1(\IDinst/n9104 ), .DIN2(\IDinst/n9103 ), 
        .Q(\IDinst/n9105 ) );
  nnd2s1 \IDinst/U9137  ( .DIN1(\IDinst/RegFile[23][1] ), .DIN2(n1226), 
        .Q(\IDinst/n9104 ) );
  nnd2s1 \IDinst/U9136  ( .DIN1(\IDinst/RegFile[22][1] ), .DIN2(n1257), 
        .Q(\IDinst/n9103 ) );
  nnd2s1 \IDinst/U9135  ( .DIN1(\IDinst/n9101 ), .DIN2(\IDinst/n9100 ), 
        .Q(\IDinst/n9102 ) );
  nnd2s1 \IDinst/U9134  ( .DIN1(\IDinst/RegFile[21][1] ), .DIN2(n1226), 
        .Q(\IDinst/n9101 ) );
  nnd2s1 \IDinst/U9133  ( .DIN1(\IDinst/RegFile[20][1] ), .DIN2(n1256), 
        .Q(\IDinst/n9100 ) );
  nnd2s1 \IDinst/U9132  ( .DIN1(\IDinst/n9098 ), .DIN2(\IDinst/n9097 ), 
        .Q(\IDinst/n9099 ) );
  nnd2s1 \IDinst/U9131  ( .DIN1(\IDinst/n9096 ), .DIN2(n1323), 
        .Q(\IDinst/n9098 ) );
  nnd2s1 \IDinst/U9130  ( .DIN1(\IDinst/n9093 ), .DIN2(n1347), 
        .Q(\IDinst/n9097 ) );
  nnd2s1 \IDinst/U9129  ( .DIN1(\IDinst/n9095 ), .DIN2(\IDinst/n9094 ), 
        .Q(\IDinst/n9096 ) );
  nnd2s1 \IDinst/U9128  ( .DIN1(\IDinst/RegFile[19][1] ), .DIN2(n1226), 
        .Q(\IDinst/n9095 ) );
  nnd2s1 \IDinst/U9127  ( .DIN1(\IDinst/RegFile[18][1] ), .DIN2(n1256), 
        .Q(\IDinst/n9094 ) );
  nnd2s1 \IDinst/U9126  ( .DIN1(\IDinst/n9092 ), .DIN2(\IDinst/n9091 ), 
        .Q(\IDinst/n9093 ) );
  nnd2s1 \IDinst/U9125  ( .DIN1(\IDinst/RegFile[17][1] ), .DIN2(n1226), 
        .Q(\IDinst/n9092 ) );
  nnd2s1 \IDinst/U9124  ( .DIN1(\IDinst/RegFile[16][1] ), .DIN2(n1256), 
        .Q(\IDinst/n9091 ) );
  nnd2s1 \IDinst/U9123  ( .DIN1(\IDinst/n9089 ), .DIN2(\IDinst/n9088 ), 
        .Q(\IDinst/n9090 ) );
  nnd2s1 \IDinst/U9122  ( .DIN1(\IDinst/n9087 ), .DIN2(n665), 
        .Q(\IDinst/n9089 ) );
  nnd2s1 \IDinst/U9121  ( .DIN1(\IDinst/n9066 ), .DIN2(n682), 
        .Q(\IDinst/n9088 ) );
  nnd2s1 \IDinst/U9120  ( .DIN1(\IDinst/n9086 ), .DIN2(\IDinst/n9085 ), 
        .Q(\IDinst/n9087 ) );
  nnd2s1 \IDinst/U9119  ( .DIN1(\IDinst/n9084 ), .DIN2(n1380), 
        .Q(\IDinst/n9086 ) );
  nnd2s1 \IDinst/U9118  ( .DIN1(\IDinst/n9075 ), .DIN2(n1365), 
        .Q(\IDinst/n9085 ) );
  nnd2s1 \IDinst/U9117  ( .DIN1(\IDinst/n9083 ), .DIN2(\IDinst/n9082 ), 
        .Q(\IDinst/n9084 ) );
  nnd2s1 \IDinst/U9116  ( .DIN1(\IDinst/n9081 ), .DIN2(n1323), 
        .Q(\IDinst/n9083 ) );
  nnd2s1 \IDinst/U9115  ( .DIN1(\IDinst/n9078 ), .DIN2(n1347), 
        .Q(\IDinst/n9082 ) );
  nnd2s1 \IDinst/U9114  ( .DIN1(\IDinst/n9080 ), .DIN2(\IDinst/n9079 ), 
        .Q(\IDinst/n9081 ) );
  nnd2s1 \IDinst/U9113  ( .DIN1(\IDinst/RegFile[15][1] ), .DIN2(n1226), 
        .Q(\IDinst/n9080 ) );
  nnd2s1 \IDinst/U9112  ( .DIN1(\IDinst/RegFile[14][1] ), .DIN2(n1256), 
        .Q(\IDinst/n9079 ) );
  nnd2s1 \IDinst/U9111  ( .DIN1(\IDinst/n9077 ), .DIN2(\IDinst/n9076 ), 
        .Q(\IDinst/n9078 ) );
  nnd2s1 \IDinst/U9110  ( .DIN1(\IDinst/RegFile[13][1] ), .DIN2(n1226), 
        .Q(\IDinst/n9077 ) );
  nnd2s1 \IDinst/U9109  ( .DIN1(\IDinst/RegFile[12][1] ), .DIN2(n1256), 
        .Q(\IDinst/n9076 ) );
  nnd2s1 \IDinst/U9108  ( .DIN1(\IDinst/n9074 ), .DIN2(\IDinst/n9073 ), 
        .Q(\IDinst/n9075 ) );
  nnd2s1 \IDinst/U9107  ( .DIN1(\IDinst/n9072 ), .DIN2(n1323), 
        .Q(\IDinst/n9074 ) );
  nnd2s1 \IDinst/U9106  ( .DIN1(\IDinst/n9069 ), .DIN2(n1347), 
        .Q(\IDinst/n9073 ) );
  nnd2s1 \IDinst/U9105  ( .DIN1(\IDinst/n9071 ), .DIN2(\IDinst/n9070 ), 
        .Q(\IDinst/n9072 ) );
  nnd2s1 \IDinst/U9104  ( .DIN1(\IDinst/RegFile[11][1] ), .DIN2(n1226), 
        .Q(\IDinst/n9071 ) );
  nnd2s1 \IDinst/U9103  ( .DIN1(\IDinst/RegFile[10][1] ), .DIN2(n1256), 
        .Q(\IDinst/n9070 ) );
  nnd2s1 \IDinst/U9102  ( .DIN1(\IDinst/n9068 ), .DIN2(\IDinst/n9067 ), 
        .Q(\IDinst/n9069 ) );
  nnd2s1 \IDinst/U9101  ( .DIN1(\IDinst/RegFile[9][1] ), .DIN2(n1226), 
        .Q(\IDinst/n9068 ) );
  nnd2s1 \IDinst/U9100  ( .DIN1(\IDinst/RegFile[8][1] ), .DIN2(n1256), 
        .Q(\IDinst/n9067 ) );
  nnd2s1 \IDinst/U9099  ( .DIN1(\IDinst/n9065 ), .DIN2(\IDinst/n9064 ), 
        .Q(\IDinst/n9066 ) );
  nnd2s1 \IDinst/U9098  ( .DIN1(\IDinst/n9063 ), .DIN2(n1380), 
        .Q(\IDinst/n9065 ) );
  nnd2s1 \IDinst/U9097  ( .DIN1(\IDinst/n9054 ), .DIN2(n1365), 
        .Q(\IDinst/n9064 ) );
  nnd2s1 \IDinst/U9096  ( .DIN1(\IDinst/n9062 ), .DIN2(\IDinst/n9061 ), 
        .Q(\IDinst/n9063 ) );
  nnd2s1 \IDinst/U9095  ( .DIN1(\IDinst/n9060 ), .DIN2(n1323), 
        .Q(\IDinst/n9062 ) );
  nnd2s1 \IDinst/U9094  ( .DIN1(\IDinst/n9057 ), .DIN2(n1347), 
        .Q(\IDinst/n9061 ) );
  nnd2s1 \IDinst/U9093  ( .DIN1(\IDinst/n9059 ), .DIN2(\IDinst/n9058 ), 
        .Q(\IDinst/n9060 ) );
  nnd2s1 \IDinst/U9092  ( .DIN1(\IDinst/RegFile[7][1] ), .DIN2(n1226), 
        .Q(\IDinst/n9059 ) );
  nnd2s1 \IDinst/U9091  ( .DIN1(\IDinst/RegFile[6][1] ), .DIN2(n1256), 
        .Q(\IDinst/n9058 ) );
  nnd2s1 \IDinst/U9090  ( .DIN1(\IDinst/n9056 ), .DIN2(\IDinst/n9055 ), 
        .Q(\IDinst/n9057 ) );
  nnd2s1 \IDinst/U9089  ( .DIN1(\IDinst/RegFile[5][1] ), .DIN2(n1226), 
        .Q(\IDinst/n9056 ) );
  nnd2s1 \IDinst/U9088  ( .DIN1(\IDinst/RegFile[4][1] ), .DIN2(n1256), 
        .Q(\IDinst/n9055 ) );
  nnd2s1 \IDinst/U9087  ( .DIN1(\IDinst/n9053 ), .DIN2(\IDinst/n9052 ), 
        .Q(\IDinst/n9054 ) );
  nnd2s1 \IDinst/U9086  ( .DIN1(\IDinst/n9051 ), .DIN2(n1322), 
        .Q(\IDinst/n9053 ) );
  nnd2s1 \IDinst/U9085  ( .DIN1(\IDinst/n9048 ), .DIN2(n1347), 
        .Q(\IDinst/n9052 ) );
  nnd2s1 \IDinst/U9084  ( .DIN1(\IDinst/n9050 ), .DIN2(\IDinst/n9049 ), 
        .Q(\IDinst/n9051 ) );
  nnd2s1 \IDinst/U9083  ( .DIN1(\IDinst/RegFile[3][1] ), .DIN2(n1226), 
        .Q(\IDinst/n9050 ) );
  nnd2s1 \IDinst/U9082  ( .DIN1(\IDinst/RegFile[2][1] ), .DIN2(n1255), 
        .Q(\IDinst/n9049 ) );
  nnd2s1 \IDinst/U9081  ( .DIN1(\IDinst/n9047 ), .DIN2(\IDinst/n9046 ), 
        .Q(\IDinst/n9048 ) );
  nnd2s1 \IDinst/U9080  ( .DIN1(\IDinst/RegFile[1][1] ), .DIN2(n1227), 
        .Q(\IDinst/n9047 ) );
  nnd2s1 \IDinst/U9079  ( .DIN1(\IDinst/RegFile[0][1] ), .DIN2(n1255), 
        .Q(\IDinst/n9046 ) );
  nnd2s1 \IDinst/U9078  ( .DIN1(n535), .DIN2(\IDinst/n9045 ), 
        .Q(\IDinst/n8892 ) );
  nnd2s1 \IDinst/U9077  ( .DIN1(\IDinst/n9000 ), .DIN2(n634), 
        .Q(\IDinst/n8893 ) );
  nnd2s1 \IDinst/U9076  ( .DIN1(\IDinst/n9044 ), .DIN2(\IDinst/n9043 ), 
        .Q(\IDinst/n9045 ) );
  nnd2s1 \IDinst/U9075  ( .DIN1(\IDinst/n9042 ), .DIN2(n668), 
        .Q(\IDinst/n9044 ) );
  nnd2s1 \IDinst/U9074  ( .DIN1(\IDinst/n9021 ), .DIN2(n680), 
        .Q(\IDinst/n9043 ) );
  nnd2s1 \IDinst/U9073  ( .DIN1(\IDinst/n9041 ), .DIN2(\IDinst/n9040 ), 
        .Q(\IDinst/n9042 ) );
  nnd2s1 \IDinst/U9072  ( .DIN1(\IDinst/n9039 ), .DIN2(n1380), 
        .Q(\IDinst/n9041 ) );
  nnd2s1 \IDinst/U9071  ( .DIN1(\IDinst/n9030 ), .DIN2(n1364), 
        .Q(\IDinst/n9040 ) );
  nnd2s1 \IDinst/U9070  ( .DIN1(\IDinst/n9038 ), .DIN2(\IDinst/n9037 ), 
        .Q(\IDinst/n9039 ) );
  nnd2s1 \IDinst/U9069  ( .DIN1(\IDinst/n9036 ), .DIN2(n1322), 
        .Q(\IDinst/n9038 ) );
  nnd2s1 \IDinst/U9068  ( .DIN1(\IDinst/n9033 ), .DIN2(n1347), 
        .Q(\IDinst/n9037 ) );
  nnd2s1 \IDinst/U9067  ( .DIN1(\IDinst/n9035 ), .DIN2(\IDinst/n9034 ), 
        .Q(\IDinst/n9036 ) );
  nnd2s1 \IDinst/U9066  ( .DIN1(\IDinst/RegFile[31][0] ), .DIN2(n1227), 
        .Q(\IDinst/n9035 ) );
  nnd2s1 \IDinst/U9065  ( .DIN1(\IDinst/RegFile[30][0] ), .DIN2(n1255), 
        .Q(\IDinst/n9034 ) );
  nnd2s1 \IDinst/U9064  ( .DIN1(\IDinst/n9032 ), .DIN2(\IDinst/n9031 ), 
        .Q(\IDinst/n9033 ) );
  nnd2s1 \IDinst/U9063  ( .DIN1(\IDinst/RegFile[29][0] ), .DIN2(n1227), 
        .Q(\IDinst/n9032 ) );
  nnd2s1 \IDinst/U9062  ( .DIN1(\IDinst/RegFile[28][0] ), .DIN2(n1255), 
        .Q(\IDinst/n9031 ) );
  nnd2s1 \IDinst/U9061  ( .DIN1(\IDinst/n9029 ), .DIN2(\IDinst/n9028 ), 
        .Q(\IDinst/n9030 ) );
  nnd2s1 \IDinst/U9060  ( .DIN1(\IDinst/n9027 ), .DIN2(n1322), 
        .Q(\IDinst/n9029 ) );
  nnd2s1 \IDinst/U9059  ( .DIN1(\IDinst/n9024 ), .DIN2(n1347), 
        .Q(\IDinst/n9028 ) );
  nnd2s1 \IDinst/U9058  ( .DIN1(\IDinst/n9026 ), .DIN2(\IDinst/n9025 ), 
        .Q(\IDinst/n9027 ) );
  nnd2s1 \IDinst/U9057  ( .DIN1(\IDinst/RegFile[27][0] ), .DIN2(n1227), 
        .Q(\IDinst/n9026 ) );
  nnd2s1 \IDinst/U9056  ( .DIN1(\IDinst/RegFile[26][0] ), .DIN2(n1255), 
        .Q(\IDinst/n9025 ) );
  nnd2s1 \IDinst/U9055  ( .DIN1(\IDinst/n9023 ), .DIN2(\IDinst/n9022 ), 
        .Q(\IDinst/n9024 ) );
  nnd2s1 \IDinst/U9054  ( .DIN1(\IDinst/RegFile[25][0] ), .DIN2(n1227), 
        .Q(\IDinst/n9023 ) );
  nnd2s1 \IDinst/U9053  ( .DIN1(\IDinst/RegFile[24][0] ), .DIN2(n1255), 
        .Q(\IDinst/n9022 ) );
  nnd2s1 \IDinst/U9052  ( .DIN1(\IDinst/n9020 ), .DIN2(\IDinst/n9019 ), 
        .Q(\IDinst/n9021 ) );
  nnd2s1 \IDinst/U9051  ( .DIN1(\IDinst/n9018 ), .DIN2(n1380), 
        .Q(\IDinst/n9020 ) );
  nnd2s1 \IDinst/U9050  ( .DIN1(\IDinst/n9009 ), .DIN2(n1364), 
        .Q(\IDinst/n9019 ) );
  nnd2s1 \IDinst/U9049  ( .DIN1(\IDinst/n9017 ), .DIN2(\IDinst/n9016 ), 
        .Q(\IDinst/n9018 ) );
  nnd2s1 \IDinst/U9048  ( .DIN1(\IDinst/n9015 ), .DIN2(n1322), 
        .Q(\IDinst/n9017 ) );
  nnd2s1 \IDinst/U9047  ( .DIN1(\IDinst/n9012 ), .DIN2(n1347), 
        .Q(\IDinst/n9016 ) );
  nnd2s1 \IDinst/U9046  ( .DIN1(\IDinst/n9014 ), .DIN2(\IDinst/n9013 ), 
        .Q(\IDinst/n9015 ) );
  nnd2s1 \IDinst/U9045  ( .DIN1(\IDinst/RegFile[23][0] ), .DIN2(n1227), 
        .Q(\IDinst/n9014 ) );
  nnd2s1 \IDinst/U9044  ( .DIN1(\IDinst/RegFile[22][0] ), .DIN2(n1255), 
        .Q(\IDinst/n9013 ) );
  nnd2s1 \IDinst/U9043  ( .DIN1(\IDinst/n9011 ), .DIN2(\IDinst/n9010 ), 
        .Q(\IDinst/n9012 ) );
  nnd2s1 \IDinst/U9042  ( .DIN1(\IDinst/RegFile[21][0] ), .DIN2(n1227), 
        .Q(\IDinst/n9011 ) );
  nnd2s1 \IDinst/U9041  ( .DIN1(\IDinst/RegFile[20][0] ), .DIN2(n1255), 
        .Q(\IDinst/n9010 ) );
  nnd2s1 \IDinst/U9040  ( .DIN1(\IDinst/n9008 ), .DIN2(\IDinst/n9007 ), 
        .Q(\IDinst/n9009 ) );
  nnd2s1 \IDinst/U9039  ( .DIN1(\IDinst/n9006 ), .DIN2(n1322), 
        .Q(\IDinst/n9008 ) );
  nnd2s1 \IDinst/U9038  ( .DIN1(\IDinst/n9003 ), .DIN2(n1348), 
        .Q(\IDinst/n9007 ) );
  nnd2s1 \IDinst/U9037  ( .DIN1(\IDinst/n9005 ), .DIN2(\IDinst/n9004 ), 
        .Q(\IDinst/n9006 ) );
  nnd2s1 \IDinst/U9036  ( .DIN1(\IDinst/RegFile[19][0] ), .DIN2(n1227), 
        .Q(\IDinst/n9005 ) );
  nnd2s1 \IDinst/U9035  ( .DIN1(\IDinst/RegFile[18][0] ), .DIN2(n1255), 
        .Q(\IDinst/n9004 ) );
  nnd2s1 \IDinst/U9034  ( .DIN1(\IDinst/n9002 ), .DIN2(\IDinst/n9001 ), 
        .Q(\IDinst/n9003 ) );
  nnd2s1 \IDinst/U9033  ( .DIN1(\IDinst/RegFile[17][0] ), .DIN2(n1227), 
        .Q(\IDinst/n9002 ) );
  nnd2s1 \IDinst/U9032  ( .DIN1(\IDinst/RegFile[16][0] ), .DIN2(n1254), 
        .Q(\IDinst/n9001 ) );
  nnd2s1 \IDinst/U9031  ( .DIN1(\IDinst/n8999 ), .DIN2(\IDinst/n8998 ), 
        .Q(\IDinst/n9000 ) );
  nnd2s1 \IDinst/U9030  ( .DIN1(n667), .DIN2(\IDinst/n8997 ), 
        .Q(\IDinst/n8999 ) );
  nnd2s1 \IDinst/U9029  ( .DIN1(\IDinst/n8976 ), .DIN2(n681), 
        .Q(\IDinst/n8998 ) );
  nnd2s1 \IDinst/U9028  ( .DIN1(\IDinst/n8996 ), .DIN2(\IDinst/n8995 ), 
        .Q(\IDinst/n8997 ) );
  nnd2s1 \IDinst/U9027  ( .DIN1(\IDinst/n8994 ), .DIN2(\IDinst/N46 ), 
        .Q(\IDinst/n8996 ) );
  nnd2s1 \IDinst/U9026  ( .DIN1(\IDinst/n8985 ), .DIN2(n1364), 
        .Q(\IDinst/n8995 ) );
  nnd2s1 \IDinst/U9025  ( .DIN1(\IDinst/n8993 ), .DIN2(\IDinst/n8992 ), 
        .Q(\IDinst/n8994 ) );
  nnd2s1 \IDinst/U9024  ( .DIN1(\IDinst/n8991 ), .DIN2(n1322), 
        .Q(\IDinst/n8993 ) );
  nnd2s1 \IDinst/U9023  ( .DIN1(\IDinst/n8988 ), .DIN2(n1348), 
        .Q(\IDinst/n8992 ) );
  nnd2s1 \IDinst/U9022  ( .DIN1(\IDinst/n8990 ), .DIN2(\IDinst/n8989 ), 
        .Q(\IDinst/n8991 ) );
  nnd2s1 \IDinst/U9021  ( .DIN1(\IDinst/RegFile[15][0] ), .DIN2(n1227), 
        .Q(\IDinst/n8990 ) );
  nnd2s1 \IDinst/U9020  ( .DIN1(\IDinst/RegFile[14][0] ), .DIN2(n1254), 
        .Q(\IDinst/n8989 ) );
  nnd2s1 \IDinst/U9019  ( .DIN1(\IDinst/n8987 ), .DIN2(\IDinst/n8986 ), 
        .Q(\IDinst/n8988 ) );
  nnd2s1 \IDinst/U9018  ( .DIN1(\IDinst/RegFile[13][0] ), .DIN2(n1227), 
        .Q(\IDinst/n8987 ) );
  nnd2s1 \IDinst/U9017  ( .DIN1(\IDinst/RegFile[12][0] ), .DIN2(n1254), 
        .Q(\IDinst/n8986 ) );
  nnd2s1 \IDinst/U9016  ( .DIN1(\IDinst/n8984 ), .DIN2(\IDinst/n8983 ), 
        .Q(\IDinst/n8985 ) );
  nnd2s1 \IDinst/U9015  ( .DIN1(\IDinst/n8982 ), .DIN2(n1327), 
        .Q(\IDinst/n8984 ) );
  nnd2s1 \IDinst/U9014  ( .DIN1(\IDinst/n8979 ), .DIN2(n1348), 
        .Q(\IDinst/n8983 ) );
  nnd2s1 \IDinst/U9013  ( .DIN1(\IDinst/n8981 ), .DIN2(\IDinst/n8980 ), 
        .Q(\IDinst/n8982 ) );
  nnd2s1 \IDinst/U9012  ( .DIN1(\IDinst/RegFile[11][0] ), .DIN2(n1227), 
        .Q(\IDinst/n8981 ) );
  nnd2s1 \IDinst/U9011  ( .DIN1(\IDinst/RegFile[10][0] ), .DIN2(n1254), 
        .Q(\IDinst/n8980 ) );
  nnd2s1 \IDinst/U9010  ( .DIN1(\IDinst/n8978 ), .DIN2(\IDinst/n8977 ), 
        .Q(\IDinst/n8979 ) );
  nnd2s1 \IDinst/U9009  ( .DIN1(\IDinst/RegFile[9][0] ), .DIN2(n1227), 
        .Q(\IDinst/n8978 ) );
  nnd2s1 \IDinst/U9008  ( .DIN1(\IDinst/RegFile[8][0] ), .DIN2(n1254), 
        .Q(\IDinst/n8977 ) );
  nnd2s1 \IDinst/U9007  ( .DIN1(\IDinst/n8975 ), .DIN2(\IDinst/n8974 ), 
        .Q(\IDinst/n8976 ) );
  nnd2s1 \IDinst/U9006  ( .DIN1(n1372), .DIN2(\IDinst/n8973 ), 
        .Q(\IDinst/n8975 ) );
  nnd2s1 \IDinst/U9005  ( .DIN1(\IDinst/n8964 ), .DIN2(n1368), 
        .Q(\IDinst/n8974 ) );
  nnd2s1 \IDinst/U9004  ( .DIN1(\IDinst/n8972 ), .DIN2(\IDinst/n8971 ), 
        .Q(\IDinst/n8973 ) );
  nnd2s1 \IDinst/U9003  ( .DIN1(\IDinst/n8970 ), .DIN2(n1312), 
        .Q(\IDinst/n8972 ) );
  nnd2s1 \IDinst/U9002  ( .DIN1(\IDinst/n8967 ), .DIN2(n1333), 
        .Q(\IDinst/n8971 ) );
  nnd2s1 \IDinst/U9001  ( .DIN1(\IDinst/n8969 ), .DIN2(\IDinst/n8968 ), 
        .Q(\IDinst/n8970 ) );
  nnd2s1 \IDinst/U9000  ( .DIN1(\IDinst/RegFile[7][0] ), .DIN2(n1228), 
        .Q(\IDinst/n8969 ) );
  nnd2s1 \IDinst/U8999  ( .DIN1(\IDinst/RegFile[6][0] ), .DIN2(n1254), 
        .Q(\IDinst/n8968 ) );
  nnd2s1 \IDinst/U8998  ( .DIN1(\IDinst/n8966 ), .DIN2(\IDinst/n8965 ), 
        .Q(\IDinst/n8967 ) );
  nnd2s1 \IDinst/U8997  ( .DIN1(\IDinst/RegFile[5][0] ), .DIN2(n1228), 
        .Q(\IDinst/n8966 ) );
  nnd2s1 \IDinst/U8996  ( .DIN1(\IDinst/RegFile[4][0] ), .DIN2(n1261), 
        .Q(\IDinst/n8965 ) );
  nnd2s1 \IDinst/U8995  ( .DIN1(\IDinst/n8963 ), .DIN2(\IDinst/n8962 ), 
        .Q(\IDinst/n8964 ) );
  nnd2s1 \IDinst/U8994  ( .DIN1(n1312), .DIN2(\IDinst/n8961 ), 
        .Q(\IDinst/n8963 ) );
  nnd2s1 \IDinst/U8993  ( .DIN1(\IDinst/n8958 ), .DIN2(n1353), 
        .Q(\IDinst/n8962 ) );
  nnd2s1 \IDinst/U8992  ( .DIN1(\IDinst/n8960 ), .DIN2(\IDinst/n8959 ), 
        .Q(\IDinst/n8961 ) );
  nnd2s1 \IDinst/U8991  ( .DIN1(\IDinst/RegFile[3][0] ), .DIN2(n1228), 
        .Q(\IDinst/n8960 ) );
  nnd2s1 \IDinst/U8990  ( .DIN1(\IDinst/RegFile[2][0] ), .DIN2(n1239), 
        .Q(\IDinst/n8959 ) );
  nnd2s1 \IDinst/U8989  ( .DIN1(\IDinst/n8957 ), .DIN2(\IDinst/n8956 ), 
        .Q(\IDinst/n8958 ) );
  nnd2s1 \IDinst/U8988  ( .DIN1(\IDinst/RegFile[1][0] ), .DIN2(n1198), 
        .Q(\IDinst/n8957 ) );
  nnd2s1 \IDinst/U8987  ( .DIN1(\IDinst/RegFile[0][0] ), .DIN2(n1292), 
        .Q(\IDinst/n8956 ) );
  nnd2s1 \IDinst/U8986  ( .DIN1(\IDinst/n8954 ), .DIN2(\IDinst/n8955 ), 
        .Q(\IDinst/N89 ) );
  nnd2s1 \IDinst/U8985  ( .DIN1(\IDinst/n8952 ), .DIN2(\IDinst/n8953 ), 
        .Q(\IDinst/N90 ) );
  nnd2s1 \IDinst/U8984  ( .DIN1(\IDinst/n8950 ), .DIN2(\IDinst/n8951 ), 
        .Q(\IDinst/N91 ) );
  nnd2s1 \IDinst/U8983  ( .DIN1(\IDinst/n8948 ), .DIN2(\IDinst/n8949 ), 
        .Q(\IDinst/N92 ) );
  nnd2s1 \IDinst/U8982  ( .DIN1(\IDinst/n8946 ), .DIN2(\IDinst/n8947 ), 
        .Q(\IDinst/N93 ) );
  nnd2s1 \IDinst/U8981  ( .DIN1(\IDinst/n8944 ), .DIN2(\IDinst/n8945 ), 
        .Q(\IDinst/N94 ) );
  nnd2s1 \IDinst/U8980  ( .DIN1(\IDinst/n8942 ), .DIN2(\IDinst/n8943 ), 
        .Q(\IDinst/N95 ) );
  nnd2s1 \IDinst/U8979  ( .DIN1(\IDinst/n8940 ), .DIN2(\IDinst/n8941 ), 
        .Q(\IDinst/N96 ) );
  nnd2s1 \IDinst/U8978  ( .DIN1(\IDinst/n8938 ), .DIN2(\IDinst/n8939 ), 
        .Q(\IDinst/N97 ) );
  nnd2s1 \IDinst/U8977  ( .DIN1(\IDinst/n8936 ), .DIN2(\IDinst/n8937 ), 
        .Q(\IDinst/N98 ) );
  nnd2s1 \IDinst/U8976  ( .DIN1(\IDinst/n8934 ), .DIN2(\IDinst/n8935 ), 
        .Q(\IDinst/N99 ) );
  nnd2s1 \IDinst/U8975  ( .DIN1(\IDinst/n8932 ), .DIN2(\IDinst/n8933 ), 
        .Q(\IDinst/N100 ) );
  nnd2s1 \IDinst/U8974  ( .DIN1(\IDinst/n8930 ), .DIN2(\IDinst/n8931 ), 
        .Q(\IDinst/N101 ) );
  nnd2s1 \IDinst/U8973  ( .DIN1(\IDinst/n8928 ), .DIN2(\IDinst/n8929 ), 
        .Q(\IDinst/N102 ) );
  nnd2s1 \IDinst/U8972  ( .DIN1(\IDinst/n8926 ), .DIN2(\IDinst/n8927 ), 
        .Q(\IDinst/N103 ) );
  nnd2s1 \IDinst/U8971  ( .DIN1(\IDinst/n8924 ), .DIN2(\IDinst/n8925 ), 
        .Q(\IDinst/N104 ) );
  nnd2s1 \IDinst/U8970  ( .DIN1(\IDinst/n8922 ), .DIN2(\IDinst/n8923 ), 
        .Q(\IDinst/N105 ) );
  nnd2s1 \IDinst/U8969  ( .DIN1(\IDinst/n8920 ), .DIN2(\IDinst/n8921 ), 
        .Q(\IDinst/N106 ) );
  nnd2s1 \IDinst/U8968  ( .DIN1(\IDinst/n8918 ), .DIN2(\IDinst/n8919 ), 
        .Q(\IDinst/N107 ) );
  nnd2s1 \IDinst/U8967  ( .DIN1(\IDinst/n8916 ), .DIN2(\IDinst/n8917 ), 
        .Q(\IDinst/N108 ) );
  nnd2s1 \IDinst/U8966  ( .DIN1(\IDinst/n8914 ), .DIN2(\IDinst/n8915 ), 
        .Q(\IDinst/N109 ) );
  nnd2s1 \IDinst/U8965  ( .DIN1(\IDinst/n8912 ), .DIN2(\IDinst/n8913 ), 
        .Q(\IDinst/N110 ) );
  nnd2s1 \IDinst/U8964  ( .DIN1(\IDinst/n8910 ), .DIN2(\IDinst/n8911 ), 
        .Q(\IDinst/N111 ) );
  nnd2s1 \IDinst/U8963  ( .DIN1(\IDinst/n8908 ), .DIN2(\IDinst/n8909 ), 
        .Q(\IDinst/N112 ) );
  nnd2s1 \IDinst/U8962  ( .DIN1(\IDinst/n8906 ), .DIN2(\IDinst/n8907 ), 
        .Q(\IDinst/N113 ) );
  nnd2s1 \IDinst/U8961  ( .DIN1(\IDinst/n8904 ), .DIN2(\IDinst/n8905 ), 
        .Q(\IDinst/N114 ) );
  nnd2s1 \IDinst/U8960  ( .DIN1(\IDinst/n8902 ), .DIN2(\IDinst/n8903 ), 
        .Q(\IDinst/N115 ) );
  nnd2s1 \IDinst/U8959  ( .DIN1(\IDinst/n8900 ), .DIN2(\IDinst/n8901 ), 
        .Q(\IDinst/N116 ) );
  nnd2s1 \IDinst/U8958  ( .DIN1(\IDinst/n8898 ), .DIN2(\IDinst/n8899 ), 
        .Q(\IDinst/N117 ) );
  nnd2s1 \IDinst/U8957  ( .DIN1(\IDinst/n8896 ), .DIN2(\IDinst/n8897 ), 
        .Q(\IDinst/N118 ) );
  nnd2s1 \IDinst/U8956  ( .DIN1(\IDinst/n8894 ), .DIN2(\IDinst/n8895 ), 
        .Q(\IDinst/N119 ) );
  nnd2s1 \IDinst/U8955  ( .DIN1(\IDinst/n8892 ), .DIN2(\IDinst/n8893 ), 
        .Q(\IDinst/N120 ) );
  nnd2s1 \IDinst/U8954  ( .DIN1(\IDinst/n8891 ), .DIN2(n539), 
        .Q(\IDinst/n6010 ) );
  nnd2s1 \IDinst/U8953  ( .DIN1(\IDinst/n8846 ), .DIN2(n635), 
        .Q(\IDinst/n6011 ) );
  nnd2s1 \IDinst/U8952  ( .DIN1(\IDinst/n8890 ), .DIN2(\IDinst/n8889 ), 
        .Q(\IDinst/n8891 ) );
  nnd2s1 \IDinst/U8951  ( .DIN1(\IDinst/n8888 ), .DIN2(n643), 
        .Q(\IDinst/n8890 ) );
  nnd2s1 \IDinst/U8950  ( .DIN1(\IDinst/n8867 ), .DIN2(n673), 
        .Q(\IDinst/n8889 ) );
  nnd2s1 \IDinst/U8949  ( .DIN1(\IDinst/n8887 ), .DIN2(\IDinst/n8886 ), 
        .Q(\IDinst/n8888 ) );
  nnd2s1 \IDinst/U8948  ( .DIN1(\IDinst/n8885 ), .DIN2(n1191), 
        .Q(\IDinst/n8887 ) );
  nnd2s1 \IDinst/U8947  ( .DIN1(\IDinst/n8876 ), .DIN2(n1189), 
        .Q(\IDinst/n8886 ) );
  nnd2s1 \IDinst/U8946  ( .DIN1(\IDinst/n8884 ), .DIN2(\IDinst/n8883 ), 
        .Q(\IDinst/n8885 ) );
  nnd2s1 \IDinst/U8945  ( .DIN1(\IDinst/n8882 ), .DIN2(\IDinst/N40 ), 
        .Q(\IDinst/n8884 ) );
  nnd2s1 \IDinst/U8944  ( .DIN1(\IDinst/n8879 ), .DIN2(n1143), 
        .Q(\IDinst/n8883 ) );
  nnd2s1 \IDinst/U8943  ( .DIN1(\IDinst/n8881 ), .DIN2(\IDinst/n8880 ), 
        .Q(\IDinst/n8882 ) );
  nnd2s1 \IDinst/U8942  ( .DIN1(\IDinst/RegFile[31][31] ), .DIN2(n1119), 
        .Q(\IDinst/n8881 ) );
  nnd2s1 \IDinst/U8941  ( .DIN1(\IDinst/RegFile[30][31] ), .DIN2(n1055), 
        .Q(\IDinst/n8880 ) );
  nnd2s1 \IDinst/U8940  ( .DIN1(\IDinst/n8878 ), .DIN2(\IDinst/n8877 ), 
        .Q(\IDinst/n8879 ) );
  nnd2s1 \IDinst/U8939  ( .DIN1(\IDinst/RegFile[29][31] ), .DIN2(n1065), 
        .Q(\IDinst/n8878 ) );
  nnd2s1 \IDinst/U8938  ( .DIN1(\IDinst/RegFile[28][31] ), .DIN2(n1055), 
        .Q(\IDinst/n8877 ) );
  nnd2s1 \IDinst/U8937  ( .DIN1(\IDinst/n8875 ), .DIN2(\IDinst/n8874 ), 
        .Q(\IDinst/n8876 ) );
  nnd2s1 \IDinst/U8936  ( .DIN1(\IDinst/n8873 ), .DIN2(n1155), 
        .Q(\IDinst/n8875 ) );
  nnd2s1 \IDinst/U8935  ( .DIN1(\IDinst/n8870 ), .DIN2(n1143), 
        .Q(\IDinst/n8874 ) );
  nnd2s1 \IDinst/U8934  ( .DIN1(\IDinst/n8872 ), .DIN2(\IDinst/n8871 ), 
        .Q(\IDinst/n8873 ) );
  nnd2s1 \IDinst/U8933  ( .DIN1(\IDinst/RegFile[27][31] ), .DIN2(n1088), 
        .Q(\IDinst/n8872 ) );
  nnd2s1 \IDinst/U8932  ( .DIN1(\IDinst/RegFile[26][31] ), .DIN2(n1055), 
        .Q(\IDinst/n8871 ) );
  nnd2s1 \IDinst/U8931  ( .DIN1(\IDinst/n8869 ), .DIN2(\IDinst/n8868 ), 
        .Q(\IDinst/n8870 ) );
  nnd2s1 \IDinst/U8930  ( .DIN1(\IDinst/RegFile[25][31] ), .DIN2(n1081), 
        .Q(\IDinst/n8869 ) );
  nnd2s1 \IDinst/U8929  ( .DIN1(\IDinst/RegFile[24][31] ), .DIN2(n1054), 
        .Q(\IDinst/n8868 ) );
  nnd2s1 \IDinst/U8928  ( .DIN1(\IDinst/n8866 ), .DIN2(\IDinst/n8865 ), 
        .Q(\IDinst/n8867 ) );
  nnd2s1 \IDinst/U8927  ( .DIN1(\IDinst/n8864 ), .DIN2(n1193), 
        .Q(\IDinst/n8866 ) );
  nnd2s1 \IDinst/U8926  ( .DIN1(\IDinst/n8855 ), .DIN2(n1188), 
        .Q(\IDinst/n8865 ) );
  nnd2s1 \IDinst/U8925  ( .DIN1(\IDinst/n8863 ), .DIN2(\IDinst/n8862 ), 
        .Q(\IDinst/n8864 ) );
  nnd2s1 \IDinst/U8924  ( .DIN1(\IDinst/n8861 ), .DIN2(n1166), 
        .Q(\IDinst/n8863 ) );
  nnd2s1 \IDinst/U8923  ( .DIN1(\IDinst/n8858 ), .DIN2(n1143), 
        .Q(\IDinst/n8862 ) );
  nnd2s1 \IDinst/U8922  ( .DIN1(\IDinst/n8860 ), .DIN2(\IDinst/n8859 ), 
        .Q(\IDinst/n8861 ) );
  nnd2s1 \IDinst/U8921  ( .DIN1(\IDinst/RegFile[23][31] ), .DIN2(n1081), 
        .Q(\IDinst/n8860 ) );
  nnd2s1 \IDinst/U8920  ( .DIN1(\IDinst/RegFile[22][31] ), .DIN2(n1054), 
        .Q(\IDinst/n8859 ) );
  nnd2s1 \IDinst/U8919  ( .DIN1(\IDinst/n8857 ), .DIN2(\IDinst/n8856 ), 
        .Q(\IDinst/n8858 ) );
  nnd2s1 \IDinst/U8918  ( .DIN1(\IDinst/RegFile[21][31] ), .DIN2(n1081), 
        .Q(\IDinst/n8857 ) );
  nnd2s1 \IDinst/U8917  ( .DIN1(\IDinst/RegFile[20][31] ), .DIN2(n1054), 
        .Q(\IDinst/n8856 ) );
  nnd2s1 \IDinst/U8916  ( .DIN1(\IDinst/n8854 ), .DIN2(\IDinst/n8853 ), 
        .Q(\IDinst/n8855 ) );
  nnd2s1 \IDinst/U8915  ( .DIN1(\IDinst/n8852 ), .DIN2(n1166), 
        .Q(\IDinst/n8854 ) );
  nnd2s1 \IDinst/U8914  ( .DIN1(\IDinst/n8849 ), .DIN2(n1143), 
        .Q(\IDinst/n8853 ) );
  nnd2s1 \IDinst/U8913  ( .DIN1(\IDinst/n8851 ), .DIN2(\IDinst/n8850 ), 
        .Q(\IDinst/n8852 ) );
  nnd2s1 \IDinst/U8912  ( .DIN1(\IDinst/RegFile[19][31] ), .DIN2(n1081), 
        .Q(\IDinst/n8851 ) );
  nnd2s1 \IDinst/U8911  ( .DIN1(\IDinst/RegFile[18][31] ), .DIN2(n1054), 
        .Q(\IDinst/n8850 ) );
  nnd2s1 \IDinst/U8910  ( .DIN1(\IDinst/n8848 ), .DIN2(\IDinst/n8847 ), 
        .Q(\IDinst/n8849 ) );
  nnd2s1 \IDinst/U8909  ( .DIN1(\IDinst/RegFile[17][31] ), .DIN2(n1081), 
        .Q(\IDinst/n8848 ) );
  nnd2s1 \IDinst/U8908  ( .DIN1(\IDinst/RegFile[16][31] ), .DIN2(n1054), 
        .Q(\IDinst/n8847 ) );
  nnd2s1 \IDinst/U8907  ( .DIN1(\IDinst/n8845 ), .DIN2(\IDinst/n8844 ), 
        .Q(\IDinst/n8846 ) );
  nnd2s1 \IDinst/U8906  ( .DIN1(\IDinst/n8843 ), .DIN2(n642), 
        .Q(\IDinst/n8845 ) );
  nnd2s1 \IDinst/U8905  ( .DIN1(\IDinst/n8822 ), .DIN2(n670), 
        .Q(\IDinst/n8844 ) );
  nnd2s1 \IDinst/U8904  ( .DIN1(\IDinst/n8842 ), .DIN2(\IDinst/n8841 ), 
        .Q(\IDinst/n8843 ) );
  nnd2s1 \IDinst/U8903  ( .DIN1(\IDinst/n8840 ), .DIN2(n1190), 
        .Q(\IDinst/n8842 ) );
  nnd2s1 \IDinst/U8902  ( .DIN1(\IDinst/n8831 ), .DIN2(n1187), 
        .Q(\IDinst/n8841 ) );
  nnd2s1 \IDinst/U8901  ( .DIN1(\IDinst/n8839 ), .DIN2(\IDinst/n8838 ), 
        .Q(\IDinst/n8840 ) );
  nnd2s1 \IDinst/U8900  ( .DIN1(\IDinst/n8837 ), .DIN2(n1156), 
        .Q(\IDinst/n8839 ) );
  nnd2s1 \IDinst/U8899  ( .DIN1(\IDinst/n8834 ), .DIN2(n1143), 
        .Q(\IDinst/n8838 ) );
  nnd2s1 \IDinst/U8898  ( .DIN1(\IDinst/n8836 ), .DIN2(\IDinst/n8835 ), 
        .Q(\IDinst/n8837 ) );
  nnd2s1 \IDinst/U8897  ( .DIN1(\IDinst/RegFile[15][31] ), .DIN2(n1081), 
        .Q(\IDinst/n8836 ) );
  nnd2s1 \IDinst/U8896  ( .DIN1(\IDinst/RegFile[14][31] ), .DIN2(n1054), 
        .Q(\IDinst/n8835 ) );
  nnd2s1 \IDinst/U8895  ( .DIN1(\IDinst/n8833 ), .DIN2(\IDinst/n8832 ), 
        .Q(\IDinst/n8834 ) );
  nnd2s1 \IDinst/U8894  ( .DIN1(\IDinst/RegFile[13][31] ), .DIN2(n1081), 
        .Q(\IDinst/n8833 ) );
  nnd2s1 \IDinst/U8893  ( .DIN1(\IDinst/RegFile[12][31] ), .DIN2(n1054), 
        .Q(\IDinst/n8832 ) );
  nnd2s1 \IDinst/U8892  ( .DIN1(\IDinst/n8830 ), .DIN2(\IDinst/n8829 ), 
        .Q(\IDinst/n8831 ) );
  nnd2s1 \IDinst/U8891  ( .DIN1(\IDinst/n8828 ), .DIN2(n1161), 
        .Q(\IDinst/n8830 ) );
  nnd2s1 \IDinst/U8890  ( .DIN1(\IDinst/n8825 ), .DIN2(n1144), 
        .Q(\IDinst/n8829 ) );
  nnd2s1 \IDinst/U8889  ( .DIN1(\IDinst/n8827 ), .DIN2(\IDinst/n8826 ), 
        .Q(\IDinst/n8828 ) );
  nnd2s1 \IDinst/U8888  ( .DIN1(\IDinst/RegFile[11][31] ), .DIN2(n1082), 
        .Q(\IDinst/n8827 ) );
  nnd2s1 \IDinst/U8887  ( .DIN1(\IDinst/RegFile[10][31] ), .DIN2(n1054), 
        .Q(\IDinst/n8826 ) );
  nnd2s1 \IDinst/U8886  ( .DIN1(\IDinst/n8824 ), .DIN2(\IDinst/n8823 ), 
        .Q(\IDinst/n8825 ) );
  nnd2s1 \IDinst/U8885  ( .DIN1(\IDinst/RegFile[9][31] ), .DIN2(n1082), 
        .Q(\IDinst/n8824 ) );
  nnd2s1 \IDinst/U8884  ( .DIN1(\IDinst/RegFile[8][31] ), .DIN2(n1054), 
        .Q(\IDinst/n8823 ) );
  nnd2s1 \IDinst/U8883  ( .DIN1(\IDinst/n8821 ), .DIN2(\IDinst/n8820 ), 
        .Q(\IDinst/n8822 ) );
  nnd2s1 \IDinst/U8882  ( .DIN1(\IDinst/n8819 ), .DIN2(n1195), 
        .Q(\IDinst/n8821 ) );
  nnd2s1 \IDinst/U8881  ( .DIN1(\IDinst/n8810 ), .DIN2(n1186), 
        .Q(\IDinst/n8820 ) );
  nnd2s1 \IDinst/U8880  ( .DIN1(\IDinst/n8818 ), .DIN2(\IDinst/n8817 ), 
        .Q(\IDinst/n8819 ) );
  nnd2s1 \IDinst/U8879  ( .DIN1(\IDinst/n8816 ), .DIN2(n1171), 
        .Q(\IDinst/n8818 ) );
  nnd2s1 \IDinst/U8878  ( .DIN1(\IDinst/n8813 ), .DIN2(n1144), 
        .Q(\IDinst/n8817 ) );
  nnd2s1 \IDinst/U8877  ( .DIN1(\IDinst/n8815 ), .DIN2(\IDinst/n8814 ), 
        .Q(\IDinst/n8816 ) );
  nnd2s1 \IDinst/U8876  ( .DIN1(\IDinst/RegFile[7][31] ), .DIN2(n1082), 
        .Q(\IDinst/n8815 ) );
  nnd2s1 \IDinst/U8875  ( .DIN1(\IDinst/RegFile[6][31] ), .DIN2(n1054), 
        .Q(\IDinst/n8814 ) );
  nnd2s1 \IDinst/U8874  ( .DIN1(\IDinst/n8812 ), .DIN2(\IDinst/n8811 ), 
        .Q(\IDinst/n8813 ) );
  nnd2s1 \IDinst/U8873  ( .DIN1(\IDinst/RegFile[5][31] ), .DIN2(n1082), 
        .Q(\IDinst/n8812 ) );
  nnd2s1 \IDinst/U8872  ( .DIN1(\IDinst/RegFile[4][31] ), .DIN2(n1054), 
        .Q(\IDinst/n8811 ) );
  nnd2s1 \IDinst/U8871  ( .DIN1(\IDinst/n8809 ), .DIN2(\IDinst/n8808 ), 
        .Q(\IDinst/n8810 ) );
  nnd2s1 \IDinst/U8870  ( .DIN1(\IDinst/n8807 ), .DIN2(n1169), 
        .Q(\IDinst/n8809 ) );
  nnd2s1 \IDinst/U8869  ( .DIN1(\IDinst/n8804 ), .DIN2(n1144), 
        .Q(\IDinst/n8808 ) );
  nnd2s1 \IDinst/U8868  ( .DIN1(\IDinst/n8806 ), .DIN2(\IDinst/n8805 ), 
        .Q(\IDinst/n8807 ) );
  nnd2s1 \IDinst/U8867  ( .DIN1(\IDinst/RegFile[3][31] ), .DIN2(n1082), 
        .Q(\IDinst/n8806 ) );
  nnd2s1 \IDinst/U8866  ( .DIN1(\IDinst/RegFile[2][31] ), .DIN2(n1054), 
        .Q(\IDinst/n8805 ) );
  nnd2s1 \IDinst/U8865  ( .DIN1(\IDinst/n8803 ), .DIN2(\IDinst/n8802 ), 
        .Q(\IDinst/n8804 ) );
  nnd2s1 \IDinst/U8864  ( .DIN1(\IDinst/RegFile[1][31] ), .DIN2(n1082), 
        .Q(\IDinst/n8803 ) );
  nnd2s1 \IDinst/U8863  ( .DIN1(\IDinst/RegFile[0][31] ), .DIN2(n1054), 
        .Q(\IDinst/n8802 ) );
  nnd2s1 \IDinst/U8862  ( .DIN1(\IDinst/n8801 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n6008 ) );
  nnd2s1 \IDinst/U8861  ( .DIN1(\IDinst/n8756 ), .DIN2(n636), 
        .Q(\IDinst/n6009 ) );
  nnd2s1 \IDinst/U8860  ( .DIN1(\IDinst/n8800 ), .DIN2(\IDinst/n8799 ), 
        .Q(\IDinst/n8801 ) );
  nnd2s1 \IDinst/U8859  ( .DIN1(\IDinst/n8798 ), .DIN2(n641), 
        .Q(\IDinst/n8800 ) );
  nnd2s1 \IDinst/U8858  ( .DIN1(\IDinst/n8777 ), .DIN2(n673), 
        .Q(\IDinst/n8799 ) );
  nnd2s1 \IDinst/U8857  ( .DIN1(\IDinst/n8797 ), .DIN2(\IDinst/n8796 ), 
        .Q(\IDinst/n8798 ) );
  nnd2s1 \IDinst/U8856  ( .DIN1(\IDinst/n8795 ), .DIN2(n1192), 
        .Q(\IDinst/n8797 ) );
  nnd2s1 \IDinst/U8855  ( .DIN1(\IDinst/n8786 ), .DIN2(n1185), 
        .Q(\IDinst/n8796 ) );
  nnd2s1 \IDinst/U8854  ( .DIN1(\IDinst/n8794 ), .DIN2(\IDinst/n8793 ), 
        .Q(\IDinst/n8795 ) );
  nnd2s1 \IDinst/U8853  ( .DIN1(\IDinst/n8792 ), .DIN2(n1174), 
        .Q(\IDinst/n8794 ) );
  nnd2s1 \IDinst/U8852  ( .DIN1(\IDinst/n8789 ), .DIN2(n1144), 
        .Q(\IDinst/n8793 ) );
  nnd2s1 \IDinst/U8851  ( .DIN1(\IDinst/n8791 ), .DIN2(\IDinst/n8790 ), 
        .Q(\IDinst/n8792 ) );
  nnd2s1 \IDinst/U8850  ( .DIN1(\IDinst/RegFile[31][30] ), .DIN2(n1082), 
        .Q(\IDinst/n8791 ) );
  nnd2s1 \IDinst/U8849  ( .DIN1(\IDinst/RegFile[30][30] ), .DIN2(n1053), 
        .Q(\IDinst/n8790 ) );
  nnd2s1 \IDinst/U8848  ( .DIN1(\IDinst/n8788 ), .DIN2(\IDinst/n8787 ), 
        .Q(\IDinst/n8789 ) );
  nnd2s1 \IDinst/U8847  ( .DIN1(\IDinst/RegFile[29][30] ), .DIN2(n1082), 
        .Q(\IDinst/n8788 ) );
  nnd2s1 \IDinst/U8846  ( .DIN1(\IDinst/RegFile[28][30] ), .DIN2(n1053), 
        .Q(\IDinst/n8787 ) );
  nnd2s1 \IDinst/U8845  ( .DIN1(\IDinst/n8785 ), .DIN2(\IDinst/n8784 ), 
        .Q(\IDinst/n8786 ) );
  nnd2s1 \IDinst/U8844  ( .DIN1(\IDinst/n8783 ), .DIN2(n1162), 
        .Q(\IDinst/n8785 ) );
  nnd2s1 \IDinst/U8843  ( .DIN1(\IDinst/n8780 ), .DIN2(n1144), 
        .Q(\IDinst/n8784 ) );
  nnd2s1 \IDinst/U8842  ( .DIN1(\IDinst/n8782 ), .DIN2(\IDinst/n8781 ), 
        .Q(\IDinst/n8783 ) );
  nnd2s1 \IDinst/U8841  ( .DIN1(\IDinst/RegFile[27][30] ), .DIN2(n1082), 
        .Q(\IDinst/n8782 ) );
  nnd2s1 \IDinst/U8840  ( .DIN1(\IDinst/RegFile[26][30] ), .DIN2(n1053), 
        .Q(\IDinst/n8781 ) );
  nnd2s1 \IDinst/U8839  ( .DIN1(\IDinst/n8779 ), .DIN2(\IDinst/n8778 ), 
        .Q(\IDinst/n8780 ) );
  nnd2s1 \IDinst/U8838  ( .DIN1(\IDinst/RegFile[25][30] ), .DIN2(n1083), 
        .Q(\IDinst/n8779 ) );
  nnd2s1 \IDinst/U8837  ( .DIN1(\IDinst/RegFile[24][30] ), .DIN2(n1053), 
        .Q(\IDinst/n8778 ) );
  nnd2s1 \IDinst/U8836  ( .DIN1(\IDinst/n8776 ), .DIN2(\IDinst/n8775 ), 
        .Q(\IDinst/n8777 ) );
  nnd2s1 \IDinst/U8835  ( .DIN1(\IDinst/n8774 ), .DIN2(n1191), 
        .Q(\IDinst/n8776 ) );
  nnd2s1 \IDinst/U8834  ( .DIN1(\IDinst/n8765 ), .DIN2(n1184), 
        .Q(\IDinst/n8775 ) );
  nnd2s1 \IDinst/U8833  ( .DIN1(\IDinst/n8773 ), .DIN2(\IDinst/n8772 ), 
        .Q(\IDinst/n8774 ) );
  nnd2s1 \IDinst/U8832  ( .DIN1(\IDinst/n8771 ), .DIN2(n1167), 
        .Q(\IDinst/n8773 ) );
  nnd2s1 \IDinst/U8831  ( .DIN1(\IDinst/n8768 ), .DIN2(n1144), 
        .Q(\IDinst/n8772 ) );
  nnd2s1 \IDinst/U8830  ( .DIN1(\IDinst/n8770 ), .DIN2(\IDinst/n8769 ), 
        .Q(\IDinst/n8771 ) );
  nnd2s1 \IDinst/U8829  ( .DIN1(\IDinst/RegFile[23][30] ), .DIN2(n1083), 
        .Q(\IDinst/n8770 ) );
  nnd2s1 \IDinst/U8828  ( .DIN1(\IDinst/RegFile[22][30] ), .DIN2(n1053), 
        .Q(\IDinst/n8769 ) );
  nnd2s1 \IDinst/U8827  ( .DIN1(\IDinst/n8767 ), .DIN2(\IDinst/n8766 ), 
        .Q(\IDinst/n8768 ) );
  nnd2s1 \IDinst/U8826  ( .DIN1(\IDinst/RegFile[21][30] ), .DIN2(n1083), 
        .Q(\IDinst/n8767 ) );
  nnd2s1 \IDinst/U8825  ( .DIN1(\IDinst/RegFile[20][30] ), .DIN2(n1053), 
        .Q(\IDinst/n8766 ) );
  nnd2s1 \IDinst/U8824  ( .DIN1(\IDinst/n8764 ), .DIN2(\IDinst/n8763 ), 
        .Q(\IDinst/n8765 ) );
  nnd2s1 \IDinst/U8823  ( .DIN1(\IDinst/n8762 ), .DIN2(n1172), 
        .Q(\IDinst/n8764 ) );
  nnd2s1 \IDinst/U8822  ( .DIN1(\IDinst/n8759 ), .DIN2(n1144), 
        .Q(\IDinst/n8763 ) );
  nnd2s1 \IDinst/U8821  ( .DIN1(\IDinst/n8761 ), .DIN2(\IDinst/n8760 ), 
        .Q(\IDinst/n8762 ) );
  nnd2s1 \IDinst/U8820  ( .DIN1(\IDinst/RegFile[19][30] ), .DIN2(n1083), 
        .Q(\IDinst/n8761 ) );
  nnd2s1 \IDinst/U8819  ( .DIN1(\IDinst/RegFile[18][30] ), .DIN2(n1053), 
        .Q(\IDinst/n8760 ) );
  nnd2s1 \IDinst/U8818  ( .DIN1(\IDinst/n8758 ), .DIN2(\IDinst/n8757 ), 
        .Q(\IDinst/n8759 ) );
  nnd2s1 \IDinst/U8817  ( .DIN1(\IDinst/RegFile[17][30] ), .DIN2(n1083), 
        .Q(\IDinst/n8758 ) );
  nnd2s1 \IDinst/U8816  ( .DIN1(\IDinst/RegFile[16][30] ), .DIN2(n1053), 
        .Q(\IDinst/n8757 ) );
  nnd2s1 \IDinst/U8815  ( .DIN1(\IDinst/n8755 ), .DIN2(\IDinst/n8754 ), 
        .Q(\IDinst/n8756 ) );
  nnd2s1 \IDinst/U8814  ( .DIN1(\IDinst/n8753 ), .DIN2(n644), 
        .Q(\IDinst/n8755 ) );
  nnd2s1 \IDinst/U8813  ( .DIN1(\IDinst/n8732 ), .DIN2(n670), 
        .Q(\IDinst/n8754 ) );
  nnd2s1 \IDinst/U8812  ( .DIN1(\IDinst/n8752 ), .DIN2(\IDinst/n8751 ), 
        .Q(\IDinst/n8753 ) );
  nnd2s1 \IDinst/U8811  ( .DIN1(\IDinst/n8750 ), .DIN2(\IDinst/N41 ), 
        .Q(\IDinst/n8752 ) );
  nnd2s1 \IDinst/U8810  ( .DIN1(\IDinst/n8741 ), .DIN2(n1189), 
        .Q(\IDinst/n8751 ) );
  nnd2s1 \IDinst/U8809  ( .DIN1(\IDinst/n8749 ), .DIN2(\IDinst/n8748 ), 
        .Q(\IDinst/n8750 ) );
  nnd2s1 \IDinst/U8808  ( .DIN1(\IDinst/n8747 ), .DIN2(n1160), 
        .Q(\IDinst/n8749 ) );
  nnd2s1 \IDinst/U8807  ( .DIN1(\IDinst/n8744 ), .DIN2(n1144), 
        .Q(\IDinst/n8748 ) );
  nnd2s1 \IDinst/U8806  ( .DIN1(\IDinst/n8746 ), .DIN2(\IDinst/n8745 ), 
        .Q(\IDinst/n8747 ) );
  nnd2s1 \IDinst/U8805  ( .DIN1(\IDinst/RegFile[15][30] ), .DIN2(n1083), 
        .Q(\IDinst/n8746 ) );
  nnd2s1 \IDinst/U8804  ( .DIN1(\IDinst/RegFile[14][30] ), .DIN2(n1053), 
        .Q(\IDinst/n8745 ) );
  nnd2s1 \IDinst/U8803  ( .DIN1(\IDinst/n8743 ), .DIN2(\IDinst/n8742 ), 
        .Q(\IDinst/n8744 ) );
  nnd2s1 \IDinst/U8802  ( .DIN1(\IDinst/RegFile[13][30] ), .DIN2(n1083), 
        .Q(\IDinst/n8743 ) );
  nnd2s1 \IDinst/U8801  ( .DIN1(\IDinst/RegFile[12][30] ), .DIN2(n1053), 
        .Q(\IDinst/n8742 ) );
  nnd2s1 \IDinst/U8800  ( .DIN1(\IDinst/n8740 ), .DIN2(\IDinst/n8739 ), 
        .Q(\IDinst/n8741 ) );
  nnd2s1 \IDinst/U8799  ( .DIN1(\IDinst/n8738 ), .DIN2(n1165), 
        .Q(\IDinst/n8740 ) );
  nnd2s1 \IDinst/U8798  ( .DIN1(\IDinst/n8735 ), .DIN2(n1144), 
        .Q(\IDinst/n8739 ) );
  nnd2s1 \IDinst/U8797  ( .DIN1(\IDinst/n8737 ), .DIN2(\IDinst/n8736 ), 
        .Q(\IDinst/n8738 ) );
  nnd2s1 \IDinst/U8796  ( .DIN1(\IDinst/RegFile[11][30] ), .DIN2(n1083), 
        .Q(\IDinst/n8737 ) );
  nnd2s1 \IDinst/U8795  ( .DIN1(\IDinst/RegFile[10][30] ), .DIN2(n1053), 
        .Q(\IDinst/n8736 ) );
  nnd2s1 \IDinst/U8794  ( .DIN1(\IDinst/n8734 ), .DIN2(\IDinst/n8733 ), 
        .Q(\IDinst/n8735 ) );
  nnd2s1 \IDinst/U8793  ( .DIN1(\IDinst/RegFile[9][30] ), .DIN2(n1083), 
        .Q(\IDinst/n8734 ) );
  nnd2s1 \IDinst/U8792  ( .DIN1(\IDinst/RegFile[8][30] ), .DIN2(n1053), 
        .Q(\IDinst/n8733 ) );
  nnd2s1 \IDinst/U8791  ( .DIN1(\IDinst/n8731 ), .DIN2(\IDinst/n8730 ), 
        .Q(\IDinst/n8732 ) );
  nnd2s1 \IDinst/U8790  ( .DIN1(\IDinst/n8729 ), .DIN2(\IDinst/N41 ), 
        .Q(\IDinst/n8731 ) );
  nnd2s1 \IDinst/U8789  ( .DIN1(\IDinst/n8720 ), .DIN2(n1189), 
        .Q(\IDinst/n8730 ) );
  nnd2s1 \IDinst/U8788  ( .DIN1(\IDinst/n8728 ), .DIN2(\IDinst/n8727 ), 
        .Q(\IDinst/n8729 ) );
  nnd2s1 \IDinst/U8787  ( .DIN1(\IDinst/n8726 ), .DIN2(n1165), 
        .Q(\IDinst/n8728 ) );
  nnd2s1 \IDinst/U8786  ( .DIN1(\IDinst/n8723 ), .DIN2(n1144), 
        .Q(\IDinst/n8727 ) );
  nnd2s1 \IDinst/U8785  ( .DIN1(\IDinst/n8725 ), .DIN2(\IDinst/n8724 ), 
        .Q(\IDinst/n8726 ) );
  nnd2s1 \IDinst/U8784  ( .DIN1(\IDinst/RegFile[7][30] ), .DIN2(n1084), 
        .Q(\IDinst/n8725 ) );
  nnd2s1 \IDinst/U8783  ( .DIN1(\IDinst/RegFile[6][30] ), .DIN2(n1053), 
        .Q(\IDinst/n8724 ) );
  nnd2s1 \IDinst/U8782  ( .DIN1(\IDinst/n8722 ), .DIN2(\IDinst/n8721 ), 
        .Q(\IDinst/n8723 ) );
  nnd2s1 \IDinst/U8781  ( .DIN1(\IDinst/RegFile[5][30] ), .DIN2(n1084), 
        .Q(\IDinst/n8722 ) );
  nnd2s1 \IDinst/U8780  ( .DIN1(\IDinst/RegFile[4][30] ), .DIN2(n1052), 
        .Q(\IDinst/n8721 ) );
  nnd2s1 \IDinst/U8779  ( .DIN1(\IDinst/n8719 ), .DIN2(\IDinst/n8718 ), 
        .Q(\IDinst/n8720 ) );
  nnd2s1 \IDinst/U8778  ( .DIN1(\IDinst/n8717 ), .DIN2(n1165), 
        .Q(\IDinst/n8719 ) );
  nnd2s1 \IDinst/U8777  ( .DIN1(\IDinst/n8714 ), .DIN2(n1144), 
        .Q(\IDinst/n8718 ) );
  nnd2s1 \IDinst/U8776  ( .DIN1(\IDinst/n8716 ), .DIN2(\IDinst/n8715 ), 
        .Q(\IDinst/n8717 ) );
  nnd2s1 \IDinst/U8775  ( .DIN1(\IDinst/RegFile[3][30] ), .DIN2(n1084), 
        .Q(\IDinst/n8716 ) );
  nnd2s1 \IDinst/U8774  ( .DIN1(\IDinst/RegFile[2][30] ), .DIN2(n1052), 
        .Q(\IDinst/n8715 ) );
  nnd2s1 \IDinst/U8773  ( .DIN1(\IDinst/n8713 ), .DIN2(\IDinst/n8712 ), 
        .Q(\IDinst/n8714 ) );
  nnd2s1 \IDinst/U8772  ( .DIN1(\IDinst/RegFile[1][30] ), .DIN2(n1084), 
        .Q(\IDinst/n8713 ) );
  nnd2s1 \IDinst/U8771  ( .DIN1(\IDinst/RegFile[0][30] ), .DIN2(n1052), 
        .Q(\IDinst/n8712 ) );
  nnd2s1 \IDinst/U8770  ( .DIN1(\IDinst/n8711 ), .DIN2(n539), 
        .Q(\IDinst/n6006 ) );
  nnd2s1 \IDinst/U8769  ( .DIN1(\IDinst/n8666 ), .DIN2(n635), 
        .Q(\IDinst/n6007 ) );
  nnd2s1 \IDinst/U8768  ( .DIN1(\IDinst/n8710 ), .DIN2(\IDinst/n8709 ), 
        .Q(\IDinst/n8711 ) );
  nnd2s1 \IDinst/U8767  ( .DIN1(\IDinst/n8708 ), .DIN2(n643), 
        .Q(\IDinst/n8710 ) );
  nnd2s1 \IDinst/U8766  ( .DIN1(\IDinst/n8687 ), .DIN2(n673), 
        .Q(\IDinst/n8709 ) );
  nnd2s1 \IDinst/U8765  ( .DIN1(\IDinst/n8707 ), .DIN2(\IDinst/n8706 ), 
        .Q(\IDinst/n8708 ) );
  nnd2s1 \IDinst/U8764  ( .DIN1(\IDinst/n8705 ), .DIN2(n1192), 
        .Q(\IDinst/n8707 ) );
  nnd2s1 \IDinst/U8763  ( .DIN1(\IDinst/n8696 ), .DIN2(n1189), 
        .Q(\IDinst/n8706 ) );
  nnd2s1 \IDinst/U8762  ( .DIN1(\IDinst/n8704 ), .DIN2(\IDinst/n8703 ), 
        .Q(\IDinst/n8705 ) );
  nnd2s1 \IDinst/U8761  ( .DIN1(\IDinst/n8702 ), .DIN2(n1165), 
        .Q(\IDinst/n8704 ) );
  nnd2s1 \IDinst/U8760  ( .DIN1(\IDinst/n8699 ), .DIN2(n1144), 
        .Q(\IDinst/n8703 ) );
  nnd2s1 \IDinst/U8759  ( .DIN1(\IDinst/n8701 ), .DIN2(\IDinst/n8700 ), 
        .Q(\IDinst/n8702 ) );
  nnd2s1 \IDinst/U8758  ( .DIN1(\IDinst/RegFile[31][29] ), .DIN2(n1084), 
        .Q(\IDinst/n8701 ) );
  nnd2s1 \IDinst/U8757  ( .DIN1(\IDinst/RegFile[30][29] ), .DIN2(n1052), 
        .Q(\IDinst/n8700 ) );
  nnd2s1 \IDinst/U8756  ( .DIN1(\IDinst/n8698 ), .DIN2(\IDinst/n8697 ), 
        .Q(\IDinst/n8699 ) );
  nnd2s1 \IDinst/U8755  ( .DIN1(\IDinst/RegFile[29][29] ), .DIN2(n1084), 
        .Q(\IDinst/n8698 ) );
  nnd2s1 \IDinst/U8754  ( .DIN1(\IDinst/RegFile[28][29] ), .DIN2(n1052), 
        .Q(\IDinst/n8697 ) );
  nnd2s1 \IDinst/U8753  ( .DIN1(\IDinst/n8695 ), .DIN2(\IDinst/n8694 ), 
        .Q(\IDinst/n8696 ) );
  nnd2s1 \IDinst/U8752  ( .DIN1(\IDinst/n8693 ), .DIN2(n1165), 
        .Q(\IDinst/n8695 ) );
  nnd2s1 \IDinst/U8751  ( .DIN1(\IDinst/n8690 ), .DIN2(n1144), 
        .Q(\IDinst/n8694 ) );
  nnd2s1 \IDinst/U8750  ( .DIN1(\IDinst/n8692 ), .DIN2(\IDinst/n8691 ), 
        .Q(\IDinst/n8693 ) );
  nnd2s1 \IDinst/U8749  ( .DIN1(\IDinst/RegFile[27][29] ), .DIN2(n1084), 
        .Q(\IDinst/n8692 ) );
  nnd2s1 \IDinst/U8748  ( .DIN1(\IDinst/RegFile[26][29] ), .DIN2(n1052), 
        .Q(\IDinst/n8691 ) );
  nnd2s1 \IDinst/U8747  ( .DIN1(\IDinst/n8689 ), .DIN2(\IDinst/n8688 ), 
        .Q(\IDinst/n8690 ) );
  nnd2s1 \IDinst/U8746  ( .DIN1(\IDinst/RegFile[25][29] ), .DIN2(n1084), 
        .Q(\IDinst/n8689 ) );
  nnd2s1 \IDinst/U8745  ( .DIN1(\IDinst/RegFile[24][29] ), .DIN2(n1052), 
        .Q(\IDinst/n8688 ) );
  nnd2s1 \IDinst/U8744  ( .DIN1(\IDinst/n8686 ), .DIN2(\IDinst/n8685 ), 
        .Q(\IDinst/n8687 ) );
  nnd2s1 \IDinst/U8743  ( .DIN1(\IDinst/n8684 ), .DIN2(n1193), 
        .Q(\IDinst/n8686 ) );
  nnd2s1 \IDinst/U8742  ( .DIN1(\IDinst/n8675 ), .DIN2(n1189), 
        .Q(\IDinst/n8685 ) );
  nnd2s1 \IDinst/U8741  ( .DIN1(\IDinst/n8683 ), .DIN2(\IDinst/n8682 ), 
        .Q(\IDinst/n8684 ) );
  nnd2s1 \IDinst/U8740  ( .DIN1(\IDinst/n8681 ), .DIN2(n1165), 
        .Q(\IDinst/n8683 ) );
  nnd2s1 \IDinst/U8739  ( .DIN1(\IDinst/n8678 ), .DIN2(n1145), 
        .Q(\IDinst/n8682 ) );
  nnd2s1 \IDinst/U8738  ( .DIN1(\IDinst/n8680 ), .DIN2(\IDinst/n8679 ), 
        .Q(\IDinst/n8681 ) );
  nnd2s1 \IDinst/U8737  ( .DIN1(\IDinst/RegFile[23][29] ), .DIN2(n1084), 
        .Q(\IDinst/n8680 ) );
  nnd2s1 \IDinst/U8736  ( .DIN1(\IDinst/RegFile[22][29] ), .DIN2(n1052), 
        .Q(\IDinst/n8679 ) );
  nnd2s1 \IDinst/U8735  ( .DIN1(\IDinst/n8677 ), .DIN2(\IDinst/n8676 ), 
        .Q(\IDinst/n8678 ) );
  nnd2s1 \IDinst/U8734  ( .DIN1(\IDinst/RegFile[21][29] ), .DIN2(n1085), 
        .Q(\IDinst/n8677 ) );
  nnd2s1 \IDinst/U8733  ( .DIN1(\IDinst/RegFile[20][29] ), .DIN2(n1052), 
        .Q(\IDinst/n8676 ) );
  nnd2s1 \IDinst/U8732  ( .DIN1(\IDinst/n8674 ), .DIN2(\IDinst/n8673 ), 
        .Q(\IDinst/n8675 ) );
  nnd2s1 \IDinst/U8731  ( .DIN1(\IDinst/n8672 ), .DIN2(n1165), 
        .Q(\IDinst/n8674 ) );
  nnd2s1 \IDinst/U8730  ( .DIN1(\IDinst/n8669 ), .DIN2(n1145), 
        .Q(\IDinst/n8673 ) );
  nnd2s1 \IDinst/U8729  ( .DIN1(\IDinst/n8671 ), .DIN2(\IDinst/n8670 ), 
        .Q(\IDinst/n8672 ) );
  nnd2s1 \IDinst/U8728  ( .DIN1(\IDinst/RegFile[19][29] ), .DIN2(n1085), 
        .Q(\IDinst/n8671 ) );
  nnd2s1 \IDinst/U8727  ( .DIN1(\IDinst/RegFile[18][29] ), .DIN2(n1052), 
        .Q(\IDinst/n8670 ) );
  nnd2s1 \IDinst/U8726  ( .DIN1(\IDinst/n8668 ), .DIN2(\IDinst/n8667 ), 
        .Q(\IDinst/n8669 ) );
  nnd2s1 \IDinst/U8725  ( .DIN1(\IDinst/RegFile[17][29] ), .DIN2(n1085), 
        .Q(\IDinst/n8668 ) );
  nnd2s1 \IDinst/U8724  ( .DIN1(\IDinst/RegFile[16][29] ), .DIN2(n1052), 
        .Q(\IDinst/n8667 ) );
  nnd2s1 \IDinst/U8723  ( .DIN1(\IDinst/n8665 ), .DIN2(\IDinst/n8664 ), 
        .Q(\IDinst/n8666 ) );
  nnd2s1 \IDinst/U8722  ( .DIN1(\IDinst/n8663 ), .DIN2(n642), 
        .Q(\IDinst/n8665 ) );
  nnd2s1 \IDinst/U8721  ( .DIN1(\IDinst/n8642 ), .DIN2(n670), 
        .Q(\IDinst/n8664 ) );
  nnd2s1 \IDinst/U8720  ( .DIN1(\IDinst/n8662 ), .DIN2(\IDinst/n8661 ), 
        .Q(\IDinst/n8663 ) );
  nnd2s1 \IDinst/U8719  ( .DIN1(\IDinst/n8660 ), .DIN2(n1194), 
        .Q(\IDinst/n8662 ) );
  nnd2s1 \IDinst/U8718  ( .DIN1(\IDinst/n8651 ), .DIN2(n1189), 
        .Q(\IDinst/n8661 ) );
  nnd2s1 \IDinst/U8717  ( .DIN1(\IDinst/n8659 ), .DIN2(\IDinst/n8658 ), 
        .Q(\IDinst/n8660 ) );
  nnd2s1 \IDinst/U8716  ( .DIN1(\IDinst/n8657 ), .DIN2(n1165), 
        .Q(\IDinst/n8659 ) );
  nnd2s1 \IDinst/U8715  ( .DIN1(\IDinst/n8654 ), .DIN2(n1145), 
        .Q(\IDinst/n8658 ) );
  nnd2s1 \IDinst/U8714  ( .DIN1(\IDinst/n8656 ), .DIN2(\IDinst/n8655 ), 
        .Q(\IDinst/n8657 ) );
  nnd2s1 \IDinst/U8713  ( .DIN1(\IDinst/RegFile[15][29] ), .DIN2(n1085), 
        .Q(\IDinst/n8656 ) );
  nnd2s1 \IDinst/U8712  ( .DIN1(\IDinst/RegFile[14][29] ), .DIN2(n1052), 
        .Q(\IDinst/n8655 ) );
  nnd2s1 \IDinst/U8711  ( .DIN1(\IDinst/n8653 ), .DIN2(\IDinst/n8652 ), 
        .Q(\IDinst/n8654 ) );
  nnd2s1 \IDinst/U8710  ( .DIN1(\IDinst/RegFile[13][29] ), .DIN2(n1085), 
        .Q(\IDinst/n8653 ) );
  nnd2s1 \IDinst/U8709  ( .DIN1(\IDinst/RegFile[12][29] ), .DIN2(n1052), 
        .Q(\IDinst/n8652 ) );
  nnd2s1 \IDinst/U8708  ( .DIN1(\IDinst/n8650 ), .DIN2(\IDinst/n8649 ), 
        .Q(\IDinst/n8651 ) );
  nnd2s1 \IDinst/U8707  ( .DIN1(\IDinst/n8648 ), .DIN2(n1165), 
        .Q(\IDinst/n8650 ) );
  nnd2s1 \IDinst/U8706  ( .DIN1(\IDinst/n8645 ), .DIN2(n1145), 
        .Q(\IDinst/n8649 ) );
  nnd2s1 \IDinst/U8705  ( .DIN1(\IDinst/n8647 ), .DIN2(\IDinst/n8646 ), 
        .Q(\IDinst/n8648 ) );
  nnd2s1 \IDinst/U8704  ( .DIN1(\IDinst/RegFile[11][29] ), .DIN2(n1085), 
        .Q(\IDinst/n8647 ) );
  nnd2s1 \IDinst/U8703  ( .DIN1(\IDinst/RegFile[10][29] ), .DIN2(n1051), 
        .Q(\IDinst/n8646 ) );
  nnd2s1 \IDinst/U8702  ( .DIN1(\IDinst/n8644 ), .DIN2(\IDinst/n8643 ), 
        .Q(\IDinst/n8645 ) );
  nnd2s1 \IDinst/U8701  ( .DIN1(\IDinst/RegFile[9][29] ), .DIN2(n1085), 
        .Q(\IDinst/n8644 ) );
  nnd2s1 \IDinst/U8700  ( .DIN1(\IDinst/RegFile[8][29] ), .DIN2(n1051), 
        .Q(\IDinst/n8643 ) );
  nnd2s1 \IDinst/U8699  ( .DIN1(\IDinst/n8641 ), .DIN2(\IDinst/n8640 ), 
        .Q(\IDinst/n8642 ) );
  nnd2s1 \IDinst/U8698  ( .DIN1(\IDinst/n8639 ), .DIN2(n1196), 
        .Q(\IDinst/n8641 ) );
  nnd2s1 \IDinst/U8697  ( .DIN1(\IDinst/n8630 ), .DIN2(n1189), 
        .Q(\IDinst/n8640 ) );
  nnd2s1 \IDinst/U8696  ( .DIN1(\IDinst/n8638 ), .DIN2(\IDinst/n8637 ), 
        .Q(\IDinst/n8639 ) );
  nnd2s1 \IDinst/U8695  ( .DIN1(\IDinst/n8636 ), .DIN2(n1164), 
        .Q(\IDinst/n8638 ) );
  nnd2s1 \IDinst/U8694  ( .DIN1(\IDinst/n8633 ), .DIN2(n1145), 
        .Q(\IDinst/n8637 ) );
  nnd2s1 \IDinst/U8693  ( .DIN1(\IDinst/n8635 ), .DIN2(\IDinst/n8634 ), 
        .Q(\IDinst/n8636 ) );
  nnd2s1 \IDinst/U8692  ( .DIN1(\IDinst/RegFile[7][29] ), .DIN2(n1085), 
        .Q(\IDinst/n8635 ) );
  nnd2s1 \IDinst/U8691  ( .DIN1(\IDinst/RegFile[6][29] ), .DIN2(n1051), 
        .Q(\IDinst/n8634 ) );
  nnd2s1 \IDinst/U8690  ( .DIN1(\IDinst/n8632 ), .DIN2(\IDinst/n8631 ), 
        .Q(\IDinst/n8633 ) );
  nnd2s1 \IDinst/U8689  ( .DIN1(\IDinst/RegFile[5][29] ), .DIN2(n1085), 
        .Q(\IDinst/n8632 ) );
  nnd2s1 \IDinst/U8688  ( .DIN1(\IDinst/RegFile[4][29] ), .DIN2(n1051), 
        .Q(\IDinst/n8631 ) );
  nnd2s1 \IDinst/U8687  ( .DIN1(\IDinst/n8629 ), .DIN2(\IDinst/n8628 ), 
        .Q(\IDinst/n8630 ) );
  nnd2s1 \IDinst/U8686  ( .DIN1(\IDinst/n8627 ), .DIN2(n1164), 
        .Q(\IDinst/n8629 ) );
  nnd2s1 \IDinst/U8685  ( .DIN1(\IDinst/n8624 ), .DIN2(n1145), 
        .Q(\IDinst/n8628 ) );
  nnd2s1 \IDinst/U8684  ( .DIN1(\IDinst/n8626 ), .DIN2(\IDinst/n8625 ), 
        .Q(\IDinst/n8627 ) );
  nnd2s1 \IDinst/U8683  ( .DIN1(\IDinst/RegFile[3][29] ), .DIN2(n1086), 
        .Q(\IDinst/n8626 ) );
  nnd2s1 \IDinst/U8682  ( .DIN1(\IDinst/RegFile[2][29] ), .DIN2(n1051), 
        .Q(\IDinst/n8625 ) );
  nnd2s1 \IDinst/U8681  ( .DIN1(\IDinst/n8623 ), .DIN2(\IDinst/n8622 ), 
        .Q(\IDinst/n8624 ) );
  nnd2s1 \IDinst/U8680  ( .DIN1(\IDinst/RegFile[1][29] ), .DIN2(n1086), 
        .Q(\IDinst/n8623 ) );
  nnd2s1 \IDinst/U8679  ( .DIN1(\IDinst/RegFile[0][29] ), .DIN2(n1051), 
        .Q(\IDinst/n8622 ) );
  nnd2s1 \IDinst/U8678  ( .DIN1(\IDinst/n8621 ), .DIN2(n539), 
        .Q(\IDinst/n6004 ) );
  nnd2s1 \IDinst/U8677  ( .DIN1(\IDinst/n8576 ), .DIN2(n636), 
        .Q(\IDinst/n6005 ) );
  nnd2s1 \IDinst/U8676  ( .DIN1(\IDinst/n8620 ), .DIN2(\IDinst/n8619 ), 
        .Q(\IDinst/n8621 ) );
  nnd2s1 \IDinst/U8675  ( .DIN1(\IDinst/n8618 ), .DIN2(n641), 
        .Q(\IDinst/n8620 ) );
  nnd2s1 \IDinst/U8674  ( .DIN1(\IDinst/n8597 ), .DIN2(n673), 
        .Q(\IDinst/n8619 ) );
  nnd2s1 \IDinst/U8673  ( .DIN1(\IDinst/n8617 ), .DIN2(\IDinst/n8616 ), 
        .Q(\IDinst/n8618 ) );
  nnd2s1 \IDinst/U8672  ( .DIN1(\IDinst/n8615 ), .DIN2(n1193), 
        .Q(\IDinst/n8617 ) );
  nnd2s1 \IDinst/U8671  ( .DIN1(\IDinst/n8606 ), .DIN2(n1189), 
        .Q(\IDinst/n8616 ) );
  nnd2s1 \IDinst/U8670  ( .DIN1(\IDinst/n8614 ), .DIN2(\IDinst/n8613 ), 
        .Q(\IDinst/n8615 ) );
  nnd2s1 \IDinst/U8669  ( .DIN1(\IDinst/n8612 ), .DIN2(n1164), 
        .Q(\IDinst/n8614 ) );
  nnd2s1 \IDinst/U8668  ( .DIN1(\IDinst/n8609 ), .DIN2(n1145), 
        .Q(\IDinst/n8613 ) );
  nnd2s1 \IDinst/U8667  ( .DIN1(\IDinst/n8611 ), .DIN2(\IDinst/n8610 ), 
        .Q(\IDinst/n8612 ) );
  nnd2s1 \IDinst/U8666  ( .DIN1(\IDinst/RegFile[31][28] ), .DIN2(n1086), 
        .Q(\IDinst/n8611 ) );
  nnd2s1 \IDinst/U8665  ( .DIN1(\IDinst/RegFile[30][28] ), .DIN2(n1051), 
        .Q(\IDinst/n8610 ) );
  nnd2s1 \IDinst/U8664  ( .DIN1(\IDinst/n8608 ), .DIN2(\IDinst/n8607 ), 
        .Q(\IDinst/n8609 ) );
  nnd2s1 \IDinst/U8663  ( .DIN1(\IDinst/RegFile[29][28] ), .DIN2(n1086), 
        .Q(\IDinst/n8608 ) );
  nnd2s1 \IDinst/U8662  ( .DIN1(\IDinst/RegFile[28][28] ), .DIN2(n1051), 
        .Q(\IDinst/n8607 ) );
  nnd2s1 \IDinst/U8661  ( .DIN1(\IDinst/n8605 ), .DIN2(\IDinst/n8604 ), 
        .Q(\IDinst/n8606 ) );
  nnd2s1 \IDinst/U8660  ( .DIN1(\IDinst/n8603 ), .DIN2(n1164), 
        .Q(\IDinst/n8605 ) );
  nnd2s1 \IDinst/U8659  ( .DIN1(\IDinst/n8600 ), .DIN2(n1145), 
        .Q(\IDinst/n8604 ) );
  nnd2s1 \IDinst/U8658  ( .DIN1(\IDinst/n8602 ), .DIN2(\IDinst/n8601 ), 
        .Q(\IDinst/n8603 ) );
  nnd2s1 \IDinst/U8657  ( .DIN1(\IDinst/RegFile[27][28] ), .DIN2(n1086), 
        .Q(\IDinst/n8602 ) );
  nnd2s1 \IDinst/U8656  ( .DIN1(\IDinst/RegFile[26][28] ), .DIN2(n1051), 
        .Q(\IDinst/n8601 ) );
  nnd2s1 \IDinst/U8655  ( .DIN1(\IDinst/n8599 ), .DIN2(\IDinst/n8598 ), 
        .Q(\IDinst/n8600 ) );
  nnd2s1 \IDinst/U8654  ( .DIN1(\IDinst/RegFile[25][28] ), .DIN2(n1086), 
        .Q(\IDinst/n8599 ) );
  nnd2s1 \IDinst/U8653  ( .DIN1(\IDinst/RegFile[24][28] ), .DIN2(n1051), 
        .Q(\IDinst/n8598 ) );
  nnd2s1 \IDinst/U8652  ( .DIN1(\IDinst/n8596 ), .DIN2(\IDinst/n8595 ), 
        .Q(\IDinst/n8597 ) );
  nnd2s1 \IDinst/U8651  ( .DIN1(\IDinst/n8594 ), .DIN2(n1193), 
        .Q(\IDinst/n8596 ) );
  nnd2s1 \IDinst/U8650  ( .DIN1(\IDinst/n8585 ), .DIN2(n1189), 
        .Q(\IDinst/n8595 ) );
  nnd2s1 \IDinst/U8649  ( .DIN1(\IDinst/n8593 ), .DIN2(\IDinst/n8592 ), 
        .Q(\IDinst/n8594 ) );
  nnd2s1 \IDinst/U8648  ( .DIN1(\IDinst/n8591 ), .DIN2(n1164), 
        .Q(\IDinst/n8593 ) );
  nnd2s1 \IDinst/U8647  ( .DIN1(\IDinst/n8588 ), .DIN2(n1145), 
        .Q(\IDinst/n8592 ) );
  nnd2s1 \IDinst/U8646  ( .DIN1(\IDinst/n8590 ), .DIN2(\IDinst/n8589 ), 
        .Q(\IDinst/n8591 ) );
  nnd2s1 \IDinst/U8645  ( .DIN1(\IDinst/RegFile[23][28] ), .DIN2(n1086), 
        .Q(\IDinst/n8590 ) );
  nnd2s1 \IDinst/U8644  ( .DIN1(\IDinst/RegFile[22][28] ), .DIN2(n1051), 
        .Q(\IDinst/n8589 ) );
  nnd2s1 \IDinst/U8643  ( .DIN1(\IDinst/n8587 ), .DIN2(\IDinst/n8586 ), 
        .Q(\IDinst/n8588 ) );
  nnd2s1 \IDinst/U8642  ( .DIN1(\IDinst/RegFile[21][28] ), .DIN2(n1086), 
        .Q(\IDinst/n8587 ) );
  nnd2s1 \IDinst/U8641  ( .DIN1(\IDinst/RegFile[20][28] ), .DIN2(n1051), 
        .Q(\IDinst/n8586 ) );
  nnd2s1 \IDinst/U8640  ( .DIN1(\IDinst/n8584 ), .DIN2(\IDinst/n8583 ), 
        .Q(\IDinst/n8585 ) );
  nnd2s1 \IDinst/U8639  ( .DIN1(\IDinst/n8582 ), .DIN2(n1164), 
        .Q(\IDinst/n8584 ) );
  nnd2s1 \IDinst/U8638  ( .DIN1(\IDinst/n8579 ), .DIN2(n1145), 
        .Q(\IDinst/n8583 ) );
  nnd2s1 \IDinst/U8637  ( .DIN1(\IDinst/n8581 ), .DIN2(\IDinst/n8580 ), 
        .Q(\IDinst/n8582 ) );
  nnd2s1 \IDinst/U8636  ( .DIN1(\IDinst/RegFile[19][28] ), .DIN2(n1086), 
        .Q(\IDinst/n8581 ) );
  nnd2s1 \IDinst/U8635  ( .DIN1(\IDinst/RegFile[18][28] ), .DIN2(n1051), 
        .Q(\IDinst/n8580 ) );
  nnd2s1 \IDinst/U8634  ( .DIN1(\IDinst/n8578 ), .DIN2(\IDinst/n8577 ), 
        .Q(\IDinst/n8579 ) );
  nnd2s1 \IDinst/U8633  ( .DIN1(\IDinst/RegFile[17][28] ), .DIN2(n1087), 
        .Q(\IDinst/n8578 ) );
  nnd2s1 \IDinst/U8632  ( .DIN1(\IDinst/RegFile[16][28] ), .DIN2(n1050), 
        .Q(\IDinst/n8577 ) );
  nnd2s1 \IDinst/U8631  ( .DIN1(\IDinst/n8575 ), .DIN2(\IDinst/n8574 ), 
        .Q(\IDinst/n8576 ) );
  nnd2s1 \IDinst/U8630  ( .DIN1(\IDinst/n8573 ), .DIN2(n644), 
        .Q(\IDinst/n8575 ) );
  nnd2s1 \IDinst/U8629  ( .DIN1(\IDinst/n8552 ), .DIN2(n670), 
        .Q(\IDinst/n8574 ) );
  nnd2s1 \IDinst/U8628  ( .DIN1(\IDinst/n8572 ), .DIN2(\IDinst/n8571 ), 
        .Q(\IDinst/n8573 ) );
  nnd2s1 \IDinst/U8627  ( .DIN1(\IDinst/n8570 ), .DIN2(n1192), 
        .Q(\IDinst/n8572 ) );
  nnd2s1 \IDinst/U8626  ( .DIN1(\IDinst/n8561 ), .DIN2(n1189), 
        .Q(\IDinst/n8571 ) );
  nnd2s1 \IDinst/U8625  ( .DIN1(\IDinst/n8569 ), .DIN2(\IDinst/n8568 ), 
        .Q(\IDinst/n8570 ) );
  nnd2s1 \IDinst/U8624  ( .DIN1(\IDinst/n8567 ), .DIN2(n1164), 
        .Q(\IDinst/n8569 ) );
  nnd2s1 \IDinst/U8623  ( .DIN1(\IDinst/n8564 ), .DIN2(n1145), 
        .Q(\IDinst/n8568 ) );
  nnd2s1 \IDinst/U8622  ( .DIN1(\IDinst/n8566 ), .DIN2(\IDinst/n8565 ), 
        .Q(\IDinst/n8567 ) );
  nnd2s1 \IDinst/U8621  ( .DIN1(\IDinst/RegFile[15][28] ), .DIN2(n1087), 
        .Q(\IDinst/n8566 ) );
  nnd2s1 \IDinst/U8620  ( .DIN1(\IDinst/RegFile[14][28] ), .DIN2(n1050), 
        .Q(\IDinst/n8565 ) );
  nnd2s1 \IDinst/U8619  ( .DIN1(\IDinst/n8563 ), .DIN2(\IDinst/n8562 ), 
        .Q(\IDinst/n8564 ) );
  nnd2s1 \IDinst/U8618  ( .DIN1(\IDinst/RegFile[13][28] ), .DIN2(n1087), 
        .Q(\IDinst/n8563 ) );
  nnd2s1 \IDinst/U8617  ( .DIN1(\IDinst/RegFile[12][28] ), .DIN2(n1050), 
        .Q(\IDinst/n8562 ) );
  nnd2s1 \IDinst/U8616  ( .DIN1(\IDinst/n8560 ), .DIN2(\IDinst/n8559 ), 
        .Q(\IDinst/n8561 ) );
  nnd2s1 \IDinst/U8615  ( .DIN1(\IDinst/n8558 ), .DIN2(n1164), 
        .Q(\IDinst/n8560 ) );
  nnd2s1 \IDinst/U8614  ( .DIN1(\IDinst/n8555 ), .DIN2(n1145), 
        .Q(\IDinst/n8559 ) );
  nnd2s1 \IDinst/U8613  ( .DIN1(\IDinst/n8557 ), .DIN2(\IDinst/n8556 ), 
        .Q(\IDinst/n8558 ) );
  nnd2s1 \IDinst/U8612  ( .DIN1(\IDinst/RegFile[11][28] ), .DIN2(n1087), 
        .Q(\IDinst/n8557 ) );
  nnd2s1 \IDinst/U8611  ( .DIN1(\IDinst/RegFile[10][28] ), .DIN2(n1050), 
        .Q(\IDinst/n8556 ) );
  nnd2s1 \IDinst/U8610  ( .DIN1(\IDinst/n8554 ), .DIN2(\IDinst/n8553 ), 
        .Q(\IDinst/n8555 ) );
  nnd2s1 \IDinst/U8609  ( .DIN1(\IDinst/RegFile[9][28] ), .DIN2(n1087), 
        .Q(\IDinst/n8554 ) );
  nnd2s1 \IDinst/U8608  ( .DIN1(\IDinst/RegFile[8][28] ), .DIN2(n1050), 
        .Q(\IDinst/n8553 ) );
  nnd2s1 \IDinst/U8607  ( .DIN1(\IDinst/n8551 ), .DIN2(\IDinst/n8550 ), 
        .Q(\IDinst/n8552 ) );
  nnd2s1 \IDinst/U8606  ( .DIN1(\IDinst/n8549 ), .DIN2(n1191), 
        .Q(\IDinst/n8551 ) );
  nnd2s1 \IDinst/U8605  ( .DIN1(\IDinst/n8540 ), .DIN2(n1189), 
        .Q(\IDinst/n8550 ) );
  nnd2s1 \IDinst/U8604  ( .DIN1(\IDinst/n8548 ), .DIN2(\IDinst/n8547 ), 
        .Q(\IDinst/n8549 ) );
  nnd2s1 \IDinst/U8603  ( .DIN1(\IDinst/n8546 ), .DIN2(n1164), 
        .Q(\IDinst/n8548 ) );
  nnd2s1 \IDinst/U8602  ( .DIN1(\IDinst/n8543 ), .DIN2(n1145), 
        .Q(\IDinst/n8547 ) );
  nnd2s1 \IDinst/U8601  ( .DIN1(\IDinst/n8545 ), .DIN2(\IDinst/n8544 ), 
        .Q(\IDinst/n8546 ) );
  nnd2s1 \IDinst/U8600  ( .DIN1(\IDinst/RegFile[7][28] ), .DIN2(n1087), 
        .Q(\IDinst/n8545 ) );
  nnd2s1 \IDinst/U8599  ( .DIN1(\IDinst/RegFile[6][28] ), .DIN2(n1050), 
        .Q(\IDinst/n8544 ) );
  nnd2s1 \IDinst/U8598  ( .DIN1(\IDinst/n8542 ), .DIN2(\IDinst/n8541 ), 
        .Q(\IDinst/n8543 ) );
  nnd2s1 \IDinst/U8597  ( .DIN1(\IDinst/RegFile[5][28] ), .DIN2(n1087), 
        .Q(\IDinst/n8542 ) );
  nnd2s1 \IDinst/U8596  ( .DIN1(\IDinst/RegFile[4][28] ), .DIN2(n1050), 
        .Q(\IDinst/n8541 ) );
  nnd2s1 \IDinst/U8595  ( .DIN1(\IDinst/n8539 ), .DIN2(\IDinst/n8538 ), 
        .Q(\IDinst/n8540 ) );
  nnd2s1 \IDinst/U8594  ( .DIN1(\IDinst/n8537 ), .DIN2(n1163), 
        .Q(\IDinst/n8539 ) );
  nnd2s1 \IDinst/U8593  ( .DIN1(\IDinst/n8534 ), .DIN2(n1148), 
        .Q(\IDinst/n8538 ) );
  nnd2s1 \IDinst/U8592  ( .DIN1(\IDinst/n8536 ), .DIN2(\IDinst/n8535 ), 
        .Q(\IDinst/n8537 ) );
  nnd2s1 \IDinst/U8591  ( .DIN1(\IDinst/RegFile[3][28] ), .DIN2(n1087), 
        .Q(\IDinst/n8536 ) );
  nnd2s1 \IDinst/U8590  ( .DIN1(\IDinst/RegFile[2][28] ), .DIN2(n1050), 
        .Q(\IDinst/n8535 ) );
  nnd2s1 \IDinst/U8589  ( .DIN1(\IDinst/n8533 ), .DIN2(\IDinst/n8532 ), 
        .Q(\IDinst/n8534 ) );
  nnd2s1 \IDinst/U8588  ( .DIN1(\IDinst/RegFile[1][28] ), .DIN2(n1087), 
        .Q(\IDinst/n8533 ) );
  nnd2s1 \IDinst/U8587  ( .DIN1(\IDinst/RegFile[0][28] ), .DIN2(n1055), 
        .Q(\IDinst/n8532 ) );
  nnd2s1 \IDinst/U8586  ( .DIN1(\IDinst/n8531 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n6002 ) );
  nnd2s1 \IDinst/U8585  ( .DIN1(\IDinst/n8486 ), .DIN2(n635), 
        .Q(\IDinst/n6003 ) );
  nnd2s1 \IDinst/U8584  ( .DIN1(\IDinst/n8530 ), .DIN2(\IDinst/n8529 ), 
        .Q(\IDinst/n8531 ) );
  nnd2s1 \IDinst/U8583  ( .DIN1(\IDinst/n8528 ), .DIN2(n643), 
        .Q(\IDinst/n8530 ) );
  nnd2s1 \IDinst/U8582  ( .DIN1(\IDinst/n8507 ), .DIN2(n670), 
        .Q(\IDinst/n8529 ) );
  nnd2s1 \IDinst/U8581  ( .DIN1(\IDinst/n8527 ), .DIN2(\IDinst/n8526 ), 
        .Q(\IDinst/n8528 ) );
  nnd2s1 \IDinst/U8580  ( .DIN1(\IDinst/n8525 ), .DIN2(n1194), 
        .Q(\IDinst/n8527 ) );
  nnd2s1 \IDinst/U8579  ( .DIN1(\IDinst/n8516 ), .DIN2(n1189), 
        .Q(\IDinst/n8526 ) );
  nnd2s1 \IDinst/U8578  ( .DIN1(\IDinst/n8524 ), .DIN2(\IDinst/n8523 ), 
        .Q(\IDinst/n8525 ) );
  nnd2s1 \IDinst/U8577  ( .DIN1(\IDinst/n8522 ), .DIN2(n1163), 
        .Q(\IDinst/n8524 ) );
  nnd2s1 \IDinst/U8576  ( .DIN1(\IDinst/n8519 ), .DIN2(n1146), 
        .Q(\IDinst/n8523 ) );
  nnd2s1 \IDinst/U8575  ( .DIN1(\IDinst/n8521 ), .DIN2(\IDinst/n8520 ), 
        .Q(\IDinst/n8522 ) );
  nnd2s1 \IDinst/U8574  ( .DIN1(\IDinst/RegFile[31][27] ), .DIN2(n1088), 
        .Q(\IDinst/n8521 ) );
  nnd2s1 \IDinst/U8573  ( .DIN1(\IDinst/RegFile[30][27] ), .DIN2(n1050), 
        .Q(\IDinst/n8520 ) );
  nnd2s1 \IDinst/U8572  ( .DIN1(\IDinst/n8518 ), .DIN2(\IDinst/n8517 ), 
        .Q(\IDinst/n8519 ) );
  nnd2s1 \IDinst/U8571  ( .DIN1(\IDinst/RegFile[29][27] ), .DIN2(n1088), 
        .Q(\IDinst/n8518 ) );
  nnd2s1 \IDinst/U8570  ( .DIN1(\IDinst/RegFile[28][27] ), .DIN2(n1050), 
        .Q(\IDinst/n8517 ) );
  nnd2s1 \IDinst/U8569  ( .DIN1(\IDinst/n8515 ), .DIN2(\IDinst/n8514 ), 
        .Q(\IDinst/n8516 ) );
  nnd2s1 \IDinst/U8568  ( .DIN1(\IDinst/n8513 ), .DIN2(n1163), 
        .Q(\IDinst/n8515 ) );
  nnd2s1 \IDinst/U8567  ( .DIN1(\IDinst/n8510 ), .DIN2(n1146), 
        .Q(\IDinst/n8514 ) );
  nnd2s1 \IDinst/U8566  ( .DIN1(\IDinst/n8512 ), .DIN2(\IDinst/n8511 ), 
        .Q(\IDinst/n8513 ) );
  nnd2s1 \IDinst/U8565  ( .DIN1(\IDinst/RegFile[27][27] ), .DIN2(n1088), 
        .Q(\IDinst/n8512 ) );
  nnd2s1 \IDinst/U8564  ( .DIN1(\IDinst/RegFile[26][27] ), .DIN2(n1050), 
        .Q(\IDinst/n8511 ) );
  nnd2s1 \IDinst/U8563  ( .DIN1(\IDinst/n8509 ), .DIN2(\IDinst/n8508 ), 
        .Q(\IDinst/n8510 ) );
  nnd2s1 \IDinst/U8562  ( .DIN1(\IDinst/RegFile[25][27] ), .DIN2(n1088), 
        .Q(\IDinst/n8509 ) );
  nnd2s1 \IDinst/U8561  ( .DIN1(\IDinst/RegFile[24][27] ), .DIN2(n1050), 
        .Q(\IDinst/n8508 ) );
  nnd2s1 \IDinst/U8560  ( .DIN1(\IDinst/n8506 ), .DIN2(\IDinst/n8505 ), 
        .Q(\IDinst/n8507 ) );
  nnd2s1 \IDinst/U8559  ( .DIN1(\IDinst/n8504 ), .DIN2(n1197), 
        .Q(\IDinst/n8506 ) );
  nnd2s1 \IDinst/U8558  ( .DIN1(\IDinst/n8495 ), .DIN2(n1189), 
        .Q(\IDinst/n8505 ) );
  nnd2s1 \IDinst/U8557  ( .DIN1(\IDinst/n8503 ), .DIN2(\IDinst/n8502 ), 
        .Q(\IDinst/n8504 ) );
  nnd2s1 \IDinst/U8556  ( .DIN1(\IDinst/n8501 ), .DIN2(n1163), 
        .Q(\IDinst/n8503 ) );
  nnd2s1 \IDinst/U8555  ( .DIN1(\IDinst/n8498 ), .DIN2(n1146), 
        .Q(\IDinst/n8502 ) );
  nnd2s1 \IDinst/U8554  ( .DIN1(\IDinst/n8500 ), .DIN2(\IDinst/n8499 ), 
        .Q(\IDinst/n8501 ) );
  nnd2s1 \IDinst/U8553  ( .DIN1(\IDinst/RegFile[23][27] ), .DIN2(n1088), 
        .Q(\IDinst/n8500 ) );
  nnd2s1 \IDinst/U8552  ( .DIN1(\IDinst/RegFile[22][27] ), .DIN2(n1049), 
        .Q(\IDinst/n8499 ) );
  nnd2s1 \IDinst/U8551  ( .DIN1(\IDinst/n8497 ), .DIN2(\IDinst/n8496 ), 
        .Q(\IDinst/n8498 ) );
  nnd2s1 \IDinst/U8550  ( .DIN1(\IDinst/RegFile[21][27] ), .DIN2(n1088), 
        .Q(\IDinst/n8497 ) );
  nnd2s1 \IDinst/U8549  ( .DIN1(\IDinst/RegFile[20][27] ), .DIN2(n1049), 
        .Q(\IDinst/n8496 ) );
  nnd2s1 \IDinst/U8548  ( .DIN1(\IDinst/n8494 ), .DIN2(\IDinst/n8493 ), 
        .Q(\IDinst/n8495 ) );
  nnd2s1 \IDinst/U8547  ( .DIN1(\IDinst/n8492 ), .DIN2(n1163), 
        .Q(\IDinst/n8494 ) );
  nnd2s1 \IDinst/U8546  ( .DIN1(\IDinst/n8489 ), .DIN2(n1146), 
        .Q(\IDinst/n8493 ) );
  nnd2s1 \IDinst/U8545  ( .DIN1(\IDinst/n8491 ), .DIN2(\IDinst/n8490 ), 
        .Q(\IDinst/n8492 ) );
  nnd2s1 \IDinst/U8544  ( .DIN1(\IDinst/RegFile[19][27] ), .DIN2(n1088), 
        .Q(\IDinst/n8491 ) );
  nnd2s1 \IDinst/U8543  ( .DIN1(\IDinst/RegFile[18][27] ), .DIN2(n1049), 
        .Q(\IDinst/n8490 ) );
  nnd2s1 \IDinst/U8542  ( .DIN1(\IDinst/n8488 ), .DIN2(\IDinst/n8487 ), 
        .Q(\IDinst/n8489 ) );
  nnd2s1 \IDinst/U8541  ( .DIN1(\IDinst/RegFile[17][27] ), .DIN2(n1088), 
        .Q(\IDinst/n8488 ) );
  nnd2s1 \IDinst/U8540  ( .DIN1(\IDinst/RegFile[16][27] ), .DIN2(n1049), 
        .Q(\IDinst/n8487 ) );
  nnd2s1 \IDinst/U8539  ( .DIN1(\IDinst/n8485 ), .DIN2(\IDinst/n8484 ), 
        .Q(\IDinst/n8486 ) );
  nnd2s1 \IDinst/U8538  ( .DIN1(\IDinst/n8483 ), .DIN2(n642), 
        .Q(\IDinst/n8485 ) );
  nnd2s1 \IDinst/U8537  ( .DIN1(\IDinst/n8462 ), .DIN2(n673), 
        .Q(\IDinst/n8484 ) );
  nnd2s1 \IDinst/U8536  ( .DIN1(\IDinst/n8482 ), .DIN2(\IDinst/n8481 ), 
        .Q(\IDinst/n8483 ) );
  nnd2s1 \IDinst/U8535  ( .DIN1(\IDinst/n8480 ), .DIN2(n1196), 
        .Q(\IDinst/n8482 ) );
  nnd2s1 \IDinst/U8534  ( .DIN1(\IDinst/n8471 ), .DIN2(n1189), 
        .Q(\IDinst/n8481 ) );
  nnd2s1 \IDinst/U8533  ( .DIN1(\IDinst/n8479 ), .DIN2(\IDinst/n8478 ), 
        .Q(\IDinst/n8480 ) );
  nnd2s1 \IDinst/U8532  ( .DIN1(\IDinst/n8477 ), .DIN2(n1163), 
        .Q(\IDinst/n8479 ) );
  nnd2s1 \IDinst/U8531  ( .DIN1(\IDinst/n8474 ), .DIN2(n1146), 
        .Q(\IDinst/n8478 ) );
  nnd2s1 \IDinst/U8530  ( .DIN1(\IDinst/n8476 ), .DIN2(\IDinst/n8475 ), 
        .Q(\IDinst/n8477 ) );
  nnd2s1 \IDinst/U8529  ( .DIN1(\IDinst/RegFile[15][27] ), .DIN2(n1089), 
        .Q(\IDinst/n8476 ) );
  nnd2s1 \IDinst/U8528  ( .DIN1(\IDinst/RegFile[14][27] ), .DIN2(n1049), 
        .Q(\IDinst/n8475 ) );
  nnd2s1 \IDinst/U8527  ( .DIN1(\IDinst/n8473 ), .DIN2(\IDinst/n8472 ), 
        .Q(\IDinst/n8474 ) );
  nnd2s1 \IDinst/U8526  ( .DIN1(\IDinst/RegFile[13][27] ), .DIN2(n1089), 
        .Q(\IDinst/n8473 ) );
  nnd2s1 \IDinst/U8525  ( .DIN1(\IDinst/RegFile[12][27] ), .DIN2(n1049), 
        .Q(\IDinst/n8472 ) );
  nnd2s1 \IDinst/U8524  ( .DIN1(\IDinst/n8470 ), .DIN2(\IDinst/n8469 ), 
        .Q(\IDinst/n8471 ) );
  nnd2s1 \IDinst/U8523  ( .DIN1(\IDinst/n8468 ), .DIN2(n1163), 
        .Q(\IDinst/n8470 ) );
  nnd2s1 \IDinst/U8522  ( .DIN1(\IDinst/n8465 ), .DIN2(n1146), 
        .Q(\IDinst/n8469 ) );
  nnd2s1 \IDinst/U8521  ( .DIN1(\IDinst/n8467 ), .DIN2(\IDinst/n8466 ), 
        .Q(\IDinst/n8468 ) );
  nnd2s1 \IDinst/U8520  ( .DIN1(\IDinst/RegFile[11][27] ), .DIN2(n1089), 
        .Q(\IDinst/n8467 ) );
  nnd2s1 \IDinst/U8519  ( .DIN1(\IDinst/RegFile[10][27] ), .DIN2(n1049), 
        .Q(\IDinst/n8466 ) );
  nnd2s1 \IDinst/U8518  ( .DIN1(\IDinst/n8464 ), .DIN2(\IDinst/n8463 ), 
        .Q(\IDinst/n8465 ) );
  nnd2s1 \IDinst/U8517  ( .DIN1(\IDinst/RegFile[9][27] ), .DIN2(n1089), 
        .Q(\IDinst/n8464 ) );
  nnd2s1 \IDinst/U8516  ( .DIN1(\IDinst/RegFile[8][27] ), .DIN2(n1049), 
        .Q(\IDinst/n8463 ) );
  nnd2s1 \IDinst/U8515  ( .DIN1(\IDinst/n8461 ), .DIN2(\IDinst/n8460 ), 
        .Q(\IDinst/n8462 ) );
  nnd2s1 \IDinst/U8514  ( .DIN1(\IDinst/n8459 ), .DIN2(\IDinst/N41 ), 
        .Q(\IDinst/n8461 ) );
  nnd2s1 \IDinst/U8513  ( .DIN1(\IDinst/n8450 ), .DIN2(n1188), 
        .Q(\IDinst/n8460 ) );
  nnd2s1 \IDinst/U8512  ( .DIN1(\IDinst/n8458 ), .DIN2(\IDinst/n8457 ), 
        .Q(\IDinst/n8459 ) );
  nnd2s1 \IDinst/U8511  ( .DIN1(\IDinst/n8456 ), .DIN2(n1163), 
        .Q(\IDinst/n8458 ) );
  nnd2s1 \IDinst/U8510  ( .DIN1(\IDinst/n8453 ), .DIN2(n1146), 
        .Q(\IDinst/n8457 ) );
  nnd2s1 \IDinst/U8509  ( .DIN1(\IDinst/n8455 ), .DIN2(\IDinst/n8454 ), 
        .Q(\IDinst/n8456 ) );
  nnd2s1 \IDinst/U8508  ( .DIN1(\IDinst/RegFile[7][27] ), .DIN2(n1089), 
        .Q(\IDinst/n8455 ) );
  nnd2s1 \IDinst/U8507  ( .DIN1(\IDinst/RegFile[6][27] ), .DIN2(n1049), 
        .Q(\IDinst/n8454 ) );
  nnd2s1 \IDinst/U8506  ( .DIN1(\IDinst/n8452 ), .DIN2(\IDinst/n8451 ), 
        .Q(\IDinst/n8453 ) );
  nnd2s1 \IDinst/U8505  ( .DIN1(\IDinst/RegFile[5][27] ), .DIN2(n1089), 
        .Q(\IDinst/n8452 ) );
  nnd2s1 \IDinst/U8504  ( .DIN1(\IDinst/RegFile[4][27] ), .DIN2(n1049), 
        .Q(\IDinst/n8451 ) );
  nnd2s1 \IDinst/U8503  ( .DIN1(\IDinst/n8449 ), .DIN2(\IDinst/n8448 ), 
        .Q(\IDinst/n8450 ) );
  nnd2s1 \IDinst/U8502  ( .DIN1(\IDinst/n8447 ), .DIN2(n1163), 
        .Q(\IDinst/n8449 ) );
  nnd2s1 \IDinst/U8501  ( .DIN1(\IDinst/n8444 ), .DIN2(n1146), 
        .Q(\IDinst/n8448 ) );
  nnd2s1 \IDinst/U8500  ( .DIN1(\IDinst/n8446 ), .DIN2(\IDinst/n8445 ), 
        .Q(\IDinst/n8447 ) );
  nnd2s1 \IDinst/U8499  ( .DIN1(\IDinst/RegFile[3][27] ), .DIN2(n1089), 
        .Q(\IDinst/n8446 ) );
  nnd2s1 \IDinst/U8498  ( .DIN1(\IDinst/RegFile[2][27] ), .DIN2(n1049), 
        .Q(\IDinst/n8445 ) );
  nnd2s1 \IDinst/U8497  ( .DIN1(\IDinst/n8443 ), .DIN2(\IDinst/n8442 ), 
        .Q(\IDinst/n8444 ) );
  nnd2s1 \IDinst/U8496  ( .DIN1(\IDinst/RegFile[1][27] ), .DIN2(n1089), 
        .Q(\IDinst/n8443 ) );
  nnd2s1 \IDinst/U8495  ( .DIN1(\IDinst/RegFile[0][27] ), .DIN2(n1049), 
        .Q(\IDinst/n8442 ) );
  nnd2s1 \IDinst/U8494  ( .DIN1(\IDinst/n8441 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n6000 ) );
  nnd2s1 \IDinst/U8493  ( .DIN1(\IDinst/n8396 ), .DIN2(n636), 
        .Q(\IDinst/n6001 ) );
  nnd2s1 \IDinst/U8492  ( .DIN1(\IDinst/n8440 ), .DIN2(\IDinst/n8439 ), 
        .Q(\IDinst/n8441 ) );
  nnd2s1 \IDinst/U8491  ( .DIN1(\IDinst/n8438 ), .DIN2(n641), 
        .Q(\IDinst/n8440 ) );
  nnd2s1 \IDinst/U8490  ( .DIN1(\IDinst/n8417 ), .DIN2(n671), 
        .Q(\IDinst/n8439 ) );
  nnd2s1 \IDinst/U8489  ( .DIN1(\IDinst/n8437 ), .DIN2(\IDinst/n8436 ), 
        .Q(\IDinst/n8438 ) );
  nnd2s1 \IDinst/U8488  ( .DIN1(\IDinst/n8435 ), .DIN2(n1195), 
        .Q(\IDinst/n8437 ) );
  nnd2s1 \IDinst/U8487  ( .DIN1(\IDinst/n8426 ), .DIN2(n1188), 
        .Q(\IDinst/n8436 ) );
  nnd2s1 \IDinst/U8486  ( .DIN1(\IDinst/n8434 ), .DIN2(\IDinst/n8433 ), 
        .Q(\IDinst/n8435 ) );
  nnd2s1 \IDinst/U8485  ( .DIN1(\IDinst/n8432 ), .DIN2(n1162), 
        .Q(\IDinst/n8434 ) );
  nnd2s1 \IDinst/U8484  ( .DIN1(\IDinst/n8429 ), .DIN2(n1146), 
        .Q(\IDinst/n8433 ) );
  nnd2s1 \IDinst/U8483  ( .DIN1(\IDinst/n8431 ), .DIN2(\IDinst/n8430 ), 
        .Q(\IDinst/n8432 ) );
  nnd2s1 \IDinst/U8482  ( .DIN1(\IDinst/RegFile[31][26] ), .DIN2(n1089), 
        .Q(\IDinst/n8431 ) );
  nnd2s1 \IDinst/U8481  ( .DIN1(\IDinst/RegFile[30][26] ), .DIN2(n1049), 
        .Q(\IDinst/n8430 ) );
  nnd2s1 \IDinst/U8480  ( .DIN1(\IDinst/n8428 ), .DIN2(\IDinst/n8427 ), 
        .Q(\IDinst/n8429 ) );
  nnd2s1 \IDinst/U8479  ( .DIN1(\IDinst/RegFile[29][26] ), .DIN2(n1090), 
        .Q(\IDinst/n8428 ) );
  nnd2s1 \IDinst/U8478  ( .DIN1(\IDinst/RegFile[28][26] ), .DIN2(n1048), 
        .Q(\IDinst/n8427 ) );
  nnd2s1 \IDinst/U8477  ( .DIN1(\IDinst/n8425 ), .DIN2(\IDinst/n8424 ), 
        .Q(\IDinst/n8426 ) );
  nnd2s1 \IDinst/U8476  ( .DIN1(\IDinst/n8423 ), .DIN2(n1162), 
        .Q(\IDinst/n8425 ) );
  nnd2s1 \IDinst/U8475  ( .DIN1(\IDinst/n8420 ), .DIN2(n1146), 
        .Q(\IDinst/n8424 ) );
  nnd2s1 \IDinst/U8474  ( .DIN1(\IDinst/n8422 ), .DIN2(\IDinst/n8421 ), 
        .Q(\IDinst/n8423 ) );
  nnd2s1 \IDinst/U8473  ( .DIN1(\IDinst/RegFile[27][26] ), .DIN2(n1090), 
        .Q(\IDinst/n8422 ) );
  nnd2s1 \IDinst/U8472  ( .DIN1(\IDinst/RegFile[26][26] ), .DIN2(n1048), 
        .Q(\IDinst/n8421 ) );
  nnd2s1 \IDinst/U8471  ( .DIN1(\IDinst/n8419 ), .DIN2(\IDinst/n8418 ), 
        .Q(\IDinst/n8420 ) );
  nnd2s1 \IDinst/U8470  ( .DIN1(\IDinst/RegFile[25][26] ), .DIN2(n1090), 
        .Q(\IDinst/n8419 ) );
  nnd2s1 \IDinst/U8469  ( .DIN1(\IDinst/RegFile[24][26] ), .DIN2(n1048), 
        .Q(\IDinst/n8418 ) );
  nnd2s1 \IDinst/U8468  ( .DIN1(\IDinst/n8416 ), .DIN2(\IDinst/n8415 ), 
        .Q(\IDinst/n8417 ) );
  nnd2s1 \IDinst/U8467  ( .DIN1(\IDinst/n8414 ), .DIN2(n1191), 
        .Q(\IDinst/n8416 ) );
  nnd2s1 \IDinst/U8466  ( .DIN1(\IDinst/n8405 ), .DIN2(n1188), 
        .Q(\IDinst/n8415 ) );
  nnd2s1 \IDinst/U8465  ( .DIN1(\IDinst/n8413 ), .DIN2(\IDinst/n8412 ), 
        .Q(\IDinst/n8414 ) );
  nnd2s1 \IDinst/U8464  ( .DIN1(\IDinst/n8411 ), .DIN2(n1162), 
        .Q(\IDinst/n8413 ) );
  nnd2s1 \IDinst/U8463  ( .DIN1(\IDinst/n8408 ), .DIN2(n1146), 
        .Q(\IDinst/n8412 ) );
  nnd2s1 \IDinst/U8462  ( .DIN1(\IDinst/n8410 ), .DIN2(\IDinst/n8409 ), 
        .Q(\IDinst/n8411 ) );
  nnd2s1 \IDinst/U8461  ( .DIN1(\IDinst/RegFile[23][26] ), .DIN2(n1090), 
        .Q(\IDinst/n8410 ) );
  nnd2s1 \IDinst/U8460  ( .DIN1(\IDinst/RegFile[22][26] ), .DIN2(n1048), 
        .Q(\IDinst/n8409 ) );
  nnd2s1 \IDinst/U8459  ( .DIN1(\IDinst/n8407 ), .DIN2(\IDinst/n8406 ), 
        .Q(\IDinst/n8408 ) );
  nnd2s1 \IDinst/U8458  ( .DIN1(\IDinst/RegFile[21][26] ), .DIN2(n1090), 
        .Q(\IDinst/n8407 ) );
  nnd2s1 \IDinst/U8457  ( .DIN1(\IDinst/RegFile[20][26] ), .DIN2(n1048), 
        .Q(\IDinst/n8406 ) );
  nnd2s1 \IDinst/U8456  ( .DIN1(\IDinst/n8404 ), .DIN2(\IDinst/n8403 ), 
        .Q(\IDinst/n8405 ) );
  nnd2s1 \IDinst/U8455  ( .DIN1(\IDinst/n8402 ), .DIN2(n1162), 
        .Q(\IDinst/n8404 ) );
  nnd2s1 \IDinst/U8454  ( .DIN1(\IDinst/n8399 ), .DIN2(n1146), 
        .Q(\IDinst/n8403 ) );
  nnd2s1 \IDinst/U8453  ( .DIN1(\IDinst/n8401 ), .DIN2(\IDinst/n8400 ), 
        .Q(\IDinst/n8402 ) );
  nnd2s1 \IDinst/U8452  ( .DIN1(\IDinst/RegFile[19][26] ), .DIN2(n1090), 
        .Q(\IDinst/n8401 ) );
  nnd2s1 \IDinst/U8451  ( .DIN1(\IDinst/RegFile[18][26] ), .DIN2(n1048), 
        .Q(\IDinst/n8400 ) );
  nnd2s1 \IDinst/U8450  ( .DIN1(\IDinst/n8398 ), .DIN2(\IDinst/n8397 ), 
        .Q(\IDinst/n8399 ) );
  nnd2s1 \IDinst/U8449  ( .DIN1(\IDinst/RegFile[17][26] ), .DIN2(n1090), 
        .Q(\IDinst/n8398 ) );
  nnd2s1 \IDinst/U8448  ( .DIN1(\IDinst/RegFile[16][26] ), .DIN2(n1048), 
        .Q(\IDinst/n8397 ) );
  nnd2s1 \IDinst/U8447  ( .DIN1(\IDinst/n8395 ), .DIN2(\IDinst/n8394 ), 
        .Q(\IDinst/n8396 ) );
  nnd2s1 \IDinst/U8446  ( .DIN1(\IDinst/n8393 ), .DIN2(n644), 
        .Q(\IDinst/n8395 ) );
  nnd2s1 \IDinst/U8445  ( .DIN1(\IDinst/n8372 ), .DIN2(n672), 
        .Q(\IDinst/n8394 ) );
  nnd2s1 \IDinst/U8444  ( .DIN1(\IDinst/n8392 ), .DIN2(\IDinst/n8391 ), 
        .Q(\IDinst/n8393 ) );
  nnd2s1 \IDinst/U8443  ( .DIN1(\IDinst/n8390 ), .DIN2(n1190), 
        .Q(\IDinst/n8392 ) );
  nnd2s1 \IDinst/U8442  ( .DIN1(\IDinst/n8381 ), .DIN2(n1188), 
        .Q(\IDinst/n8391 ) );
  nnd2s1 \IDinst/U8441  ( .DIN1(\IDinst/n8389 ), .DIN2(\IDinst/n8388 ), 
        .Q(\IDinst/n8390 ) );
  nnd2s1 \IDinst/U8440  ( .DIN1(\IDinst/n8387 ), .DIN2(n1162), 
        .Q(\IDinst/n8389 ) );
  nnd2s1 \IDinst/U8439  ( .DIN1(\IDinst/n8384 ), .DIN2(n1146), 
        .Q(\IDinst/n8388 ) );
  nnd2s1 \IDinst/U8438  ( .DIN1(\IDinst/n8386 ), .DIN2(\IDinst/n8385 ), 
        .Q(\IDinst/n8387 ) );
  nnd2s1 \IDinst/U8437  ( .DIN1(\IDinst/RegFile[15][26] ), .DIN2(n1090), 
        .Q(\IDinst/n8386 ) );
  nnd2s1 \IDinst/U8436  ( .DIN1(\IDinst/RegFile[14][26] ), .DIN2(n1048), 
        .Q(\IDinst/n8385 ) );
  nnd2s1 \IDinst/U8435  ( .DIN1(\IDinst/n8383 ), .DIN2(\IDinst/n8382 ), 
        .Q(\IDinst/n8384 ) );
  nnd2s1 \IDinst/U8434  ( .DIN1(\IDinst/RegFile[13][26] ), .DIN2(n1090), 
        .Q(\IDinst/n8383 ) );
  nnd2s1 \IDinst/U8433  ( .DIN1(\IDinst/RegFile[12][26] ), .DIN2(n1048), 
        .Q(\IDinst/n8382 ) );
  nnd2s1 \IDinst/U8432  ( .DIN1(\IDinst/n8380 ), .DIN2(\IDinst/n8379 ), 
        .Q(\IDinst/n8381 ) );
  nnd2s1 \IDinst/U8431  ( .DIN1(\IDinst/n8378 ), .DIN2(n1162), 
        .Q(\IDinst/n8380 ) );
  nnd2s1 \IDinst/U8430  ( .DIN1(\IDinst/n8375 ), .DIN2(n1147), 
        .Q(\IDinst/n8379 ) );
  nnd2s1 \IDinst/U8429  ( .DIN1(\IDinst/n8377 ), .DIN2(\IDinst/n8376 ), 
        .Q(\IDinst/n8378 ) );
  nnd2s1 \IDinst/U8428  ( .DIN1(\IDinst/RegFile[11][26] ), .DIN2(n1091), 
        .Q(\IDinst/n8377 ) );
  nnd2s1 \IDinst/U8427  ( .DIN1(\IDinst/RegFile[10][26] ), .DIN2(n1048), 
        .Q(\IDinst/n8376 ) );
  nnd2s1 \IDinst/U8426  ( .DIN1(\IDinst/n8374 ), .DIN2(\IDinst/n8373 ), 
        .Q(\IDinst/n8375 ) );
  nnd2s1 \IDinst/U8425  ( .DIN1(\IDinst/RegFile[9][26] ), .DIN2(n1091), 
        .Q(\IDinst/n8374 ) );
  nnd2s1 \IDinst/U8424  ( .DIN1(\IDinst/RegFile[8][26] ), .DIN2(n1048), 
        .Q(\IDinst/n8373 ) );
  nnd2s1 \IDinst/U8423  ( .DIN1(\IDinst/n8371 ), .DIN2(\IDinst/n8370 ), 
        .Q(\IDinst/n8372 ) );
  nnd2s1 \IDinst/U8422  ( .DIN1(\IDinst/n8369 ), .DIN2(n1195), 
        .Q(\IDinst/n8371 ) );
  nnd2s1 \IDinst/U8421  ( .DIN1(\IDinst/n8360 ), .DIN2(n1188), 
        .Q(\IDinst/n8370 ) );
  nnd2s1 \IDinst/U8420  ( .DIN1(\IDinst/n8368 ), .DIN2(\IDinst/n8367 ), 
        .Q(\IDinst/n8369 ) );
  nnd2s1 \IDinst/U8419  ( .DIN1(\IDinst/n8366 ), .DIN2(n1162), 
        .Q(\IDinst/n8368 ) );
  nnd2s1 \IDinst/U8418  ( .DIN1(\IDinst/n8363 ), .DIN2(n1147), 
        .Q(\IDinst/n8367 ) );
  nnd2s1 \IDinst/U8417  ( .DIN1(\IDinst/n8365 ), .DIN2(\IDinst/n8364 ), 
        .Q(\IDinst/n8366 ) );
  nnd2s1 \IDinst/U8416  ( .DIN1(\IDinst/RegFile[7][26] ), .DIN2(n1091), 
        .Q(\IDinst/n8365 ) );
  nnd2s1 \IDinst/U8415  ( .DIN1(\IDinst/RegFile[6][26] ), .DIN2(n1048), 
        .Q(\IDinst/n8364 ) );
  nnd2s1 \IDinst/U8414  ( .DIN1(\IDinst/n8362 ), .DIN2(\IDinst/n8361 ), 
        .Q(\IDinst/n8363 ) );
  nnd2s1 \IDinst/U8413  ( .DIN1(\IDinst/RegFile[5][26] ), .DIN2(n1091), 
        .Q(\IDinst/n8362 ) );
  nnd2s1 \IDinst/U8412  ( .DIN1(\IDinst/RegFile[4][26] ), .DIN2(n1048), 
        .Q(\IDinst/n8361 ) );
  nnd2s1 \IDinst/U8411  ( .DIN1(\IDinst/n8359 ), .DIN2(\IDinst/n8358 ), 
        .Q(\IDinst/n8360 ) );
  nnd2s1 \IDinst/U8410  ( .DIN1(\IDinst/n8357 ), .DIN2(n1162), 
        .Q(\IDinst/n8359 ) );
  nnd2s1 \IDinst/U8409  ( .DIN1(\IDinst/n8354 ), .DIN2(n1147), 
        .Q(\IDinst/n8358 ) );
  nnd2s1 \IDinst/U8408  ( .DIN1(\IDinst/n8356 ), .DIN2(\IDinst/n8355 ), 
        .Q(\IDinst/n8357 ) );
  nnd2s1 \IDinst/U8407  ( .DIN1(\IDinst/RegFile[3][26] ), .DIN2(n1091), 
        .Q(\IDinst/n8356 ) );
  nnd2s1 \IDinst/U8406  ( .DIN1(\IDinst/RegFile[2][26] ), .DIN2(n1047), 
        .Q(\IDinst/n8355 ) );
  nnd2s1 \IDinst/U8405  ( .DIN1(\IDinst/n8353 ), .DIN2(\IDinst/n8352 ), 
        .Q(\IDinst/n8354 ) );
  nnd2s1 \IDinst/U8404  ( .DIN1(\IDinst/RegFile[1][26] ), .DIN2(n1091), 
        .Q(\IDinst/n8353 ) );
  nnd2s1 \IDinst/U8403  ( .DIN1(\IDinst/RegFile[0][26] ), .DIN2(n1047), 
        .Q(\IDinst/n8352 ) );
  nnd2s1 \IDinst/U8402  ( .DIN1(\IDinst/n8351 ), .DIN2(n539), 
        .Q(\IDinst/n5998 ) );
  nnd2s1 \IDinst/U8401  ( .DIN1(\IDinst/n8306 ), .DIN2(n635), 
        .Q(\IDinst/n5999 ) );
  nnd2s1 \IDinst/U8400  ( .DIN1(\IDinst/n8350 ), .DIN2(\IDinst/n8349 ), 
        .Q(\IDinst/n8351 ) );
  nnd2s1 \IDinst/U8399  ( .DIN1(\IDinst/n8348 ), .DIN2(n643), 
        .Q(\IDinst/n8350 ) );
  nnd2s1 \IDinst/U8398  ( .DIN1(\IDinst/n8327 ), .DIN2(n670), 
        .Q(\IDinst/n8349 ) );
  nnd2s1 \IDinst/U8397  ( .DIN1(\IDinst/n8347 ), .DIN2(\IDinst/n8346 ), 
        .Q(\IDinst/n8348 ) );
  nnd2s1 \IDinst/U8396  ( .DIN1(\IDinst/n8345 ), .DIN2(n1193), 
        .Q(\IDinst/n8347 ) );
  nnd2s1 \IDinst/U8395  ( .DIN1(\IDinst/n8336 ), .DIN2(n1188), 
        .Q(\IDinst/n8346 ) );
  nnd2s1 \IDinst/U8394  ( .DIN1(\IDinst/n8344 ), .DIN2(\IDinst/n8343 ), 
        .Q(\IDinst/n8345 ) );
  nnd2s1 \IDinst/U8393  ( .DIN1(\IDinst/n8342 ), .DIN2(n1162), 
        .Q(\IDinst/n8344 ) );
  nnd2s1 \IDinst/U8392  ( .DIN1(\IDinst/n8339 ), .DIN2(n1147), 
        .Q(\IDinst/n8343 ) );
  nnd2s1 \IDinst/U8391  ( .DIN1(\IDinst/n8341 ), .DIN2(\IDinst/n8340 ), 
        .Q(\IDinst/n8342 ) );
  nnd2s1 \IDinst/U8390  ( .DIN1(\IDinst/RegFile[31][25] ), .DIN2(n1091), 
        .Q(\IDinst/n8341 ) );
  nnd2s1 \IDinst/U8389  ( .DIN1(\IDinst/RegFile[30][25] ), .DIN2(n1047), 
        .Q(\IDinst/n8340 ) );
  nnd2s1 \IDinst/U8388  ( .DIN1(\IDinst/n8338 ), .DIN2(\IDinst/n8337 ), 
        .Q(\IDinst/n8339 ) );
  nnd2s1 \IDinst/U8387  ( .DIN1(\IDinst/RegFile[29][25] ), .DIN2(n1091), 
        .Q(\IDinst/n8338 ) );
  nnd2s1 \IDinst/U8386  ( .DIN1(\IDinst/RegFile[28][25] ), .DIN2(n1047), 
        .Q(\IDinst/n8337 ) );
  nnd2s1 \IDinst/U8385  ( .DIN1(\IDinst/n8335 ), .DIN2(\IDinst/n8334 ), 
        .Q(\IDinst/n8336 ) );
  nnd2s1 \IDinst/U8384  ( .DIN1(\IDinst/n8333 ), .DIN2(n1161), 
        .Q(\IDinst/n8335 ) );
  nnd2s1 \IDinst/U8383  ( .DIN1(\IDinst/n8330 ), .DIN2(n1147), 
        .Q(\IDinst/n8334 ) );
  nnd2s1 \IDinst/U8382  ( .DIN1(\IDinst/n8332 ), .DIN2(\IDinst/n8331 ), 
        .Q(\IDinst/n8333 ) );
  nnd2s1 \IDinst/U8381  ( .DIN1(\IDinst/RegFile[27][25] ), .DIN2(n1091), 
        .Q(\IDinst/n8332 ) );
  nnd2s1 \IDinst/U8380  ( .DIN1(\IDinst/RegFile[26][25] ), .DIN2(n1047), 
        .Q(\IDinst/n8331 ) );
  nnd2s1 \IDinst/U8379  ( .DIN1(\IDinst/n8329 ), .DIN2(\IDinst/n8328 ), 
        .Q(\IDinst/n8330 ) );
  nnd2s1 \IDinst/U8378  ( .DIN1(\IDinst/RegFile[25][25] ), .DIN2(n1092), 
        .Q(\IDinst/n8329 ) );
  nnd2s1 \IDinst/U8377  ( .DIN1(\IDinst/RegFile[24][25] ), .DIN2(n1047), 
        .Q(\IDinst/n8328 ) );
  nnd2s1 \IDinst/U8376  ( .DIN1(\IDinst/n8326 ), .DIN2(\IDinst/n8325 ), 
        .Q(\IDinst/n8327 ) );
  nnd2s1 \IDinst/U8375  ( .DIN1(\IDinst/n8324 ), .DIN2(n1192), 
        .Q(\IDinst/n8326 ) );
  nnd2s1 \IDinst/U8374  ( .DIN1(\IDinst/n8315 ), .DIN2(n1188), 
        .Q(\IDinst/n8325 ) );
  nnd2s1 \IDinst/U8373  ( .DIN1(\IDinst/n8323 ), .DIN2(\IDinst/n8322 ), 
        .Q(\IDinst/n8324 ) );
  nnd2s1 \IDinst/U8372  ( .DIN1(\IDinst/n8321 ), .DIN2(n1161), 
        .Q(\IDinst/n8323 ) );
  nnd2s1 \IDinst/U8371  ( .DIN1(\IDinst/n8318 ), .DIN2(n1147), 
        .Q(\IDinst/n8322 ) );
  nnd2s1 \IDinst/U8370  ( .DIN1(\IDinst/n8320 ), .DIN2(\IDinst/n8319 ), 
        .Q(\IDinst/n8321 ) );
  nnd2s1 \IDinst/U8369  ( .DIN1(\IDinst/RegFile[23][25] ), .DIN2(n1092), 
        .Q(\IDinst/n8320 ) );
  nnd2s1 \IDinst/U8368  ( .DIN1(\IDinst/RegFile[22][25] ), .DIN2(n1047), 
        .Q(\IDinst/n8319 ) );
  nnd2s1 \IDinst/U8367  ( .DIN1(\IDinst/n8317 ), .DIN2(\IDinst/n8316 ), 
        .Q(\IDinst/n8318 ) );
  nnd2s1 \IDinst/U8366  ( .DIN1(\IDinst/RegFile[21][25] ), .DIN2(n1092), 
        .Q(\IDinst/n8317 ) );
  nnd2s1 \IDinst/U8365  ( .DIN1(\IDinst/RegFile[20][25] ), .DIN2(n1047), 
        .Q(\IDinst/n8316 ) );
  nnd2s1 \IDinst/U8364  ( .DIN1(\IDinst/n8314 ), .DIN2(\IDinst/n8313 ), 
        .Q(\IDinst/n8315 ) );
  nnd2s1 \IDinst/U8363  ( .DIN1(\IDinst/n8312 ), .DIN2(n1161), 
        .Q(\IDinst/n8314 ) );
  nnd2s1 \IDinst/U8362  ( .DIN1(\IDinst/n8309 ), .DIN2(n1147), 
        .Q(\IDinst/n8313 ) );
  nnd2s1 \IDinst/U8361  ( .DIN1(\IDinst/n8311 ), .DIN2(\IDinst/n8310 ), 
        .Q(\IDinst/n8312 ) );
  nnd2s1 \IDinst/U8360  ( .DIN1(\IDinst/RegFile[19][25] ), .DIN2(n1092), 
        .Q(\IDinst/n8311 ) );
  nnd2s1 \IDinst/U8359  ( .DIN1(\IDinst/RegFile[18][25] ), .DIN2(n1047), 
        .Q(\IDinst/n8310 ) );
  nnd2s1 \IDinst/U8358  ( .DIN1(\IDinst/n8308 ), .DIN2(\IDinst/n8307 ), 
        .Q(\IDinst/n8309 ) );
  nnd2s1 \IDinst/U8357  ( .DIN1(\IDinst/RegFile[17][25] ), .DIN2(n1092), 
        .Q(\IDinst/n8308 ) );
  nnd2s1 \IDinst/U8356  ( .DIN1(\IDinst/RegFile[16][25] ), .DIN2(n1047), 
        .Q(\IDinst/n8307 ) );
  nnd2s1 \IDinst/U8355  ( .DIN1(\IDinst/n8305 ), .DIN2(\IDinst/n8304 ), 
        .Q(\IDinst/n8306 ) );
  nnd2s1 \IDinst/U8354  ( .DIN1(\IDinst/n8303 ), .DIN2(n642), 
        .Q(\IDinst/n8305 ) );
  nnd2s1 \IDinst/U8353  ( .DIN1(\IDinst/n8282 ), .DIN2(n673), 
        .Q(\IDinst/n8304 ) );
  nnd2s1 \IDinst/U8352  ( .DIN1(\IDinst/n8302 ), .DIN2(\IDinst/n8301 ), 
        .Q(\IDinst/n8303 ) );
  nnd2s1 \IDinst/U8351  ( .DIN1(\IDinst/n8300 ), .DIN2(n1195), 
        .Q(\IDinst/n8302 ) );
  nnd2s1 \IDinst/U8350  ( .DIN1(\IDinst/n8291 ), .DIN2(n1188), 
        .Q(\IDinst/n8301 ) );
  nnd2s1 \IDinst/U8349  ( .DIN1(\IDinst/n8299 ), .DIN2(\IDinst/n8298 ), 
        .Q(\IDinst/n8300 ) );
  nnd2s1 \IDinst/U8348  ( .DIN1(\IDinst/n8297 ), .DIN2(n1161), 
        .Q(\IDinst/n8299 ) );
  nnd2s1 \IDinst/U8347  ( .DIN1(\IDinst/n8294 ), .DIN2(n1147), 
        .Q(\IDinst/n8298 ) );
  nnd2s1 \IDinst/U8346  ( .DIN1(\IDinst/n8296 ), .DIN2(\IDinst/n8295 ), 
        .Q(\IDinst/n8297 ) );
  nnd2s1 \IDinst/U8345  ( .DIN1(\IDinst/RegFile[15][25] ), .DIN2(n1092), 
        .Q(\IDinst/n8296 ) );
  nnd2s1 \IDinst/U8344  ( .DIN1(\IDinst/RegFile[14][25] ), .DIN2(n1047), 
        .Q(\IDinst/n8295 ) );
  nnd2s1 \IDinst/U8343  ( .DIN1(\IDinst/n8293 ), .DIN2(\IDinst/n8292 ), 
        .Q(\IDinst/n8294 ) );
  nnd2s1 \IDinst/U8342  ( .DIN1(\IDinst/RegFile[13][25] ), .DIN2(n1092), 
        .Q(\IDinst/n8293 ) );
  nnd2s1 \IDinst/U8341  ( .DIN1(\IDinst/RegFile[12][25] ), .DIN2(n1047), 
        .Q(\IDinst/n8292 ) );
  nnd2s1 \IDinst/U8340  ( .DIN1(\IDinst/n8290 ), .DIN2(\IDinst/n8289 ), 
        .Q(\IDinst/n8291 ) );
  nnd2s1 \IDinst/U8339  ( .DIN1(\IDinst/n8288 ), .DIN2(n1161), 
        .Q(\IDinst/n8290 ) );
  nnd2s1 \IDinst/U8338  ( .DIN1(\IDinst/n8285 ), .DIN2(n1147), 
        .Q(\IDinst/n8289 ) );
  nnd2s1 \IDinst/U8337  ( .DIN1(\IDinst/n8287 ), .DIN2(\IDinst/n8286 ), 
        .Q(\IDinst/n8288 ) );
  nnd2s1 \IDinst/U8336  ( .DIN1(\IDinst/RegFile[11][25] ), .DIN2(n1092), 
        .Q(\IDinst/n8287 ) );
  nnd2s1 \IDinst/U8335  ( .DIN1(\IDinst/RegFile[10][25] ), .DIN2(n1047), 
        .Q(\IDinst/n8286 ) );
  nnd2s1 \IDinst/U8334  ( .DIN1(\IDinst/n8284 ), .DIN2(\IDinst/n8283 ), 
        .Q(\IDinst/n8285 ) );
  nnd2s1 \IDinst/U8333  ( .DIN1(\IDinst/RegFile[9][25] ), .DIN2(n1092), 
        .Q(\IDinst/n8284 ) );
  nnd2s1 \IDinst/U8332  ( .DIN1(\IDinst/RegFile[8][25] ), .DIN2(n1046), 
        .Q(\IDinst/n8283 ) );
  nnd2s1 \IDinst/U8331  ( .DIN1(\IDinst/n8281 ), .DIN2(\IDinst/n8280 ), 
        .Q(\IDinst/n8282 ) );
  nnd2s1 \IDinst/U8330  ( .DIN1(\IDinst/n8279 ), .DIN2(n1194), 
        .Q(\IDinst/n8281 ) );
  nnd2s1 \IDinst/U8329  ( .DIN1(\IDinst/n8270 ), .DIN2(n1188), 
        .Q(\IDinst/n8280 ) );
  nnd2s1 \IDinst/U8328  ( .DIN1(\IDinst/n8278 ), .DIN2(\IDinst/n8277 ), 
        .Q(\IDinst/n8279 ) );
  nnd2s1 \IDinst/U8327  ( .DIN1(\IDinst/n8276 ), .DIN2(n1161), 
        .Q(\IDinst/n8278 ) );
  nnd2s1 \IDinst/U8326  ( .DIN1(\IDinst/n8273 ), .DIN2(n1147), 
        .Q(\IDinst/n8277 ) );
  nnd2s1 \IDinst/U8325  ( .DIN1(\IDinst/n8275 ), .DIN2(\IDinst/n8274 ), 
        .Q(\IDinst/n8276 ) );
  nnd2s1 \IDinst/U8324  ( .DIN1(\IDinst/RegFile[7][25] ), .DIN2(n1093), 
        .Q(\IDinst/n8275 ) );
  nnd2s1 \IDinst/U8323  ( .DIN1(\IDinst/RegFile[6][25] ), .DIN2(n1046), 
        .Q(\IDinst/n8274 ) );
  nnd2s1 \IDinst/U8322  ( .DIN1(\IDinst/n8272 ), .DIN2(\IDinst/n8271 ), 
        .Q(\IDinst/n8273 ) );
  nnd2s1 \IDinst/U8321  ( .DIN1(\IDinst/RegFile[5][25] ), .DIN2(n1093), 
        .Q(\IDinst/n8272 ) );
  nnd2s1 \IDinst/U8320  ( .DIN1(\IDinst/RegFile[4][25] ), .DIN2(n1046), 
        .Q(\IDinst/n8271 ) );
  nnd2s1 \IDinst/U8319  ( .DIN1(\IDinst/n8269 ), .DIN2(\IDinst/n8268 ), 
        .Q(\IDinst/n8270 ) );
  nnd2s1 \IDinst/U8318  ( .DIN1(\IDinst/n8267 ), .DIN2(n1161), 
        .Q(\IDinst/n8269 ) );
  nnd2s1 \IDinst/U8317  ( .DIN1(\IDinst/n8264 ), .DIN2(n1147), 
        .Q(\IDinst/n8268 ) );
  nnd2s1 \IDinst/U8316  ( .DIN1(\IDinst/n8266 ), .DIN2(\IDinst/n8265 ), 
        .Q(\IDinst/n8267 ) );
  nnd2s1 \IDinst/U8315  ( .DIN1(\IDinst/RegFile[3][25] ), .DIN2(n1093), 
        .Q(\IDinst/n8266 ) );
  nnd2s1 \IDinst/U8314  ( .DIN1(\IDinst/RegFile[2][25] ), .DIN2(n1046), 
        .Q(\IDinst/n8265 ) );
  nnd2s1 \IDinst/U8313  ( .DIN1(\IDinst/n8263 ), .DIN2(\IDinst/n8262 ), 
        .Q(\IDinst/n8264 ) );
  nnd2s1 \IDinst/U8312  ( .DIN1(\IDinst/RegFile[1][25] ), .DIN2(n1093), 
        .Q(\IDinst/n8263 ) );
  nnd2s1 \IDinst/U8311  ( .DIN1(\IDinst/RegFile[0][25] ), .DIN2(n1046), 
        .Q(\IDinst/n8262 ) );
  nnd2s1 \IDinst/U8310  ( .DIN1(\IDinst/n8261 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n5996 ) );
  nnd2s1 \IDinst/U8309  ( .DIN1(\IDinst/n8216 ), .DIN2(n636), 
        .Q(\IDinst/n5997 ) );
  nnd2s1 \IDinst/U8308  ( .DIN1(\IDinst/n8260 ), .DIN2(\IDinst/n8259 ), 
        .Q(\IDinst/n8261 ) );
  nnd2s1 \IDinst/U8307  ( .DIN1(\IDinst/n8258 ), .DIN2(n641), 
        .Q(\IDinst/n8260 ) );
  nnd2s1 \IDinst/U8306  ( .DIN1(\IDinst/n8237 ), .DIN2(n671), 
        .Q(\IDinst/n8259 ) );
  nnd2s1 \IDinst/U8305  ( .DIN1(\IDinst/n8257 ), .DIN2(\IDinst/n8256 ), 
        .Q(\IDinst/n8258 ) );
  nnd2s1 \IDinst/U8304  ( .DIN1(\IDinst/n8255 ), .DIN2(n1197), 
        .Q(\IDinst/n8257 ) );
  nnd2s1 \IDinst/U8303  ( .DIN1(\IDinst/n8246 ), .DIN2(n1188), 
        .Q(\IDinst/n8256 ) );
  nnd2s1 \IDinst/U8302  ( .DIN1(\IDinst/n8254 ), .DIN2(\IDinst/n8253 ), 
        .Q(\IDinst/n8255 ) );
  nnd2s1 \IDinst/U8301  ( .DIN1(\IDinst/n8252 ), .DIN2(n1161), 
        .Q(\IDinst/n8254 ) );
  nnd2s1 \IDinst/U8300  ( .DIN1(\IDinst/n8249 ), .DIN2(n1147), 
        .Q(\IDinst/n8253 ) );
  nnd2s1 \IDinst/U8299  ( .DIN1(\IDinst/n8251 ), .DIN2(\IDinst/n8250 ), 
        .Q(\IDinst/n8252 ) );
  nnd2s1 \IDinst/U8298  ( .DIN1(\IDinst/RegFile[31][24] ), .DIN2(n1093), 
        .Q(\IDinst/n8251 ) );
  nnd2s1 \IDinst/U8297  ( .DIN1(\IDinst/RegFile[30][24] ), .DIN2(n1046), 
        .Q(\IDinst/n8250 ) );
  nnd2s1 \IDinst/U8296  ( .DIN1(\IDinst/n8248 ), .DIN2(\IDinst/n8247 ), 
        .Q(\IDinst/n8249 ) );
  nnd2s1 \IDinst/U8295  ( .DIN1(\IDinst/RegFile[29][24] ), .DIN2(n1093), 
        .Q(\IDinst/n8248 ) );
  nnd2s1 \IDinst/U8294  ( .DIN1(\IDinst/RegFile[28][24] ), .DIN2(n1046), 
        .Q(\IDinst/n8247 ) );
  nnd2s1 \IDinst/U8293  ( .DIN1(\IDinst/n8245 ), .DIN2(\IDinst/n8244 ), 
        .Q(\IDinst/n8246 ) );
  nnd2s1 \IDinst/U8292  ( .DIN1(\IDinst/n8243 ), .DIN2(n1161), 
        .Q(\IDinst/n8245 ) );
  nnd2s1 \IDinst/U8291  ( .DIN1(\IDinst/n8240 ), .DIN2(n1147), 
        .Q(\IDinst/n8244 ) );
  nnd2s1 \IDinst/U8290  ( .DIN1(\IDinst/n8242 ), .DIN2(\IDinst/n8241 ), 
        .Q(\IDinst/n8243 ) );
  nnd2s1 \IDinst/U8289  ( .DIN1(\IDinst/RegFile[27][24] ), .DIN2(n1093), 
        .Q(\IDinst/n8242 ) );
  nnd2s1 \IDinst/U8288  ( .DIN1(\IDinst/RegFile[26][24] ), .DIN2(n1046), 
        .Q(\IDinst/n8241 ) );
  nnd2s1 \IDinst/U8287  ( .DIN1(\IDinst/n8239 ), .DIN2(\IDinst/n8238 ), 
        .Q(\IDinst/n8240 ) );
  nnd2s1 \IDinst/U8286  ( .DIN1(\IDinst/RegFile[25][24] ), .DIN2(n1093), 
        .Q(\IDinst/n8239 ) );
  nnd2s1 \IDinst/U8285  ( .DIN1(\IDinst/RegFile[24][24] ), .DIN2(n1046), 
        .Q(\IDinst/n8238 ) );
  nnd2s1 \IDinst/U8284  ( .DIN1(\IDinst/n8236 ), .DIN2(\IDinst/n8235 ), 
        .Q(\IDinst/n8237 ) );
  nnd2s1 \IDinst/U8283  ( .DIN1(\IDinst/n8234 ), .DIN2(n1190), 
        .Q(\IDinst/n8236 ) );
  nnd2s1 \IDinst/U8282  ( .DIN1(\IDinst/n8225 ), .DIN2(n1188), 
        .Q(\IDinst/n8235 ) );
  nnd2s1 \IDinst/U8281  ( .DIN1(\IDinst/n8233 ), .DIN2(\IDinst/n8232 ), 
        .Q(\IDinst/n8234 ) );
  nnd2s1 \IDinst/U8280  ( .DIN1(\IDinst/n8231 ), .DIN2(n1160), 
        .Q(\IDinst/n8233 ) );
  nnd2s1 \IDinst/U8279  ( .DIN1(\IDinst/n8228 ), .DIN2(n1148), 
        .Q(\IDinst/n8232 ) );
  nnd2s1 \IDinst/U8278  ( .DIN1(\IDinst/n8230 ), .DIN2(\IDinst/n8229 ), 
        .Q(\IDinst/n8231 ) );
  nnd2s1 \IDinst/U8277  ( .DIN1(\IDinst/RegFile[23][24] ), .DIN2(n1093), 
        .Q(\IDinst/n8230 ) );
  nnd2s1 \IDinst/U8276  ( .DIN1(\IDinst/RegFile[22][24] ), .DIN2(n1046), 
        .Q(\IDinst/n8229 ) );
  nnd2s1 \IDinst/U8275  ( .DIN1(\IDinst/n8227 ), .DIN2(\IDinst/n8226 ), 
        .Q(\IDinst/n8228 ) );
  nnd2s1 \IDinst/U8274  ( .DIN1(\IDinst/RegFile[21][24] ), .DIN2(n1094), 
        .Q(\IDinst/n8227 ) );
  nnd2s1 \IDinst/U8273  ( .DIN1(\IDinst/RegFile[20][24] ), .DIN2(n1046), 
        .Q(\IDinst/n8226 ) );
  nnd2s1 \IDinst/U8272  ( .DIN1(\IDinst/n8224 ), .DIN2(\IDinst/n8223 ), 
        .Q(\IDinst/n8225 ) );
  nnd2s1 \IDinst/U8271  ( .DIN1(\IDinst/n8222 ), .DIN2(n1160), 
        .Q(\IDinst/n8224 ) );
  nnd2s1 \IDinst/U8270  ( .DIN1(\IDinst/n8219 ), .DIN2(n1148), 
        .Q(\IDinst/n8223 ) );
  nnd2s1 \IDinst/U8269  ( .DIN1(\IDinst/n8221 ), .DIN2(\IDinst/n8220 ), 
        .Q(\IDinst/n8222 ) );
  nnd2s1 \IDinst/U8268  ( .DIN1(\IDinst/RegFile[19][24] ), .DIN2(n1094), 
        .Q(\IDinst/n8221 ) );
  nnd2s1 \IDinst/U8267  ( .DIN1(\IDinst/RegFile[18][24] ), .DIN2(n1046), 
        .Q(\IDinst/n8220 ) );
  nnd2s1 \IDinst/U8266  ( .DIN1(\IDinst/n8218 ), .DIN2(\IDinst/n8217 ), 
        .Q(\IDinst/n8219 ) );
  nnd2s1 \IDinst/U8265  ( .DIN1(\IDinst/RegFile[17][24] ), .DIN2(n1094), 
        .Q(\IDinst/n8218 ) );
  nnd2s1 \IDinst/U8264  ( .DIN1(\IDinst/RegFile[16][24] ), .DIN2(n1046), 
        .Q(\IDinst/n8217 ) );
  nnd2s1 \IDinst/U8263  ( .DIN1(\IDinst/n8215 ), .DIN2(\IDinst/n8214 ), 
        .Q(\IDinst/n8216 ) );
  nnd2s1 \IDinst/U8262  ( .DIN1(\IDinst/n8213 ), .DIN2(n644), 
        .Q(\IDinst/n8215 ) );
  nnd2s1 \IDinst/U8261  ( .DIN1(\IDinst/n8192 ), .DIN2(n672), 
        .Q(\IDinst/n8214 ) );
  nnd2s1 \IDinst/U8260  ( .DIN1(\IDinst/n8212 ), .DIN2(\IDinst/n8211 ), 
        .Q(\IDinst/n8213 ) );
  nnd2s1 \IDinst/U8259  ( .DIN1(\IDinst/n8210 ), .DIN2(n1190), 
        .Q(\IDinst/n8212 ) );
  nnd2s1 \IDinst/U8258  ( .DIN1(\IDinst/n8201 ), .DIN2(n1188), 
        .Q(\IDinst/n8211 ) );
  nnd2s1 \IDinst/U8257  ( .DIN1(\IDinst/n8209 ), .DIN2(\IDinst/n8208 ), 
        .Q(\IDinst/n8210 ) );
  nnd2s1 \IDinst/U8256  ( .DIN1(\IDinst/n8207 ), .DIN2(n1160), 
        .Q(\IDinst/n8209 ) );
  nnd2s1 \IDinst/U8255  ( .DIN1(\IDinst/n8204 ), .DIN2(n1148), 
        .Q(\IDinst/n8208 ) );
  nnd2s1 \IDinst/U8254  ( .DIN1(\IDinst/n8206 ), .DIN2(\IDinst/n8205 ), 
        .Q(\IDinst/n8207 ) );
  nnd2s1 \IDinst/U8253  ( .DIN1(\IDinst/RegFile[15][24] ), .DIN2(n1094), 
        .Q(\IDinst/n8206 ) );
  nnd2s1 \IDinst/U8252  ( .DIN1(\IDinst/RegFile[14][24] ), .DIN2(n1045), 
        .Q(\IDinst/n8205 ) );
  nnd2s1 \IDinst/U8251  ( .DIN1(\IDinst/n8203 ), .DIN2(\IDinst/n8202 ), 
        .Q(\IDinst/n8204 ) );
  nnd2s1 \IDinst/U8250  ( .DIN1(\IDinst/RegFile[13][24] ), .DIN2(n1094), 
        .Q(\IDinst/n8203 ) );
  nnd2s1 \IDinst/U8249  ( .DIN1(\IDinst/RegFile[12][24] ), .DIN2(n1045), 
        .Q(\IDinst/n8202 ) );
  nnd2s1 \IDinst/U8248  ( .DIN1(\IDinst/n8200 ), .DIN2(\IDinst/n8199 ), 
        .Q(\IDinst/n8201 ) );
  nnd2s1 \IDinst/U8247  ( .DIN1(\IDinst/n8198 ), .DIN2(n1160), 
        .Q(\IDinst/n8200 ) );
  nnd2s1 \IDinst/U8246  ( .DIN1(\IDinst/n8195 ), .DIN2(n1148), 
        .Q(\IDinst/n8199 ) );
  nnd2s1 \IDinst/U8245  ( .DIN1(\IDinst/n8197 ), .DIN2(\IDinst/n8196 ), 
        .Q(\IDinst/n8198 ) );
  nnd2s1 \IDinst/U8244  ( .DIN1(\IDinst/RegFile[11][24] ), .DIN2(n1094), 
        .Q(\IDinst/n8197 ) );
  nnd2s1 \IDinst/U8243  ( .DIN1(\IDinst/RegFile[10][24] ), .DIN2(n1045), 
        .Q(\IDinst/n8196 ) );
  nnd2s1 \IDinst/U8242  ( .DIN1(\IDinst/n8194 ), .DIN2(\IDinst/n8193 ), 
        .Q(\IDinst/n8195 ) );
  nnd2s1 \IDinst/U8241  ( .DIN1(\IDinst/RegFile[9][24] ), .DIN2(n1094), 
        .Q(\IDinst/n8194 ) );
  nnd2s1 \IDinst/U8240  ( .DIN1(\IDinst/RegFile[8][24] ), .DIN2(n1045), 
        .Q(\IDinst/n8193 ) );
  nnd2s1 \IDinst/U8239  ( .DIN1(\IDinst/n8191 ), .DIN2(\IDinst/n8190 ), 
        .Q(\IDinst/n8192 ) );
  nnd2s1 \IDinst/U8238  ( .DIN1(\IDinst/n8189 ), .DIN2(n1190), 
        .Q(\IDinst/n8191 ) );
  nnd2s1 \IDinst/U8237  ( .DIN1(\IDinst/n8180 ), .DIN2(n1188), 
        .Q(\IDinst/n8190 ) );
  nnd2s1 \IDinst/U8236  ( .DIN1(\IDinst/n8188 ), .DIN2(\IDinst/n8187 ), 
        .Q(\IDinst/n8189 ) );
  nnd2s1 \IDinst/U8235  ( .DIN1(\IDinst/n8186 ), .DIN2(n1160), 
        .Q(\IDinst/n8188 ) );
  nnd2s1 \IDinst/U8234  ( .DIN1(\IDinst/n8183 ), .DIN2(n1148), 
        .Q(\IDinst/n8187 ) );
  nnd2s1 \IDinst/U8233  ( .DIN1(\IDinst/n8185 ), .DIN2(\IDinst/n8184 ), 
        .Q(\IDinst/n8186 ) );
  nnd2s1 \IDinst/U8232  ( .DIN1(\IDinst/RegFile[7][24] ), .DIN2(n1094), 
        .Q(\IDinst/n8185 ) );
  nnd2s1 \IDinst/U8231  ( .DIN1(\IDinst/RegFile[6][24] ), .DIN2(n1045), 
        .Q(\IDinst/n8184 ) );
  nnd2s1 \IDinst/U8230  ( .DIN1(\IDinst/n8182 ), .DIN2(\IDinst/n8181 ), 
        .Q(\IDinst/n8183 ) );
  nnd2s1 \IDinst/U8229  ( .DIN1(\IDinst/RegFile[5][24] ), .DIN2(n1094), 
        .Q(\IDinst/n8182 ) );
  nnd2s1 \IDinst/U8228  ( .DIN1(\IDinst/RegFile[4][24] ), .DIN2(n1045), 
        .Q(\IDinst/n8181 ) );
  nnd2s1 \IDinst/U8227  ( .DIN1(\IDinst/n8179 ), .DIN2(\IDinst/n8178 ), 
        .Q(\IDinst/n8180 ) );
  nnd2s1 \IDinst/U8226  ( .DIN1(\IDinst/n8177 ), .DIN2(n1160), 
        .Q(\IDinst/n8179 ) );
  nnd2s1 \IDinst/U8225  ( .DIN1(\IDinst/n8174 ), .DIN2(n1148), 
        .Q(\IDinst/n8178 ) );
  nnd2s1 \IDinst/U8224  ( .DIN1(\IDinst/n8176 ), .DIN2(\IDinst/n8175 ), 
        .Q(\IDinst/n8177 ) );
  nnd2s1 \IDinst/U8223  ( .DIN1(\IDinst/RegFile[3][24] ), .DIN2(n1095), 
        .Q(\IDinst/n8176 ) );
  nnd2s1 \IDinst/U8222  ( .DIN1(\IDinst/RegFile[2][24] ), .DIN2(n1045), 
        .Q(\IDinst/n8175 ) );
  nnd2s1 \IDinst/U8221  ( .DIN1(\IDinst/n8173 ), .DIN2(\IDinst/n8172 ), 
        .Q(\IDinst/n8174 ) );
  nnd2s1 \IDinst/U8220  ( .DIN1(\IDinst/RegFile[1][24] ), .DIN2(n1095), 
        .Q(\IDinst/n8173 ) );
  nnd2s1 \IDinst/U8219  ( .DIN1(\IDinst/RegFile[0][24] ), .DIN2(n1050), 
        .Q(\IDinst/n8172 ) );
  nnd2s1 \IDinst/U8218  ( .DIN1(\IDinst/n8171 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n5994 ) );
  nnd2s1 \IDinst/U8217  ( .DIN1(\IDinst/n8126 ), .DIN2(n635), 
        .Q(\IDinst/n5995 ) );
  nnd2s1 \IDinst/U8216  ( .DIN1(\IDinst/n8170 ), .DIN2(\IDinst/n8169 ), 
        .Q(\IDinst/n8171 ) );
  nnd2s1 \IDinst/U8215  ( .DIN1(\IDinst/n8168 ), .DIN2(n643), 
        .Q(\IDinst/n8170 ) );
  nnd2s1 \IDinst/U8214  ( .DIN1(\IDinst/n8147 ), .DIN2(n670), 
        .Q(\IDinst/n8169 ) );
  nnd2s1 \IDinst/U8213  ( .DIN1(\IDinst/n8167 ), .DIN2(\IDinst/n8166 ), 
        .Q(\IDinst/n8168 ) );
  nnd2s1 \IDinst/U8212  ( .DIN1(\IDinst/n8165 ), .DIN2(n1190), 
        .Q(\IDinst/n8167 ) );
  nnd2s1 \IDinst/U8211  ( .DIN1(\IDinst/n8156 ), .DIN2(n1187), 
        .Q(\IDinst/n8166 ) );
  nnd2s1 \IDinst/U8210  ( .DIN1(\IDinst/n8164 ), .DIN2(\IDinst/n8163 ), 
        .Q(\IDinst/n8165 ) );
  nnd2s1 \IDinst/U8209  ( .DIN1(\IDinst/n8162 ), .DIN2(n1160), 
        .Q(\IDinst/n8164 ) );
  nnd2s1 \IDinst/U8208  ( .DIN1(\IDinst/n8159 ), .DIN2(n1148), 
        .Q(\IDinst/n8163 ) );
  nnd2s1 \IDinst/U8207  ( .DIN1(\IDinst/n8161 ), .DIN2(\IDinst/n8160 ), 
        .Q(\IDinst/n8162 ) );
  nnd2s1 \IDinst/U8206  ( .DIN1(\IDinst/RegFile[31][23] ), .DIN2(n1095), 
        .Q(\IDinst/n8161 ) );
  nnd2s1 \IDinst/U8205  ( .DIN1(\IDinst/RegFile[30][23] ), .DIN2(n1131), 
        .Q(\IDinst/n8160 ) );
  nnd2s1 \IDinst/U8204  ( .DIN1(\IDinst/n8158 ), .DIN2(\IDinst/n8157 ), 
        .Q(\IDinst/n8159 ) );
  nnd2s1 \IDinst/U8203  ( .DIN1(\IDinst/RegFile[29][23] ), .DIN2(n1095), 
        .Q(\IDinst/n8158 ) );
  nnd2s1 \IDinst/U8202  ( .DIN1(\IDinst/RegFile[28][23] ), .DIN2(n1064), 
        .Q(\IDinst/n8157 ) );
  nnd2s1 \IDinst/U8201  ( .DIN1(\IDinst/n8155 ), .DIN2(\IDinst/n8154 ), 
        .Q(\IDinst/n8156 ) );
  nnd2s1 \IDinst/U8200  ( .DIN1(\IDinst/n8153 ), .DIN2(n1160), 
        .Q(\IDinst/n8155 ) );
  nnd2s1 \IDinst/U8199  ( .DIN1(\IDinst/n8150 ), .DIN2(n1148), 
        .Q(\IDinst/n8154 ) );
  nnd2s1 \IDinst/U8198  ( .DIN1(\IDinst/n8152 ), .DIN2(\IDinst/n8151 ), 
        .Q(\IDinst/n8153 ) );
  nnd2s1 \IDinst/U8197  ( .DIN1(\IDinst/RegFile[27][23] ), .DIN2(n1095), 
        .Q(\IDinst/n8152 ) );
  nnd2s1 \IDinst/U8196  ( .DIN1(\IDinst/RegFile[26][23] ), .DIN2(n1064), 
        .Q(\IDinst/n8151 ) );
  nnd2s1 \IDinst/U8195  ( .DIN1(\IDinst/n8149 ), .DIN2(\IDinst/n8148 ), 
        .Q(\IDinst/n8150 ) );
  nnd2s1 \IDinst/U8194  ( .DIN1(\IDinst/RegFile[25][23] ), .DIN2(n1095), 
        .Q(\IDinst/n8149 ) );
  nnd2s1 \IDinst/U8193  ( .DIN1(\IDinst/RegFile[24][23] ), .DIN2(n1064), 
        .Q(\IDinst/n8148 ) );
  nnd2s1 \IDinst/U8192  ( .DIN1(\IDinst/n8146 ), .DIN2(\IDinst/n8145 ), 
        .Q(\IDinst/n8147 ) );
  nnd2s1 \IDinst/U8191  ( .DIN1(\IDinst/n8144 ), .DIN2(n1190), 
        .Q(\IDinst/n8146 ) );
  nnd2s1 \IDinst/U8190  ( .DIN1(\IDinst/n8135 ), .DIN2(n1187), 
        .Q(\IDinst/n8145 ) );
  nnd2s1 \IDinst/U8189  ( .DIN1(\IDinst/n8143 ), .DIN2(\IDinst/n8142 ), 
        .Q(\IDinst/n8144 ) );
  nnd2s1 \IDinst/U8188  ( .DIN1(\IDinst/n8141 ), .DIN2(n1160), 
        .Q(\IDinst/n8143 ) );
  nnd2s1 \IDinst/U8187  ( .DIN1(\IDinst/n8138 ), .DIN2(n1148), 
        .Q(\IDinst/n8142 ) );
  nnd2s1 \IDinst/U8186  ( .DIN1(\IDinst/n8140 ), .DIN2(\IDinst/n8139 ), 
        .Q(\IDinst/n8141 ) );
  nnd2s1 \IDinst/U8185  ( .DIN1(\IDinst/RegFile[23][23] ), .DIN2(n1095), 
        .Q(\IDinst/n8140 ) );
  nnd2s1 \IDinst/U8184  ( .DIN1(\IDinst/RegFile[22][23] ), .DIN2(n1064), 
        .Q(\IDinst/n8139 ) );
  nnd2s1 \IDinst/U8183  ( .DIN1(\IDinst/n8137 ), .DIN2(\IDinst/n8136 ), 
        .Q(\IDinst/n8138 ) );
  nnd2s1 \IDinst/U8182  ( .DIN1(\IDinst/RegFile[21][23] ), .DIN2(n1095), 
        .Q(\IDinst/n8137 ) );
  nnd2s1 \IDinst/U8181  ( .DIN1(\IDinst/RegFile[20][23] ), .DIN2(n1064), 
        .Q(\IDinst/n8136 ) );
  nnd2s1 \IDinst/U8180  ( .DIN1(\IDinst/n8134 ), .DIN2(\IDinst/n8133 ), 
        .Q(\IDinst/n8135 ) );
  nnd2s1 \IDinst/U8179  ( .DIN1(\IDinst/n8132 ), .DIN2(n1159), 
        .Q(\IDinst/n8134 ) );
  nnd2s1 \IDinst/U8178  ( .DIN1(\IDinst/n8129 ), .DIN2(n1148), 
        .Q(\IDinst/n8133 ) );
  nnd2s1 \IDinst/U8177  ( .DIN1(\IDinst/n8131 ), .DIN2(\IDinst/n8130 ), 
        .Q(\IDinst/n8132 ) );
  nnd2s1 \IDinst/U8176  ( .DIN1(\IDinst/RegFile[19][23] ), .DIN2(n1095), 
        .Q(\IDinst/n8131 ) );
  nnd2s1 \IDinst/U8175  ( .DIN1(\IDinst/RegFile[18][23] ), .DIN2(n1064), 
        .Q(\IDinst/n8130 ) );
  nnd2s1 \IDinst/U8174  ( .DIN1(\IDinst/n8128 ), .DIN2(\IDinst/n8127 ), 
        .Q(\IDinst/n8129 ) );
  nnd2s1 \IDinst/U8173  ( .DIN1(\IDinst/RegFile[17][23] ), .DIN2(n1096), 
        .Q(\IDinst/n8128 ) );
  nnd2s1 \IDinst/U8172  ( .DIN1(\IDinst/RegFile[16][23] ), .DIN2(n1064), 
        .Q(\IDinst/n8127 ) );
  nnd2s1 \IDinst/U8171  ( .DIN1(\IDinst/n8125 ), .DIN2(\IDinst/n8124 ), 
        .Q(\IDinst/n8126 ) );
  nnd2s1 \IDinst/U8170  ( .DIN1(\IDinst/n8123 ), .DIN2(n642), 
        .Q(\IDinst/n8125 ) );
  nnd2s1 \IDinst/U8169  ( .DIN1(\IDinst/n8102 ), .DIN2(n673), 
        .Q(\IDinst/n8124 ) );
  nnd2s1 \IDinst/U8168  ( .DIN1(\IDinst/n8122 ), .DIN2(\IDinst/n8121 ), 
        .Q(\IDinst/n8123 ) );
  nnd2s1 \IDinst/U8167  ( .DIN1(\IDinst/n8120 ), .DIN2(n1190), 
        .Q(\IDinst/n8122 ) );
  nnd2s1 \IDinst/U8166  ( .DIN1(\IDinst/n8111 ), .DIN2(n1187), 
        .Q(\IDinst/n8121 ) );
  nnd2s1 \IDinst/U8165  ( .DIN1(\IDinst/n8119 ), .DIN2(\IDinst/n8118 ), 
        .Q(\IDinst/n8120 ) );
  nnd2s1 \IDinst/U8164  ( .DIN1(\IDinst/n8117 ), .DIN2(n1159), 
        .Q(\IDinst/n8119 ) );
  nnd2s1 \IDinst/U8163  ( .DIN1(\IDinst/n8114 ), .DIN2(n1148), 
        .Q(\IDinst/n8118 ) );
  nnd2s1 \IDinst/U8162  ( .DIN1(\IDinst/n8116 ), .DIN2(\IDinst/n8115 ), 
        .Q(\IDinst/n8117 ) );
  nnd2s1 \IDinst/U8161  ( .DIN1(\IDinst/RegFile[15][23] ), .DIN2(n1096), 
        .Q(\IDinst/n8116 ) );
  nnd2s1 \IDinst/U8160  ( .DIN1(\IDinst/RegFile[14][23] ), .DIN2(n1064), 
        .Q(\IDinst/n8115 ) );
  nnd2s1 \IDinst/U8159  ( .DIN1(\IDinst/n8113 ), .DIN2(\IDinst/n8112 ), 
        .Q(\IDinst/n8114 ) );
  nnd2s1 \IDinst/U8158  ( .DIN1(\IDinst/RegFile[13][23] ), .DIN2(n1096), 
        .Q(\IDinst/n8113 ) );
  nnd2s1 \IDinst/U8157  ( .DIN1(\IDinst/RegFile[12][23] ), .DIN2(n1064), 
        .Q(\IDinst/n8112 ) );
  nnd2s1 \IDinst/U8156  ( .DIN1(\IDinst/n8110 ), .DIN2(\IDinst/n8109 ), 
        .Q(\IDinst/n8111 ) );
  nnd2s1 \IDinst/U8155  ( .DIN1(\IDinst/n8108 ), .DIN2(n1159), 
        .Q(\IDinst/n8110 ) );
  nnd2s1 \IDinst/U8154  ( .DIN1(\IDinst/n8105 ), .DIN2(n1148), 
        .Q(\IDinst/n8109 ) );
  nnd2s1 \IDinst/U8153  ( .DIN1(\IDinst/n8107 ), .DIN2(\IDinst/n8106 ), 
        .Q(\IDinst/n8108 ) );
  nnd2s1 \IDinst/U8152  ( .DIN1(\IDinst/RegFile[11][23] ), .DIN2(n1096), 
        .Q(\IDinst/n8107 ) );
  nnd2s1 \IDinst/U8151  ( .DIN1(\IDinst/RegFile[10][23] ), .DIN2(n1064), 
        .Q(\IDinst/n8106 ) );
  nnd2s1 \IDinst/U8150  ( .DIN1(\IDinst/n8104 ), .DIN2(\IDinst/n8103 ), 
        .Q(\IDinst/n8105 ) );
  nnd2s1 \IDinst/U8149  ( .DIN1(\IDinst/RegFile[9][23] ), .DIN2(n1073), 
        .Q(\IDinst/n8104 ) );
  nnd2s1 \IDinst/U8148  ( .DIN1(\IDinst/RegFile[8][23] ), .DIN2(n1064), 
        .Q(\IDinst/n8103 ) );
  nnd2s1 \IDinst/U8147  ( .DIN1(\IDinst/n8101 ), .DIN2(\IDinst/n8100 ), 
        .Q(\IDinst/n8102 ) );
  nnd2s1 \IDinst/U8146  ( .DIN1(\IDinst/n8099 ), .DIN2(n1190), 
        .Q(\IDinst/n8101 ) );
  nnd2s1 \IDinst/U8145  ( .DIN1(\IDinst/n8090 ), .DIN2(n1187), 
        .Q(\IDinst/n8100 ) );
  nnd2s1 \IDinst/U8144  ( .DIN1(\IDinst/n8098 ), .DIN2(\IDinst/n8097 ), 
        .Q(\IDinst/n8099 ) );
  nnd2s1 \IDinst/U8143  ( .DIN1(\IDinst/n8096 ), .DIN2(n1159), 
        .Q(\IDinst/n8098 ) );
  nnd2s1 \IDinst/U8142  ( .DIN1(\IDinst/n8093 ), .DIN2(n1149), 
        .Q(\IDinst/n8097 ) );
  nnd2s1 \IDinst/U8141  ( .DIN1(\IDinst/n8095 ), .DIN2(\IDinst/n8094 ), 
        .Q(\IDinst/n8096 ) );
  nnd2s1 \IDinst/U8140  ( .DIN1(\IDinst/RegFile[7][23] ), .DIN2(n1067), 
        .Q(\IDinst/n8095 ) );
  nnd2s1 \IDinst/U8139  ( .DIN1(\IDinst/RegFile[6][23] ), .DIN2(n1064), 
        .Q(\IDinst/n8094 ) );
  nnd2s1 \IDinst/U8138  ( .DIN1(\IDinst/n8092 ), .DIN2(\IDinst/n8091 ), 
        .Q(\IDinst/n8093 ) );
  nnd2s1 \IDinst/U8137  ( .DIN1(\IDinst/RegFile[5][23] ), .DIN2(n1065), 
        .Q(\IDinst/n8092 ) );
  nnd2s1 \IDinst/U8136  ( .DIN1(\IDinst/RegFile[4][23] ), .DIN2(n1064), 
        .Q(\IDinst/n8091 ) );
  nnd2s1 \IDinst/U8135  ( .DIN1(\IDinst/n8089 ), .DIN2(\IDinst/n8088 ), 
        .Q(\IDinst/n8090 ) );
  nnd2s1 \IDinst/U8134  ( .DIN1(\IDinst/n8087 ), .DIN2(n1159), 
        .Q(\IDinst/n8089 ) );
  nnd2s1 \IDinst/U8133  ( .DIN1(\IDinst/n8084 ), .DIN2(n1149), 
        .Q(\IDinst/n8088 ) );
  nnd2s1 \IDinst/U8132  ( .DIN1(\IDinst/n8086 ), .DIN2(\IDinst/n8085 ), 
        .Q(\IDinst/n8087 ) );
  nnd2s1 \IDinst/U8131  ( .DIN1(\IDinst/RegFile[3][23] ), .DIN2(n1066), 
        .Q(\IDinst/n8086 ) );
  nnd2s1 \IDinst/U8130  ( .DIN1(\IDinst/RegFile[2][23] ), .DIN2(n1063), 
        .Q(\IDinst/n8085 ) );
  nnd2s1 \IDinst/U8129  ( .DIN1(\IDinst/n8083 ), .DIN2(\IDinst/n8082 ), 
        .Q(\IDinst/n8084 ) );
  nnd2s1 \IDinst/U8128  ( .DIN1(\IDinst/RegFile[1][23] ), .DIN2(n1066), 
        .Q(\IDinst/n8083 ) );
  nnd2s1 \IDinst/U8127  ( .DIN1(\IDinst/RegFile[0][23] ), .DIN2(n1063), 
        .Q(\IDinst/n8082 ) );
  nnd2s1 \IDinst/U8126  ( .DIN1(\IDinst/n8081 ), .DIN2(n539), 
        .Q(\IDinst/n5992 ) );
  nnd2s1 \IDinst/U8125  ( .DIN1(\IDinst/n8036 ), .DIN2(n636), 
        .Q(\IDinst/n5993 ) );
  nnd2s1 \IDinst/U8124  ( .DIN1(\IDinst/n8080 ), .DIN2(\IDinst/n8079 ), 
        .Q(\IDinst/n8081 ) );
  nnd2s1 \IDinst/U8123  ( .DIN1(\IDinst/n8078 ), .DIN2(n641), 
        .Q(\IDinst/n8080 ) );
  nnd2s1 \IDinst/U8122  ( .DIN1(\IDinst/n8057 ), .DIN2(n671), 
        .Q(\IDinst/n8079 ) );
  nnd2s1 \IDinst/U8121  ( .DIN1(\IDinst/n8077 ), .DIN2(\IDinst/n8076 ), 
        .Q(\IDinst/n8078 ) );
  nnd2s1 \IDinst/U8120  ( .DIN1(\IDinst/n8075 ), .DIN2(n1190), 
        .Q(\IDinst/n8077 ) );
  nnd2s1 \IDinst/U8119  ( .DIN1(\IDinst/n8066 ), .DIN2(n1187), 
        .Q(\IDinst/n8076 ) );
  nnd2s1 \IDinst/U8118  ( .DIN1(\IDinst/n8074 ), .DIN2(\IDinst/n8073 ), 
        .Q(\IDinst/n8075 ) );
  nnd2s1 \IDinst/U8117  ( .DIN1(\IDinst/n8072 ), .DIN2(n1159), 
        .Q(\IDinst/n8074 ) );
  nnd2s1 \IDinst/U8116  ( .DIN1(\IDinst/n8069 ), .DIN2(n1149), 
        .Q(\IDinst/n8073 ) );
  nnd2s1 \IDinst/U8115  ( .DIN1(\IDinst/n8071 ), .DIN2(\IDinst/n8070 ), 
        .Q(\IDinst/n8072 ) );
  nnd2s1 \IDinst/U8114  ( .DIN1(\IDinst/RegFile[31][22] ), .DIN2(n1066), 
        .Q(\IDinst/n8071 ) );
  nnd2s1 \IDinst/U8113  ( .DIN1(\IDinst/RegFile[30][22] ), .DIN2(n1063), 
        .Q(\IDinst/n8070 ) );
  nnd2s1 \IDinst/U8112  ( .DIN1(\IDinst/n8068 ), .DIN2(\IDinst/n8067 ), 
        .Q(\IDinst/n8069 ) );
  nnd2s1 \IDinst/U8111  ( .DIN1(\IDinst/RegFile[29][22] ), .DIN2(n1066), 
        .Q(\IDinst/n8068 ) );
  nnd2s1 \IDinst/U8110  ( .DIN1(\IDinst/RegFile[28][22] ), .DIN2(n1063), 
        .Q(\IDinst/n8067 ) );
  nnd2s1 \IDinst/U8109  ( .DIN1(\IDinst/n8065 ), .DIN2(\IDinst/n8064 ), 
        .Q(\IDinst/n8066 ) );
  nnd2s1 \IDinst/U8108  ( .DIN1(\IDinst/n8063 ), .DIN2(n1159), 
        .Q(\IDinst/n8065 ) );
  nnd2s1 \IDinst/U8107  ( .DIN1(\IDinst/n8060 ), .DIN2(n1149), 
        .Q(\IDinst/n8064 ) );
  nnd2s1 \IDinst/U8106  ( .DIN1(\IDinst/n8062 ), .DIN2(\IDinst/n8061 ), 
        .Q(\IDinst/n8063 ) );
  nnd2s1 \IDinst/U8105  ( .DIN1(\IDinst/RegFile[27][22] ), .DIN2(n1066), 
        .Q(\IDinst/n8062 ) );
  nnd2s1 \IDinst/U8104  ( .DIN1(\IDinst/RegFile[26][22] ), .DIN2(n1063), 
        .Q(\IDinst/n8061 ) );
  nnd2s1 \IDinst/U8103  ( .DIN1(\IDinst/n8059 ), .DIN2(\IDinst/n8058 ), 
        .Q(\IDinst/n8060 ) );
  nnd2s1 \IDinst/U8102  ( .DIN1(\IDinst/RegFile[25][22] ), .DIN2(n1066), 
        .Q(\IDinst/n8059 ) );
  nnd2s1 \IDinst/U8101  ( .DIN1(\IDinst/RegFile[24][22] ), .DIN2(n1063), 
        .Q(\IDinst/n8058 ) );
  nnd2s1 \IDinst/U8100  ( .DIN1(\IDinst/n8056 ), .DIN2(\IDinst/n8055 ), 
        .Q(\IDinst/n8057 ) );
  nnd2s1 \IDinst/U8099  ( .DIN1(\IDinst/n8054 ), .DIN2(n1190), 
        .Q(\IDinst/n8056 ) );
  nnd2s1 \IDinst/U8098  ( .DIN1(\IDinst/n8045 ), .DIN2(n1187), 
        .Q(\IDinst/n8055 ) );
  nnd2s1 \IDinst/U8097  ( .DIN1(\IDinst/n8053 ), .DIN2(\IDinst/n8052 ), 
        .Q(\IDinst/n8054 ) );
  nnd2s1 \IDinst/U8096  ( .DIN1(\IDinst/n8051 ), .DIN2(n1159), 
        .Q(\IDinst/n8053 ) );
  nnd2s1 \IDinst/U8095  ( .DIN1(\IDinst/n8048 ), .DIN2(n1149), 
        .Q(\IDinst/n8052 ) );
  nnd2s1 \IDinst/U8094  ( .DIN1(\IDinst/n8050 ), .DIN2(\IDinst/n8049 ), 
        .Q(\IDinst/n8051 ) );
  nnd2s1 \IDinst/U8093  ( .DIN1(\IDinst/RegFile[23][22] ), .DIN2(n1066), 
        .Q(\IDinst/n8050 ) );
  nnd2s1 \IDinst/U8092  ( .DIN1(\IDinst/RegFile[22][22] ), .DIN2(n1063), 
        .Q(\IDinst/n8049 ) );
  nnd2s1 \IDinst/U8091  ( .DIN1(\IDinst/n8047 ), .DIN2(\IDinst/n8046 ), 
        .Q(\IDinst/n8048 ) );
  nnd2s1 \IDinst/U8090  ( .DIN1(\IDinst/RegFile[21][22] ), .DIN2(n1066), 
        .Q(\IDinst/n8047 ) );
  nnd2s1 \IDinst/U8089  ( .DIN1(\IDinst/RegFile[20][22] ), .DIN2(n1063), 
        .Q(\IDinst/n8046 ) );
  nnd2s1 \IDinst/U8088  ( .DIN1(\IDinst/n8044 ), .DIN2(\IDinst/n8043 ), 
        .Q(\IDinst/n8045 ) );
  nnd2s1 \IDinst/U8087  ( .DIN1(\IDinst/n8042 ), .DIN2(n1170), 
        .Q(\IDinst/n8044 ) );
  nnd2s1 \IDinst/U8086  ( .DIN1(\IDinst/n8039 ), .DIN2(n1149), 
        .Q(\IDinst/n8043 ) );
  nnd2s1 \IDinst/U8085  ( .DIN1(\IDinst/n8041 ), .DIN2(\IDinst/n8040 ), 
        .Q(\IDinst/n8042 ) );
  nnd2s1 \IDinst/U8084  ( .DIN1(\IDinst/RegFile[19][22] ), .DIN2(n1067), 
        .Q(\IDinst/n8041 ) );
  nnd2s1 \IDinst/U8083  ( .DIN1(\IDinst/RegFile[18][22] ), .DIN2(n1063), 
        .Q(\IDinst/n8040 ) );
  nnd2s1 \IDinst/U8082  ( .DIN1(\IDinst/n8038 ), .DIN2(\IDinst/n8037 ), 
        .Q(\IDinst/n8039 ) );
  nnd2s1 \IDinst/U8081  ( .DIN1(\IDinst/RegFile[17][22] ), .DIN2(n1066), 
        .Q(\IDinst/n8038 ) );
  nnd2s1 \IDinst/U8080  ( .DIN1(\IDinst/RegFile[16][22] ), .DIN2(n1063), 
        .Q(\IDinst/n8037 ) );
  nnd2s1 \IDinst/U8079  ( .DIN1(\IDinst/n8035 ), .DIN2(\IDinst/n8034 ), 
        .Q(\IDinst/n8036 ) );
  nnd2s1 \IDinst/U8078  ( .DIN1(\IDinst/n8033 ), .DIN2(n644), 
        .Q(\IDinst/n8035 ) );
  nnd2s1 \IDinst/U8077  ( .DIN1(\IDinst/n8012 ), .DIN2(n672), 
        .Q(\IDinst/n8034 ) );
  nnd2s1 \IDinst/U8076  ( .DIN1(\IDinst/n8032 ), .DIN2(\IDinst/n8031 ), 
        .Q(\IDinst/n8033 ) );
  nnd2s1 \IDinst/U8075  ( .DIN1(\IDinst/n8030 ), .DIN2(n1191), 
        .Q(\IDinst/n8032 ) );
  nnd2s1 \IDinst/U8074  ( .DIN1(\IDinst/n8021 ), .DIN2(n1187), 
        .Q(\IDinst/n8031 ) );
  nnd2s1 \IDinst/U8073  ( .DIN1(\IDinst/n8029 ), .DIN2(\IDinst/n8028 ), 
        .Q(\IDinst/n8030 ) );
  nnd2s1 \IDinst/U8072  ( .DIN1(\IDinst/n8027 ), .DIN2(n1176), 
        .Q(\IDinst/n8029 ) );
  nnd2s1 \IDinst/U8071  ( .DIN1(\IDinst/n8024 ), .DIN2(n1149), 
        .Q(\IDinst/n8028 ) );
  nnd2s1 \IDinst/U8070  ( .DIN1(\IDinst/n8026 ), .DIN2(\IDinst/n8025 ), 
        .Q(\IDinst/n8027 ) );
  nnd2s1 \IDinst/U8069  ( .DIN1(\IDinst/RegFile[15][22] ), .DIN2(n1067), 
        .Q(\IDinst/n8026 ) );
  nnd2s1 \IDinst/U8068  ( .DIN1(\IDinst/RegFile[14][22] ), .DIN2(n1063), 
        .Q(\IDinst/n8025 ) );
  nnd2s1 \IDinst/U8067  ( .DIN1(\IDinst/n8023 ), .DIN2(\IDinst/n8022 ), 
        .Q(\IDinst/n8024 ) );
  nnd2s1 \IDinst/U8066  ( .DIN1(\IDinst/RegFile[13][22] ), .DIN2(n1067), 
        .Q(\IDinst/n8023 ) );
  nnd2s1 \IDinst/U8065  ( .DIN1(\IDinst/RegFile[12][22] ), .DIN2(n1063), 
        .Q(\IDinst/n8022 ) );
  nnd2s1 \IDinst/U8064  ( .DIN1(\IDinst/n8020 ), .DIN2(\IDinst/n8019 ), 
        .Q(\IDinst/n8021 ) );
  nnd2s1 \IDinst/U8063  ( .DIN1(\IDinst/n8018 ), .DIN2(n1157), 
        .Q(\IDinst/n8020 ) );
  nnd2s1 \IDinst/U8062  ( .DIN1(\IDinst/n8015 ), .DIN2(n1149), 
        .Q(\IDinst/n8019 ) );
  nnd2s1 \IDinst/U8061  ( .DIN1(\IDinst/n8017 ), .DIN2(\IDinst/n8016 ), 
        .Q(\IDinst/n8018 ) );
  nnd2s1 \IDinst/U8060  ( .DIN1(\IDinst/RegFile[11][22] ), .DIN2(n1069), 
        .Q(\IDinst/n8017 ) );
  nnd2s1 \IDinst/U8059  ( .DIN1(\IDinst/RegFile[10][22] ), .DIN2(n1063), 
        .Q(\IDinst/n8016 ) );
  nnd2s1 \IDinst/U8058  ( .DIN1(\IDinst/n8014 ), .DIN2(\IDinst/n8013 ), 
        .Q(\IDinst/n8015 ) );
  nnd2s1 \IDinst/U8057  ( .DIN1(\IDinst/RegFile[9][22] ), .DIN2(n1067), 
        .Q(\IDinst/n8014 ) );
  nnd2s1 \IDinst/U8056  ( .DIN1(\IDinst/RegFile[8][22] ), .DIN2(n1062), 
        .Q(\IDinst/n8013 ) );
  nnd2s1 \IDinst/U8055  ( .DIN1(\IDinst/n8011 ), .DIN2(\IDinst/n8010 ), 
        .Q(\IDinst/n8012 ) );
  nnd2s1 \IDinst/U8054  ( .DIN1(\IDinst/n8009 ), .DIN2(n1191), 
        .Q(\IDinst/n8011 ) );
  nnd2s1 \IDinst/U8053  ( .DIN1(\IDinst/n8000 ), .DIN2(n1187), 
        .Q(\IDinst/n8010 ) );
  nnd2s1 \IDinst/U8052  ( .DIN1(\IDinst/n8008 ), .DIN2(\IDinst/n8007 ), 
        .Q(\IDinst/n8009 ) );
  nnd2s1 \IDinst/U8051  ( .DIN1(\IDinst/n8006 ), .DIN2(n1158), 
        .Q(\IDinst/n8008 ) );
  nnd2s1 \IDinst/U8050  ( .DIN1(\IDinst/n8003 ), .DIN2(n1149), 
        .Q(\IDinst/n8007 ) );
  nnd2s1 \IDinst/U8049  ( .DIN1(\IDinst/n8005 ), .DIN2(\IDinst/n8004 ), 
        .Q(\IDinst/n8006 ) );
  nnd2s1 \IDinst/U8048  ( .DIN1(\IDinst/RegFile[7][22] ), .DIN2(n1068), 
        .Q(\IDinst/n8005 ) );
  nnd2s1 \IDinst/U8047  ( .DIN1(\IDinst/RegFile[6][22] ), .DIN2(n1062), 
        .Q(\IDinst/n8004 ) );
  nnd2s1 \IDinst/U8046  ( .DIN1(\IDinst/n8002 ), .DIN2(\IDinst/n8001 ), 
        .Q(\IDinst/n8003 ) );
  nnd2s1 \IDinst/U8045  ( .DIN1(\IDinst/RegFile[5][22] ), .DIN2(n1067), 
        .Q(\IDinst/n8002 ) );
  nnd2s1 \IDinst/U8044  ( .DIN1(\IDinst/RegFile[4][22] ), .DIN2(n1062), 
        .Q(\IDinst/n8001 ) );
  nnd2s1 \IDinst/U8043  ( .DIN1(\IDinst/n7999 ), .DIN2(\IDinst/n7998 ), 
        .Q(\IDinst/n8000 ) );
  nnd2s1 \IDinst/U8042  ( .DIN1(\IDinst/n7997 ), .DIN2(n1153), 
        .Q(\IDinst/n7999 ) );
  nnd2s1 \IDinst/U8041  ( .DIN1(\IDinst/n7994 ), .DIN2(n1149), 
        .Q(\IDinst/n7998 ) );
  nnd2s1 \IDinst/U8040  ( .DIN1(\IDinst/n7996 ), .DIN2(\IDinst/n7995 ), 
        .Q(\IDinst/n7997 ) );
  nnd2s1 \IDinst/U8039  ( .DIN1(\IDinst/RegFile[3][22] ), .DIN2(n1067), 
        .Q(\IDinst/n7996 ) );
  nnd2s1 \IDinst/U8038  ( .DIN1(\IDinst/RegFile[2][22] ), .DIN2(n1062), 
        .Q(\IDinst/n7995 ) );
  nnd2s1 \IDinst/U8037  ( .DIN1(\IDinst/n7993 ), .DIN2(\IDinst/n7992 ), 
        .Q(\IDinst/n7994 ) );
  nnd2s1 \IDinst/U8036  ( .DIN1(\IDinst/RegFile[1][22] ), .DIN2(n1067), 
        .Q(\IDinst/n7993 ) );
  nnd2s1 \IDinst/U8035  ( .DIN1(\IDinst/RegFile[0][22] ), .DIN2(n1062), 
        .Q(\IDinst/n7992 ) );
  nnd2s1 \IDinst/U8034  ( .DIN1(\IDinst/n7991 ), .DIN2(n539), 
        .Q(\IDinst/n5990 ) );
  nnd2s1 \IDinst/U8033  ( .DIN1(\IDinst/n7946 ), .DIN2(n635), 
        .Q(\IDinst/n5991 ) );
  nnd2s1 \IDinst/U8032  ( .DIN1(\IDinst/n7990 ), .DIN2(\IDinst/n7989 ), 
        .Q(\IDinst/n7991 ) );
  nnd2s1 \IDinst/U8031  ( .DIN1(\IDinst/n7988 ), .DIN2(n643), 
        .Q(\IDinst/n7990 ) );
  nnd2s1 \IDinst/U8030  ( .DIN1(\IDinst/n7967 ), .DIN2(n670), 
        .Q(\IDinst/n7989 ) );
  nnd2s1 \IDinst/U8029  ( .DIN1(\IDinst/n7987 ), .DIN2(\IDinst/n7986 ), 
        .Q(\IDinst/n7988 ) );
  nnd2s1 \IDinst/U8028  ( .DIN1(\IDinst/n7985 ), .DIN2(n1191), 
        .Q(\IDinst/n7987 ) );
  nnd2s1 \IDinst/U8027  ( .DIN1(\IDinst/n7976 ), .DIN2(n1187), 
        .Q(\IDinst/n7986 ) );
  nnd2s1 \IDinst/U8026  ( .DIN1(\IDinst/n7984 ), .DIN2(\IDinst/n7983 ), 
        .Q(\IDinst/n7985 ) );
  nnd2s1 \IDinst/U8025  ( .DIN1(\IDinst/n7982 ), .DIN2(n1178), 
        .Q(\IDinst/n7984 ) );
  nnd2s1 \IDinst/U8024  ( .DIN1(\IDinst/n7979 ), .DIN2(n1149), 
        .Q(\IDinst/n7983 ) );
  nnd2s1 \IDinst/U8023  ( .DIN1(\IDinst/n7981 ), .DIN2(\IDinst/n7980 ), 
        .Q(\IDinst/n7982 ) );
  nnd2s1 \IDinst/U8022  ( .DIN1(\IDinst/RegFile[31][21] ), .DIN2(n1067), 
        .Q(\IDinst/n7981 ) );
  nnd2s1 \IDinst/U8021  ( .DIN1(\IDinst/RegFile[30][21] ), .DIN2(n1062), 
        .Q(\IDinst/n7980 ) );
  nnd2s1 \IDinst/U8020  ( .DIN1(\IDinst/n7978 ), .DIN2(\IDinst/n7977 ), 
        .Q(\IDinst/n7979 ) );
  nnd2s1 \IDinst/U8019  ( .DIN1(\IDinst/RegFile[29][21] ), .DIN2(n1068), 
        .Q(\IDinst/n7978 ) );
  nnd2s1 \IDinst/U8018  ( .DIN1(\IDinst/RegFile[28][21] ), .DIN2(n1062), 
        .Q(\IDinst/n7977 ) );
  nnd2s1 \IDinst/U8017  ( .DIN1(\IDinst/n7975 ), .DIN2(\IDinst/n7974 ), 
        .Q(\IDinst/n7976 ) );
  nnd2s1 \IDinst/U8016  ( .DIN1(\IDinst/n7973 ), .DIN2(n1179), 
        .Q(\IDinst/n7975 ) );
  nnd2s1 \IDinst/U8015  ( .DIN1(\IDinst/n7970 ), .DIN2(n1149), 
        .Q(\IDinst/n7974 ) );
  nnd2s1 \IDinst/U8014  ( .DIN1(\IDinst/n7972 ), .DIN2(\IDinst/n7971 ), 
        .Q(\IDinst/n7973 ) );
  nnd2s1 \IDinst/U8013  ( .DIN1(\IDinst/RegFile[27][21] ), .DIN2(n1068), 
        .Q(\IDinst/n7972 ) );
  nnd2s1 \IDinst/U8012  ( .DIN1(\IDinst/RegFile[26][21] ), .DIN2(n1062), 
        .Q(\IDinst/n7971 ) );
  nnd2s1 \IDinst/U8011  ( .DIN1(\IDinst/n7969 ), .DIN2(\IDinst/n7968 ), 
        .Q(\IDinst/n7970 ) );
  nnd2s1 \IDinst/U8010  ( .DIN1(\IDinst/RegFile[25][21] ), .DIN2(n1068), 
        .Q(\IDinst/n7969 ) );
  nnd2s1 \IDinst/U8009  ( .DIN1(\IDinst/RegFile[24][21] ), .DIN2(n1062), 
        .Q(\IDinst/n7968 ) );
  nnd2s1 \IDinst/U8008  ( .DIN1(\IDinst/n7966 ), .DIN2(\IDinst/n7965 ), 
        .Q(\IDinst/n7967 ) );
  nnd2s1 \IDinst/U8007  ( .DIN1(\IDinst/n7964 ), .DIN2(n1191), 
        .Q(\IDinst/n7966 ) );
  nnd2s1 \IDinst/U8006  ( .DIN1(\IDinst/n7955 ), .DIN2(n1187), 
        .Q(\IDinst/n7965 ) );
  nnd2s1 \IDinst/U8005  ( .DIN1(\IDinst/n7963 ), .DIN2(\IDinst/n7962 ), 
        .Q(\IDinst/n7964 ) );
  nnd2s1 \IDinst/U8004  ( .DIN1(\IDinst/n7961 ), .DIN2(\IDinst/N40 ), 
        .Q(\IDinst/n7963 ) );
  nnd2s1 \IDinst/U8003  ( .DIN1(\IDinst/n7958 ), .DIN2(n1149), 
        .Q(\IDinst/n7962 ) );
  nnd2s1 \IDinst/U8002  ( .DIN1(\IDinst/n7960 ), .DIN2(\IDinst/n7959 ), 
        .Q(\IDinst/n7961 ) );
  nnd2s1 \IDinst/U8001  ( .DIN1(\IDinst/RegFile[23][21] ), .DIN2(n1068), 
        .Q(\IDinst/n7960 ) );
  nnd2s1 \IDinst/U8000  ( .DIN1(\IDinst/RegFile[22][21] ), .DIN2(n1062), 
        .Q(\IDinst/n7959 ) );
  nnd2s1 \IDinst/U7999  ( .DIN1(\IDinst/n7957 ), .DIN2(\IDinst/n7956 ), 
        .Q(\IDinst/n7958 ) );
  nnd2s1 \IDinst/U7998  ( .DIN1(\IDinst/RegFile[21][21] ), .DIN2(n1068), 
        .Q(\IDinst/n7957 ) );
  nnd2s1 \IDinst/U7997  ( .DIN1(\IDinst/RegFile[20][21] ), .DIN2(n1062), 
        .Q(\IDinst/n7956 ) );
  nnd2s1 \IDinst/U7996  ( .DIN1(\IDinst/n7954 ), .DIN2(\IDinst/n7953 ), 
        .Q(\IDinst/n7955 ) );
  nnd2s1 \IDinst/U7995  ( .DIN1(\IDinst/n7952 ), .DIN2(n1154), 
        .Q(\IDinst/n7954 ) );
  nnd2s1 \IDinst/U7994  ( .DIN1(\IDinst/n7949 ), .DIN2(n1150), 
        .Q(\IDinst/n7953 ) );
  nnd2s1 \IDinst/U7993  ( .DIN1(\IDinst/n7951 ), .DIN2(\IDinst/n7950 ), 
        .Q(\IDinst/n7952 ) );
  nnd2s1 \IDinst/U7992  ( .DIN1(\IDinst/RegFile[19][21] ), .DIN2(n1068), 
        .Q(\IDinst/n7951 ) );
  nnd2s1 \IDinst/U7991  ( .DIN1(\IDinst/RegFile[18][21] ), .DIN2(n1062), 
        .Q(\IDinst/n7950 ) );
  nnd2s1 \IDinst/U7990  ( .DIN1(\IDinst/n7948 ), .DIN2(\IDinst/n7947 ), 
        .Q(\IDinst/n7949 ) );
  nnd2s1 \IDinst/U7989  ( .DIN1(\IDinst/RegFile[17][21] ), .DIN2(n1068), 
        .Q(\IDinst/n7948 ) );
  nnd2s1 \IDinst/U7988  ( .DIN1(\IDinst/RegFile[16][21] ), .DIN2(n1062), 
        .Q(\IDinst/n7947 ) );
  nnd2s1 \IDinst/U7987  ( .DIN1(\IDinst/n7945 ), .DIN2(\IDinst/n7944 ), 
        .Q(\IDinst/n7946 ) );
  nnd2s1 \IDinst/U7986  ( .DIN1(\IDinst/n7943 ), .DIN2(n642), 
        .Q(\IDinst/n7945 ) );
  nnd2s1 \IDinst/U7985  ( .DIN1(\IDinst/n7922 ), .DIN2(n673), 
        .Q(\IDinst/n7944 ) );
  nnd2s1 \IDinst/U7984  ( .DIN1(\IDinst/n7942 ), .DIN2(\IDinst/n7941 ), 
        .Q(\IDinst/n7943 ) );
  nnd2s1 \IDinst/U7983  ( .DIN1(\IDinst/n7940 ), .DIN2(n1191), 
        .Q(\IDinst/n7942 ) );
  nnd2s1 \IDinst/U7982  ( .DIN1(\IDinst/n7931 ), .DIN2(n1187), 
        .Q(\IDinst/n7941 ) );
  nnd2s1 \IDinst/U7981  ( .DIN1(\IDinst/n7939 ), .DIN2(\IDinst/n7938 ), 
        .Q(\IDinst/n7940 ) );
  nnd2s1 \IDinst/U7980  ( .DIN1(\IDinst/n7937 ), .DIN2(n1158), 
        .Q(\IDinst/n7939 ) );
  nnd2s1 \IDinst/U7979  ( .DIN1(\IDinst/n7934 ), .DIN2(n1150), 
        .Q(\IDinst/n7938 ) );
  nnd2s1 \IDinst/U7978  ( .DIN1(\IDinst/n7936 ), .DIN2(\IDinst/n7935 ), 
        .Q(\IDinst/n7937 ) );
  nnd2s1 \IDinst/U7977  ( .DIN1(\IDinst/RegFile[15][21] ), .DIN2(n1070), 
        .Q(\IDinst/n7936 ) );
  nnd2s1 \IDinst/U7976  ( .DIN1(\IDinst/RegFile[14][21] ), .DIN2(n1061), 
        .Q(\IDinst/n7935 ) );
  nnd2s1 \IDinst/U7975  ( .DIN1(\IDinst/n7933 ), .DIN2(\IDinst/n7932 ), 
        .Q(\IDinst/n7934 ) );
  nnd2s1 \IDinst/U7974  ( .DIN1(\IDinst/RegFile[13][21] ), .DIN2(n1068), 
        .Q(\IDinst/n7933 ) );
  nnd2s1 \IDinst/U7973  ( .DIN1(\IDinst/RegFile[12][21] ), .DIN2(n1061), 
        .Q(\IDinst/n7932 ) );
  nnd2s1 \IDinst/U7972  ( .DIN1(\IDinst/n7930 ), .DIN2(\IDinst/n7929 ), 
        .Q(\IDinst/n7931 ) );
  nnd2s1 \IDinst/U7971  ( .DIN1(\IDinst/n7928 ), .DIN2(n1158), 
        .Q(\IDinst/n7930 ) );
  nnd2s1 \IDinst/U7970  ( .DIN1(\IDinst/n7925 ), .DIN2(n1150), 
        .Q(\IDinst/n7929 ) );
  nnd2s1 \IDinst/U7969  ( .DIN1(\IDinst/n7927 ), .DIN2(\IDinst/n7926 ), 
        .Q(\IDinst/n7928 ) );
  nnd2s1 \IDinst/U7968  ( .DIN1(\IDinst/RegFile[11][21] ), .DIN2(n1069), 
        .Q(\IDinst/n7927 ) );
  nnd2s1 \IDinst/U7967  ( .DIN1(\IDinst/RegFile[10][21] ), .DIN2(n1061), 
        .Q(\IDinst/n7926 ) );
  nnd2s1 \IDinst/U7966  ( .DIN1(\IDinst/n7924 ), .DIN2(\IDinst/n7923 ), 
        .Q(\IDinst/n7925 ) );
  nnd2s1 \IDinst/U7965  ( .DIN1(\IDinst/RegFile[9][21] ), .DIN2(n1069), 
        .Q(\IDinst/n7924 ) );
  nnd2s1 \IDinst/U7964  ( .DIN1(\IDinst/RegFile[8][21] ), .DIN2(n1061), 
        .Q(\IDinst/n7923 ) );
  nnd2s1 \IDinst/U7963  ( .DIN1(\IDinst/n7921 ), .DIN2(\IDinst/n7920 ), 
        .Q(\IDinst/n7922 ) );
  nnd2s1 \IDinst/U7962  ( .DIN1(\IDinst/n7919 ), .DIN2(n1191), 
        .Q(\IDinst/n7921 ) );
  nnd2s1 \IDinst/U7961  ( .DIN1(\IDinst/n7910 ), .DIN2(n1187), 
        .Q(\IDinst/n7920 ) );
  nnd2s1 \IDinst/U7960  ( .DIN1(\IDinst/n7918 ), .DIN2(\IDinst/n7917 ), 
        .Q(\IDinst/n7919 ) );
  nnd2s1 \IDinst/U7959  ( .DIN1(\IDinst/n7916 ), .DIN2(n1158), 
        .Q(\IDinst/n7918 ) );
  nnd2s1 \IDinst/U7958  ( .DIN1(\IDinst/n7913 ), .DIN2(n1150), 
        .Q(\IDinst/n7917 ) );
  nnd2s1 \IDinst/U7957  ( .DIN1(\IDinst/n7915 ), .DIN2(\IDinst/n7914 ), 
        .Q(\IDinst/n7916 ) );
  nnd2s1 \IDinst/U7956  ( .DIN1(\IDinst/RegFile[7][21] ), .DIN2(n1069), 
        .Q(\IDinst/n7915 ) );
  nnd2s1 \IDinst/U7955  ( .DIN1(\IDinst/RegFile[6][21] ), .DIN2(n1061), 
        .Q(\IDinst/n7914 ) );
  nnd2s1 \IDinst/U7954  ( .DIN1(\IDinst/n7912 ), .DIN2(\IDinst/n7911 ), 
        .Q(\IDinst/n7913 ) );
  nnd2s1 \IDinst/U7953  ( .DIN1(\IDinst/RegFile[5][21] ), .DIN2(n1069), 
        .Q(\IDinst/n7912 ) );
  nnd2s1 \IDinst/U7952  ( .DIN1(\IDinst/RegFile[4][21] ), .DIN2(n1061), 
        .Q(\IDinst/n7911 ) );
  nnd2s1 \IDinst/U7951  ( .DIN1(\IDinst/n7909 ), .DIN2(\IDinst/n7908 ), 
        .Q(\IDinst/n7910 ) );
  nnd2s1 \IDinst/U7950  ( .DIN1(\IDinst/n7907 ), .DIN2(n1158), 
        .Q(\IDinst/n7909 ) );
  nnd2s1 \IDinst/U7949  ( .DIN1(\IDinst/n7904 ), .DIN2(n1150), 
        .Q(\IDinst/n7908 ) );
  nnd2s1 \IDinst/U7948  ( .DIN1(\IDinst/n7906 ), .DIN2(\IDinst/n7905 ), 
        .Q(\IDinst/n7907 ) );
  nnd2s1 \IDinst/U7947  ( .DIN1(\IDinst/RegFile[3][21] ), .DIN2(n1070), 
        .Q(\IDinst/n7906 ) );
  nnd2s1 \IDinst/U7946  ( .DIN1(\IDinst/RegFile[2][21] ), .DIN2(n1061), 
        .Q(\IDinst/n7905 ) );
  nnd2s1 \IDinst/U7945  ( .DIN1(\IDinst/n7903 ), .DIN2(\IDinst/n7902 ), 
        .Q(\IDinst/n7904 ) );
  nnd2s1 \IDinst/U7944  ( .DIN1(\IDinst/RegFile[1][21] ), .DIN2(n1069), 
        .Q(\IDinst/n7903 ) );
  nnd2s1 \IDinst/U7943  ( .DIN1(\IDinst/RegFile[0][21] ), .DIN2(n1061), 
        .Q(\IDinst/n7902 ) );
  nnd2s1 \IDinst/U7942  ( .DIN1(\IDinst/n7901 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n5988 ) );
  nnd2s1 \IDinst/U7941  ( .DIN1(\IDinst/n7856 ), .DIN2(n636), 
        .Q(\IDinst/n5989 ) );
  nnd2s1 \IDinst/U7940  ( .DIN1(\IDinst/n7900 ), .DIN2(\IDinst/n7899 ), 
        .Q(\IDinst/n7901 ) );
  nnd2s1 \IDinst/U7939  ( .DIN1(\IDinst/n7898 ), .DIN2(n641), 
        .Q(\IDinst/n7900 ) );
  nnd2s1 \IDinst/U7938  ( .DIN1(\IDinst/n7877 ), .DIN2(n671), 
        .Q(\IDinst/n7899 ) );
  nnd2s1 \IDinst/U7937  ( .DIN1(\IDinst/n7897 ), .DIN2(\IDinst/n7896 ), 
        .Q(\IDinst/n7898 ) );
  nnd2s1 \IDinst/U7936  ( .DIN1(\IDinst/n7895 ), .DIN2(n1191), 
        .Q(\IDinst/n7897 ) );
  nnd2s1 \IDinst/U7935  ( .DIN1(\IDinst/n7886 ), .DIN2(n1187), 
        .Q(\IDinst/n7896 ) );
  nnd2s1 \IDinst/U7934  ( .DIN1(\IDinst/n7894 ), .DIN2(\IDinst/n7893 ), 
        .Q(\IDinst/n7895 ) );
  nnd2s1 \IDinst/U7933  ( .DIN1(\IDinst/n7892 ), .DIN2(n1158), 
        .Q(\IDinst/n7894 ) );
  nnd2s1 \IDinst/U7932  ( .DIN1(\IDinst/n7889 ), .DIN2(n1150), 
        .Q(\IDinst/n7893 ) );
  nnd2s1 \IDinst/U7931  ( .DIN1(\IDinst/n7891 ), .DIN2(\IDinst/n7890 ), 
        .Q(\IDinst/n7892 ) );
  nnd2s1 \IDinst/U7930  ( .DIN1(\IDinst/RegFile[31][20] ), .DIN2(n1069), 
        .Q(\IDinst/n7891 ) );
  nnd2s1 \IDinst/U7929  ( .DIN1(\IDinst/RegFile[30][20] ), .DIN2(n1061), 
        .Q(\IDinst/n7890 ) );
  nnd2s1 \IDinst/U7928  ( .DIN1(\IDinst/n7888 ), .DIN2(\IDinst/n7887 ), 
        .Q(\IDinst/n7889 ) );
  nnd2s1 \IDinst/U7927  ( .DIN1(\IDinst/RegFile[29][20] ), .DIN2(n1069), 
        .Q(\IDinst/n7888 ) );
  nnd2s1 \IDinst/U7926  ( .DIN1(\IDinst/RegFile[28][20] ), .DIN2(n1061), 
        .Q(\IDinst/n7887 ) );
  nnd2s1 \IDinst/U7925  ( .DIN1(\IDinst/n7885 ), .DIN2(\IDinst/n7884 ), 
        .Q(\IDinst/n7886 ) );
  nnd2s1 \IDinst/U7924  ( .DIN1(\IDinst/n7883 ), .DIN2(n1158), 
        .Q(\IDinst/n7885 ) );
  nnd2s1 \IDinst/U7923  ( .DIN1(\IDinst/n7880 ), .DIN2(n1150), 
        .Q(\IDinst/n7884 ) );
  nnd2s1 \IDinst/U7922  ( .DIN1(\IDinst/n7882 ), .DIN2(\IDinst/n7881 ), 
        .Q(\IDinst/n7883 ) );
  nnd2s1 \IDinst/U7921  ( .DIN1(\IDinst/RegFile[27][20] ), .DIN2(n1069), 
        .Q(\IDinst/n7882 ) );
  nnd2s1 \IDinst/U7920  ( .DIN1(\IDinst/RegFile[26][20] ), .DIN2(n1061), 
        .Q(\IDinst/n7881 ) );
  nnd2s1 \IDinst/U7919  ( .DIN1(\IDinst/n7879 ), .DIN2(\IDinst/n7878 ), 
        .Q(\IDinst/n7880 ) );
  nnd2s1 \IDinst/U7918  ( .DIN1(\IDinst/RegFile[25][20] ), .DIN2(n1070), 
        .Q(\IDinst/n7879 ) );
  nnd2s1 \IDinst/U7917  ( .DIN1(\IDinst/RegFile[24][20] ), .DIN2(n1061), 
        .Q(\IDinst/n7878 ) );
  nnd2s1 \IDinst/U7916  ( .DIN1(\IDinst/n7876 ), .DIN2(\IDinst/n7875 ), 
        .Q(\IDinst/n7877 ) );
  nnd2s1 \IDinst/U7915  ( .DIN1(\IDinst/n7874 ), .DIN2(n1191), 
        .Q(\IDinst/n7876 ) );
  nnd2s1 \IDinst/U7914  ( .DIN1(\IDinst/n7865 ), .DIN2(n1186), 
        .Q(\IDinst/n7875 ) );
  nnd2s1 \IDinst/U7913  ( .DIN1(\IDinst/n7873 ), .DIN2(\IDinst/n7872 ), 
        .Q(\IDinst/n7874 ) );
  nnd2s1 \IDinst/U7912  ( .DIN1(\IDinst/n7871 ), .DIN2(n1158), 
        .Q(\IDinst/n7873 ) );
  nnd2s1 \IDinst/U7911  ( .DIN1(\IDinst/n7868 ), .DIN2(n1150), 
        .Q(\IDinst/n7872 ) );
  nnd2s1 \IDinst/U7910  ( .DIN1(\IDinst/n7870 ), .DIN2(\IDinst/n7869 ), 
        .Q(\IDinst/n7871 ) );
  nnd2s1 \IDinst/U7909  ( .DIN1(\IDinst/RegFile[23][20] ), .DIN2(n1070), 
        .Q(\IDinst/n7870 ) );
  nnd2s1 \IDinst/U7908  ( .DIN1(\IDinst/RegFile[22][20] ), .DIN2(n1061), 
        .Q(\IDinst/n7869 ) );
  nnd2s1 \IDinst/U7907  ( .DIN1(\IDinst/n7867 ), .DIN2(\IDinst/n7866 ), 
        .Q(\IDinst/n7868 ) );
  nnd2s1 \IDinst/U7906  ( .DIN1(\IDinst/RegFile[21][20] ), .DIN2(n1070), 
        .Q(\IDinst/n7867 ) );
  nnd2s1 \IDinst/U7905  ( .DIN1(\IDinst/RegFile[20][20] ), .DIN2(n1060), 
        .Q(\IDinst/n7866 ) );
  nnd2s1 \IDinst/U7904  ( .DIN1(\IDinst/n7864 ), .DIN2(\IDinst/n7863 ), 
        .Q(\IDinst/n7865 ) );
  nnd2s1 \IDinst/U7903  ( .DIN1(\IDinst/n7862 ), .DIN2(n1158), 
        .Q(\IDinst/n7864 ) );
  nnd2s1 \IDinst/U7902  ( .DIN1(\IDinst/n7859 ), .DIN2(n1150), 
        .Q(\IDinst/n7863 ) );
  nnd2s1 \IDinst/U7901  ( .DIN1(\IDinst/n7861 ), .DIN2(\IDinst/n7860 ), 
        .Q(\IDinst/n7862 ) );
  nnd2s1 \IDinst/U7900  ( .DIN1(\IDinst/RegFile[19][20] ), .DIN2(n1070), 
        .Q(\IDinst/n7861 ) );
  nnd2s1 \IDinst/U7899  ( .DIN1(\IDinst/RegFile[18][20] ), .DIN2(n1060), 
        .Q(\IDinst/n7860 ) );
  nnd2s1 \IDinst/U7898  ( .DIN1(\IDinst/n7858 ), .DIN2(\IDinst/n7857 ), 
        .Q(\IDinst/n7859 ) );
  nnd2s1 \IDinst/U7897  ( .DIN1(\IDinst/RegFile[17][20] ), .DIN2(n1070), 
        .Q(\IDinst/n7858 ) );
  nnd2s1 \IDinst/U7896  ( .DIN1(\IDinst/RegFile[16][20] ), .DIN2(n1060), 
        .Q(\IDinst/n7857 ) );
  nnd2s1 \IDinst/U7895  ( .DIN1(\IDinst/n7855 ), .DIN2(\IDinst/n7854 ), 
        .Q(\IDinst/n7856 ) );
  nnd2s1 \IDinst/U7894  ( .DIN1(\IDinst/n7853 ), .DIN2(n644), 
        .Q(\IDinst/n7855 ) );
  nnd2s1 \IDinst/U7893  ( .DIN1(\IDinst/n7832 ), .DIN2(n672), 
        .Q(\IDinst/n7854 ) );
  nnd2s1 \IDinst/U7892  ( .DIN1(\IDinst/n7852 ), .DIN2(\IDinst/n7851 ), 
        .Q(\IDinst/n7853 ) );
  nnd2s1 \IDinst/U7891  ( .DIN1(\IDinst/n7850 ), .DIN2(n1191), 
        .Q(\IDinst/n7852 ) );
  nnd2s1 \IDinst/U7890  ( .DIN1(\IDinst/n7841 ), .DIN2(n1186), 
        .Q(\IDinst/n7851 ) );
  nnd2s1 \IDinst/U7889  ( .DIN1(\IDinst/n7849 ), .DIN2(\IDinst/n7848 ), 
        .Q(\IDinst/n7850 ) );
  nnd2s1 \IDinst/U7888  ( .DIN1(\IDinst/n7847 ), .DIN2(n1158), 
        .Q(\IDinst/n7849 ) );
  nnd2s1 \IDinst/U7887  ( .DIN1(\IDinst/n7844 ), .DIN2(n1150), 
        .Q(\IDinst/n7848 ) );
  nnd2s1 \IDinst/U7886  ( .DIN1(\IDinst/n7846 ), .DIN2(\IDinst/n7845 ), 
        .Q(\IDinst/n7847 ) );
  nnd2s1 \IDinst/U7885  ( .DIN1(\IDinst/RegFile[15][20] ), .DIN2(n1070), 
        .Q(\IDinst/n7846 ) );
  nnd2s1 \IDinst/U7884  ( .DIN1(\IDinst/RegFile[14][20] ), .DIN2(n1060), 
        .Q(\IDinst/n7845 ) );
  nnd2s1 \IDinst/U7883  ( .DIN1(\IDinst/n7843 ), .DIN2(\IDinst/n7842 ), 
        .Q(\IDinst/n7844 ) );
  nnd2s1 \IDinst/U7882  ( .DIN1(\IDinst/RegFile[13][20] ), .DIN2(n1070), 
        .Q(\IDinst/n7843 ) );
  nnd2s1 \IDinst/U7881  ( .DIN1(\IDinst/RegFile[12][20] ), .DIN2(n1060), 
        .Q(\IDinst/n7842 ) );
  nnd2s1 \IDinst/U7880  ( .DIN1(\IDinst/n7840 ), .DIN2(\IDinst/n7839 ), 
        .Q(\IDinst/n7841 ) );
  nnd2s1 \IDinst/U7879  ( .DIN1(\IDinst/n7838 ), .DIN2(n1157), 
        .Q(\IDinst/n7840 ) );
  nnd2s1 \IDinst/U7878  ( .DIN1(\IDinst/n7835 ), .DIN2(n1150), 
        .Q(\IDinst/n7839 ) );
  nnd2s1 \IDinst/U7877  ( .DIN1(\IDinst/n7837 ), .DIN2(\IDinst/n7836 ), 
        .Q(\IDinst/n7838 ) );
  nnd2s1 \IDinst/U7876  ( .DIN1(\IDinst/RegFile[11][20] ), .DIN2(n1071), 
        .Q(\IDinst/n7837 ) );
  nnd2s1 \IDinst/U7875  ( .DIN1(\IDinst/RegFile[10][20] ), .DIN2(n1060), 
        .Q(\IDinst/n7836 ) );
  nnd2s1 \IDinst/U7874  ( .DIN1(\IDinst/n7834 ), .DIN2(\IDinst/n7833 ), 
        .Q(\IDinst/n7835 ) );
  nnd2s1 \IDinst/U7873  ( .DIN1(\IDinst/RegFile[9][20] ), .DIN2(n1071), 
        .Q(\IDinst/n7834 ) );
  nnd2s1 \IDinst/U7872  ( .DIN1(\IDinst/RegFile[8][20] ), .DIN2(n1060), 
        .Q(\IDinst/n7833 ) );
  nnd2s1 \IDinst/U7871  ( .DIN1(\IDinst/n7831 ), .DIN2(\IDinst/n7830 ), 
        .Q(\IDinst/n7832 ) );
  nnd2s1 \IDinst/U7870  ( .DIN1(\IDinst/n7829 ), .DIN2(n1197), 
        .Q(\IDinst/n7831 ) );
  nnd2s1 \IDinst/U7869  ( .DIN1(\IDinst/n7820 ), .DIN2(n1186), 
        .Q(\IDinst/n7830 ) );
  nnd2s1 \IDinst/U7868  ( .DIN1(\IDinst/n7828 ), .DIN2(\IDinst/n7827 ), 
        .Q(\IDinst/n7829 ) );
  nnd2s1 \IDinst/U7867  ( .DIN1(\IDinst/n7826 ), .DIN2(n1157), 
        .Q(\IDinst/n7828 ) );
  nnd2s1 \IDinst/U7866  ( .DIN1(\IDinst/n7823 ), .DIN2(n1150), 
        .Q(\IDinst/n7827 ) );
  nnd2s1 \IDinst/U7865  ( .DIN1(\IDinst/n7825 ), .DIN2(\IDinst/n7824 ), 
        .Q(\IDinst/n7826 ) );
  nnd2s1 \IDinst/U7864  ( .DIN1(\IDinst/RegFile[7][20] ), .DIN2(n1071), 
        .Q(\IDinst/n7825 ) );
  nnd2s1 \IDinst/U7863  ( .DIN1(\IDinst/RegFile[6][20] ), .DIN2(n1060), 
        .Q(\IDinst/n7824 ) );
  nnd2s1 \IDinst/U7862  ( .DIN1(\IDinst/n7822 ), .DIN2(\IDinst/n7821 ), 
        .Q(\IDinst/n7823 ) );
  nnd2s1 \IDinst/U7861  ( .DIN1(\IDinst/RegFile[5][20] ), .DIN2(n1071), 
        .Q(\IDinst/n7822 ) );
  nnd2s1 \IDinst/U7860  ( .DIN1(\IDinst/RegFile[4][20] ), .DIN2(n1060), 
        .Q(\IDinst/n7821 ) );
  nnd2s1 \IDinst/U7859  ( .DIN1(\IDinst/n7819 ), .DIN2(\IDinst/n7818 ), 
        .Q(\IDinst/n7820 ) );
  nnd2s1 \IDinst/U7858  ( .DIN1(\IDinst/n7817 ), .DIN2(n1157), 
        .Q(\IDinst/n7819 ) );
  nnd2s1 \IDinst/U7857  ( .DIN1(\IDinst/n7814 ), .DIN2(n1151), 
        .Q(\IDinst/n7818 ) );
  nnd2s1 \IDinst/U7856  ( .DIN1(\IDinst/n7816 ), .DIN2(\IDinst/n7815 ), 
        .Q(\IDinst/n7817 ) );
  nnd2s1 \IDinst/U7855  ( .DIN1(\IDinst/RegFile[3][20] ), .DIN2(n1071), 
        .Q(\IDinst/n7816 ) );
  nnd2s1 \IDinst/U7854  ( .DIN1(\IDinst/RegFile[2][20] ), .DIN2(n1060), 
        .Q(\IDinst/n7815 ) );
  nnd2s1 \IDinst/U7853  ( .DIN1(\IDinst/n7813 ), .DIN2(\IDinst/n7812 ), 
        .Q(\IDinst/n7814 ) );
  nnd2s1 \IDinst/U7852  ( .DIN1(\IDinst/RegFile[1][20] ), .DIN2(n1071), 
        .Q(\IDinst/n7813 ) );
  nnd2s1 \IDinst/U7851  ( .DIN1(\IDinst/RegFile[0][20] ), .DIN2(n1060), 
        .Q(\IDinst/n7812 ) );
  nnd2s1 \IDinst/U7850  ( .DIN1(\IDinst/n7811 ), .DIN2(n539), 
        .Q(\IDinst/n5986 ) );
  nnd2s1 \IDinst/U7849  ( .DIN1(\IDinst/n7766 ), .DIN2(n635), 
        .Q(\IDinst/n5987 ) );
  nnd2s1 \IDinst/U7848  ( .DIN1(\IDinst/n7810 ), .DIN2(\IDinst/n7809 ), 
        .Q(\IDinst/n7811 ) );
  nnd2s1 \IDinst/U7847  ( .DIN1(\IDinst/n7808 ), .DIN2(n643), 
        .Q(\IDinst/n7810 ) );
  nnd2s1 \IDinst/U7846  ( .DIN1(\IDinst/n7787 ), .DIN2(n670), 
        .Q(\IDinst/n7809 ) );
  nnd2s1 \IDinst/U7845  ( .DIN1(\IDinst/n7807 ), .DIN2(\IDinst/n7806 ), 
        .Q(\IDinst/n7808 ) );
  nnd2s1 \IDinst/U7844  ( .DIN1(\IDinst/n7805 ), .DIN2(n1196), 
        .Q(\IDinst/n7807 ) );
  nnd2s1 \IDinst/U7843  ( .DIN1(\IDinst/n7796 ), .DIN2(n1186), 
        .Q(\IDinst/n7806 ) );
  nnd2s1 \IDinst/U7842  ( .DIN1(\IDinst/n7804 ), .DIN2(\IDinst/n7803 ), 
        .Q(\IDinst/n7805 ) );
  nnd2s1 \IDinst/U7841  ( .DIN1(\IDinst/n7802 ), .DIN2(n1157), 
        .Q(\IDinst/n7804 ) );
  nnd2s1 \IDinst/U7840  ( .DIN1(\IDinst/n7799 ), .DIN2(n1150), 
        .Q(\IDinst/n7803 ) );
  nnd2s1 \IDinst/U7839  ( .DIN1(\IDinst/n7801 ), .DIN2(\IDinst/n7800 ), 
        .Q(\IDinst/n7802 ) );
  nnd2s1 \IDinst/U7838  ( .DIN1(\IDinst/RegFile[31][19] ), .DIN2(n1071), 
        .Q(\IDinst/n7801 ) );
  nnd2s1 \IDinst/U7837  ( .DIN1(\IDinst/RegFile[30][19] ), .DIN2(n1060), 
        .Q(\IDinst/n7800 ) );
  nnd2s1 \IDinst/U7836  ( .DIN1(\IDinst/n7798 ), .DIN2(\IDinst/n7797 ), 
        .Q(\IDinst/n7799 ) );
  nnd2s1 \IDinst/U7835  ( .DIN1(\IDinst/RegFile[29][19] ), .DIN2(n1071), 
        .Q(\IDinst/n7798 ) );
  nnd2s1 \IDinst/U7834  ( .DIN1(\IDinst/RegFile[28][19] ), .DIN2(n1059), 
        .Q(\IDinst/n7797 ) );
  nnd2s1 \IDinst/U7833  ( .DIN1(\IDinst/n7795 ), .DIN2(\IDinst/n7794 ), 
        .Q(\IDinst/n7796 ) );
  nnd2s1 \IDinst/U7832  ( .DIN1(\IDinst/n7793 ), .DIN2(n1157), 
        .Q(\IDinst/n7795 ) );
  nnd2s1 \IDinst/U7831  ( .DIN1(\IDinst/n7790 ), .DIN2(n1151), 
        .Q(\IDinst/n7794 ) );
  nnd2s1 \IDinst/U7830  ( .DIN1(\IDinst/n7792 ), .DIN2(\IDinst/n7791 ), 
        .Q(\IDinst/n7793 ) );
  nnd2s1 \IDinst/U7829  ( .DIN1(\IDinst/RegFile[27][19] ), .DIN2(n1071), 
        .Q(\IDinst/n7792 ) );
  nnd2s1 \IDinst/U7828  ( .DIN1(\IDinst/RegFile[26][19] ), .DIN2(n1059), 
        .Q(\IDinst/n7791 ) );
  nnd2s1 \IDinst/U7827  ( .DIN1(\IDinst/n7789 ), .DIN2(\IDinst/n7788 ), 
        .Q(\IDinst/n7790 ) );
  nnd2s1 \IDinst/U7826  ( .DIN1(\IDinst/RegFile[25][19] ), .DIN2(n1072), 
        .Q(\IDinst/n7789 ) );
  nnd2s1 \IDinst/U7825  ( .DIN1(\IDinst/RegFile[24][19] ), .DIN2(n1059), 
        .Q(\IDinst/n7788 ) );
  nnd2s1 \IDinst/U7824  ( .DIN1(\IDinst/n7786 ), .DIN2(\IDinst/n7785 ), 
        .Q(\IDinst/n7787 ) );
  nnd2s1 \IDinst/U7823  ( .DIN1(\IDinst/n7784 ), .DIN2(n1191), 
        .Q(\IDinst/n7786 ) );
  nnd2s1 \IDinst/U7822  ( .DIN1(\IDinst/n7775 ), .DIN2(n1186), 
        .Q(\IDinst/n7785 ) );
  nnd2s1 \IDinst/U7821  ( .DIN1(\IDinst/n7783 ), .DIN2(\IDinst/n7782 ), 
        .Q(\IDinst/n7784 ) );
  nnd2s1 \IDinst/U7820  ( .DIN1(\IDinst/n7781 ), .DIN2(n1157), 
        .Q(\IDinst/n7783 ) );
  nnd2s1 \IDinst/U7819  ( .DIN1(\IDinst/n7778 ), .DIN2(n1151), 
        .Q(\IDinst/n7782 ) );
  nnd2s1 \IDinst/U7818  ( .DIN1(\IDinst/n7780 ), .DIN2(\IDinst/n7779 ), 
        .Q(\IDinst/n7781 ) );
  nnd2s1 \IDinst/U7817  ( .DIN1(\IDinst/RegFile[23][19] ), .DIN2(n1072), 
        .Q(\IDinst/n7780 ) );
  nnd2s1 \IDinst/U7816  ( .DIN1(\IDinst/RegFile[22][19] ), .DIN2(n1059), 
        .Q(\IDinst/n7779 ) );
  nnd2s1 \IDinst/U7815  ( .DIN1(\IDinst/n7777 ), .DIN2(\IDinst/n7776 ), 
        .Q(\IDinst/n7778 ) );
  nnd2s1 \IDinst/U7814  ( .DIN1(\IDinst/RegFile[21][19] ), .DIN2(n1072), 
        .Q(\IDinst/n7777 ) );
  nnd2s1 \IDinst/U7813  ( .DIN1(\IDinst/RegFile[20][19] ), .DIN2(n1059), 
        .Q(\IDinst/n7776 ) );
  nnd2s1 \IDinst/U7812  ( .DIN1(\IDinst/n7774 ), .DIN2(\IDinst/n7773 ), 
        .Q(\IDinst/n7775 ) );
  nnd2s1 \IDinst/U7811  ( .DIN1(\IDinst/n7772 ), .DIN2(n1157), 
        .Q(\IDinst/n7774 ) );
  nnd2s1 \IDinst/U7810  ( .DIN1(\IDinst/n7769 ), .DIN2(n1151), 
        .Q(\IDinst/n7773 ) );
  nnd2s1 \IDinst/U7809  ( .DIN1(\IDinst/n7771 ), .DIN2(\IDinst/n7770 ), 
        .Q(\IDinst/n7772 ) );
  nnd2s1 \IDinst/U7808  ( .DIN1(\IDinst/RegFile[19][19] ), .DIN2(n1072), 
        .Q(\IDinst/n7771 ) );
  nnd2s1 \IDinst/U7807  ( .DIN1(\IDinst/RegFile[18][19] ), .DIN2(n1059), 
        .Q(\IDinst/n7770 ) );
  nnd2s1 \IDinst/U7806  ( .DIN1(\IDinst/n7768 ), .DIN2(\IDinst/n7767 ), 
        .Q(\IDinst/n7769 ) );
  nnd2s1 \IDinst/U7805  ( .DIN1(\IDinst/RegFile[17][19] ), .DIN2(n1072), 
        .Q(\IDinst/n7768 ) );
  nnd2s1 \IDinst/U7804  ( .DIN1(\IDinst/RegFile[16][19] ), .DIN2(n1059), 
        .Q(\IDinst/n7767 ) );
  nnd2s1 \IDinst/U7803  ( .DIN1(\IDinst/n7765 ), .DIN2(\IDinst/n7764 ), 
        .Q(\IDinst/n7766 ) );
  nnd2s1 \IDinst/U7802  ( .DIN1(\IDinst/n7763 ), .DIN2(n642), 
        .Q(\IDinst/n7765 ) );
  nnd2s1 \IDinst/U7801  ( .DIN1(\IDinst/n7742 ), .DIN2(n673), 
        .Q(\IDinst/n7764 ) );
  nnd2s1 \IDinst/U7800  ( .DIN1(\IDinst/n7762 ), .DIN2(\IDinst/n7761 ), 
        .Q(\IDinst/n7763 ) );
  nnd2s1 \IDinst/U7799  ( .DIN1(\IDinst/n7760 ), .DIN2(n1195), 
        .Q(\IDinst/n7762 ) );
  nnd2s1 \IDinst/U7798  ( .DIN1(\IDinst/n7751 ), .DIN2(n1186), 
        .Q(\IDinst/n7761 ) );
  nnd2s1 \IDinst/U7797  ( .DIN1(\IDinst/n7759 ), .DIN2(\IDinst/n7758 ), 
        .Q(\IDinst/n7760 ) );
  nnd2s1 \IDinst/U7796  ( .DIN1(\IDinst/n7757 ), .DIN2(n1157), 
        .Q(\IDinst/n7759 ) );
  nnd2s1 \IDinst/U7795  ( .DIN1(\IDinst/n7754 ), .DIN2(n1151), 
        .Q(\IDinst/n7758 ) );
  nnd2s1 \IDinst/U7794  ( .DIN1(\IDinst/n7756 ), .DIN2(\IDinst/n7755 ), 
        .Q(\IDinst/n7757 ) );
  nnd2s1 \IDinst/U7793  ( .DIN1(\IDinst/RegFile[15][19] ), .DIN2(n1072), 
        .Q(\IDinst/n7756 ) );
  nnd2s1 \IDinst/U7792  ( .DIN1(\IDinst/RegFile[14][19] ), .DIN2(n1059), 
        .Q(\IDinst/n7755 ) );
  nnd2s1 \IDinst/U7791  ( .DIN1(\IDinst/n7753 ), .DIN2(\IDinst/n7752 ), 
        .Q(\IDinst/n7754 ) );
  nnd2s1 \IDinst/U7790  ( .DIN1(\IDinst/RegFile[13][19] ), .DIN2(n1072), 
        .Q(\IDinst/n7753 ) );
  nnd2s1 \IDinst/U7789  ( .DIN1(\IDinst/RegFile[12][19] ), .DIN2(n1059), 
        .Q(\IDinst/n7752 ) );
  nnd2s1 \IDinst/U7788  ( .DIN1(\IDinst/n7750 ), .DIN2(\IDinst/n7749 ), 
        .Q(\IDinst/n7751 ) );
  nnd2s1 \IDinst/U7787  ( .DIN1(\IDinst/n7748 ), .DIN2(n1157), 
        .Q(\IDinst/n7750 ) );
  nnd2s1 \IDinst/U7786  ( .DIN1(\IDinst/n7745 ), .DIN2(n1151), 
        .Q(\IDinst/n7749 ) );
  nnd2s1 \IDinst/U7785  ( .DIN1(\IDinst/n7747 ), .DIN2(\IDinst/n7746 ), 
        .Q(\IDinst/n7748 ) );
  nnd2s1 \IDinst/U7784  ( .DIN1(\IDinst/RegFile[11][19] ), .DIN2(n1072), 
        .Q(\IDinst/n7747 ) );
  nnd2s1 \IDinst/U7783  ( .DIN1(\IDinst/RegFile[10][19] ), .DIN2(n1059), 
        .Q(\IDinst/n7746 ) );
  nnd2s1 \IDinst/U7782  ( .DIN1(\IDinst/n7744 ), .DIN2(\IDinst/n7743 ), 
        .Q(\IDinst/n7745 ) );
  nnd2s1 \IDinst/U7781  ( .DIN1(\IDinst/RegFile[9][19] ), .DIN2(n1072), 
        .Q(\IDinst/n7744 ) );
  nnd2s1 \IDinst/U7780  ( .DIN1(\IDinst/RegFile[8][19] ), .DIN2(n1059), 
        .Q(\IDinst/n7743 ) );
  nnd2s1 \IDinst/U7779  ( .DIN1(\IDinst/n7741 ), .DIN2(\IDinst/n7740 ), 
        .Q(\IDinst/n7742 ) );
  nnd2s1 \IDinst/U7778  ( .DIN1(\IDinst/n7739 ), .DIN2(n1193), 
        .Q(\IDinst/n7741 ) );
  nnd2s1 \IDinst/U7777  ( .DIN1(\IDinst/n7730 ), .DIN2(n1186), 
        .Q(\IDinst/n7740 ) );
  nnd2s1 \IDinst/U7776  ( .DIN1(\IDinst/n7738 ), .DIN2(\IDinst/n7737 ), 
        .Q(\IDinst/n7739 ) );
  nnd2s1 \IDinst/U7775  ( .DIN1(\IDinst/n7736 ), .DIN2(n1156), 
        .Q(\IDinst/n7738 ) );
  nnd2s1 \IDinst/U7774  ( .DIN1(\IDinst/n7733 ), .DIN2(n1151), 
        .Q(\IDinst/n7737 ) );
  nnd2s1 \IDinst/U7773  ( .DIN1(\IDinst/n7735 ), .DIN2(\IDinst/n7734 ), 
        .Q(\IDinst/n7736 ) );
  nnd2s1 \IDinst/U7772  ( .DIN1(\IDinst/RegFile[7][19] ), .DIN2(n1073), 
        .Q(\IDinst/n7735 ) );
  nnd2s1 \IDinst/U7771  ( .DIN1(\IDinst/RegFile[6][19] ), .DIN2(n1059), 
        .Q(\IDinst/n7734 ) );
  nnd2s1 \IDinst/U7770  ( .DIN1(\IDinst/n7732 ), .DIN2(\IDinst/n7731 ), 
        .Q(\IDinst/n7733 ) );
  nnd2s1 \IDinst/U7769  ( .DIN1(\IDinst/RegFile[5][19] ), .DIN2(n1073), 
        .Q(\IDinst/n7732 ) );
  nnd2s1 \IDinst/U7768  ( .DIN1(\IDinst/RegFile[4][19] ), .DIN2(n1059), 
        .Q(\IDinst/n7731 ) );
  nnd2s1 \IDinst/U7767  ( .DIN1(\IDinst/n7729 ), .DIN2(\IDinst/n7728 ), 
        .Q(\IDinst/n7730 ) );
  nnd2s1 \IDinst/U7766  ( .DIN1(\IDinst/n7727 ), .DIN2(n1156), 
        .Q(\IDinst/n7729 ) );
  nnd2s1 \IDinst/U7765  ( .DIN1(\IDinst/n7724 ), .DIN2(n1151), 
        .Q(\IDinst/n7728 ) );
  nnd2s1 \IDinst/U7764  ( .DIN1(\IDinst/n7726 ), .DIN2(\IDinst/n7725 ), 
        .Q(\IDinst/n7727 ) );
  nnd2s1 \IDinst/U7763  ( .DIN1(\IDinst/RegFile[3][19] ), .DIN2(n1073), 
        .Q(\IDinst/n7726 ) );
  nnd2s1 \IDinst/U7762  ( .DIN1(\IDinst/RegFile[2][19] ), .DIN2(n1058), 
        .Q(\IDinst/n7725 ) );
  nnd2s1 \IDinst/U7761  ( .DIN1(\IDinst/n7723 ), .DIN2(\IDinst/n7722 ), 
        .Q(\IDinst/n7724 ) );
  nnd2s1 \IDinst/U7760  ( .DIN1(\IDinst/RegFile[1][19] ), .DIN2(n1073), 
        .Q(\IDinst/n7723 ) );
  nnd2s1 \IDinst/U7759  ( .DIN1(\IDinst/RegFile[0][19] ), .DIN2(n1058), 
        .Q(\IDinst/n7722 ) );
  nnd2s1 \IDinst/U7758  ( .DIN1(\IDinst/n7721 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n5984 ) );
  nnd2s1 \IDinst/U7757  ( .DIN1(\IDinst/n7676 ), .DIN2(n636), 
        .Q(\IDinst/n5985 ) );
  nnd2s1 \IDinst/U7756  ( .DIN1(\IDinst/n7720 ), .DIN2(\IDinst/n7719 ), 
        .Q(\IDinst/n7721 ) );
  nnd2s1 \IDinst/U7755  ( .DIN1(\IDinst/n7718 ), .DIN2(n641), 
        .Q(\IDinst/n7720 ) );
  nnd2s1 \IDinst/U7754  ( .DIN1(\IDinst/n7697 ), .DIN2(n671), 
        .Q(\IDinst/n7719 ) );
  nnd2s1 \IDinst/U7753  ( .DIN1(\IDinst/n7717 ), .DIN2(\IDinst/n7716 ), 
        .Q(\IDinst/n7718 ) );
  nnd2s1 \IDinst/U7752  ( .DIN1(\IDinst/n7715 ), .DIN2(n1192), 
        .Q(\IDinst/n7717 ) );
  nnd2s1 \IDinst/U7751  ( .DIN1(\IDinst/n7706 ), .DIN2(n1186), 
        .Q(\IDinst/n7716 ) );
  nnd2s1 \IDinst/U7750  ( .DIN1(\IDinst/n7714 ), .DIN2(\IDinst/n7713 ), 
        .Q(\IDinst/n7715 ) );
  nnd2s1 \IDinst/U7749  ( .DIN1(\IDinst/n7712 ), .DIN2(n1156), 
        .Q(\IDinst/n7714 ) );
  nnd2s1 \IDinst/U7748  ( .DIN1(\IDinst/n7709 ), .DIN2(n1151), 
        .Q(\IDinst/n7713 ) );
  nnd2s1 \IDinst/U7747  ( .DIN1(\IDinst/n7711 ), .DIN2(\IDinst/n7710 ), 
        .Q(\IDinst/n7712 ) );
  nnd2s1 \IDinst/U7746  ( .DIN1(\IDinst/RegFile[31][18] ), .DIN2(n1073), 
        .Q(\IDinst/n7711 ) );
  nnd2s1 \IDinst/U7745  ( .DIN1(\IDinst/RegFile[30][18] ), .DIN2(n1058), 
        .Q(\IDinst/n7710 ) );
  nnd2s1 \IDinst/U7744  ( .DIN1(\IDinst/n7708 ), .DIN2(\IDinst/n7707 ), 
        .Q(\IDinst/n7709 ) );
  nnd2s1 \IDinst/U7743  ( .DIN1(\IDinst/RegFile[29][18] ), .DIN2(n1073), 
        .Q(\IDinst/n7708 ) );
  nnd2s1 \IDinst/U7742  ( .DIN1(\IDinst/RegFile[28][18] ), .DIN2(n1058), 
        .Q(\IDinst/n7707 ) );
  nnd2s1 \IDinst/U7741  ( .DIN1(\IDinst/n7705 ), .DIN2(\IDinst/n7704 ), 
        .Q(\IDinst/n7706 ) );
  nnd2s1 \IDinst/U7740  ( .DIN1(\IDinst/n7703 ), .DIN2(n1156), 
        .Q(\IDinst/n7705 ) );
  nnd2s1 \IDinst/U7739  ( .DIN1(\IDinst/n7700 ), .DIN2(n1151), 
        .Q(\IDinst/n7704 ) );
  nnd2s1 \IDinst/U7738  ( .DIN1(\IDinst/n7702 ), .DIN2(\IDinst/n7701 ), 
        .Q(\IDinst/n7703 ) );
  nnd2s1 \IDinst/U7737  ( .DIN1(\IDinst/RegFile[27][18] ), .DIN2(n1073), 
        .Q(\IDinst/n7702 ) );
  nnd2s1 \IDinst/U7736  ( .DIN1(\IDinst/RegFile[26][18] ), .DIN2(n1058), 
        .Q(\IDinst/n7701 ) );
  nnd2s1 \IDinst/U7735  ( .DIN1(\IDinst/n7699 ), .DIN2(\IDinst/n7698 ), 
        .Q(\IDinst/n7700 ) );
  nnd2s1 \IDinst/U7734  ( .DIN1(\IDinst/RegFile[25][18] ), .DIN2(n1073), 
        .Q(\IDinst/n7699 ) );
  nnd2s1 \IDinst/U7733  ( .DIN1(\IDinst/RegFile[24][18] ), .DIN2(n1058), 
        .Q(\IDinst/n7698 ) );
  nnd2s1 \IDinst/U7732  ( .DIN1(\IDinst/n7696 ), .DIN2(\IDinst/n7695 ), 
        .Q(\IDinst/n7697 ) );
  nnd2s1 \IDinst/U7731  ( .DIN1(\IDinst/n7694 ), .DIN2(n1190), 
        .Q(\IDinst/n7696 ) );
  nnd2s1 \IDinst/U7730  ( .DIN1(\IDinst/n7685 ), .DIN2(n1186), 
        .Q(\IDinst/n7695 ) );
  nnd2s1 \IDinst/U7729  ( .DIN1(\IDinst/n7693 ), .DIN2(\IDinst/n7692 ), 
        .Q(\IDinst/n7694 ) );
  nnd2s1 \IDinst/U7728  ( .DIN1(\IDinst/n7691 ), .DIN2(n1156), 
        .Q(\IDinst/n7693 ) );
  nnd2s1 \IDinst/U7727  ( .DIN1(\IDinst/n7688 ), .DIN2(n1151), 
        .Q(\IDinst/n7692 ) );
  nnd2s1 \IDinst/U7726  ( .DIN1(\IDinst/n7690 ), .DIN2(\IDinst/n7689 ), 
        .Q(\IDinst/n7691 ) );
  nnd2s1 \IDinst/U7725  ( .DIN1(\IDinst/RegFile[23][18] ), .DIN2(n1074), 
        .Q(\IDinst/n7690 ) );
  nnd2s1 \IDinst/U7724  ( .DIN1(\IDinst/RegFile[22][18] ), .DIN2(n1058), 
        .Q(\IDinst/n7689 ) );
  nnd2s1 \IDinst/U7723  ( .DIN1(\IDinst/n7687 ), .DIN2(\IDinst/n7686 ), 
        .Q(\IDinst/n7688 ) );
  nnd2s1 \IDinst/U7722  ( .DIN1(\IDinst/RegFile[21][18] ), .DIN2(n1074), 
        .Q(\IDinst/n7687 ) );
  nnd2s1 \IDinst/U7721  ( .DIN1(\IDinst/RegFile[20][18] ), .DIN2(n1058), 
        .Q(\IDinst/n7686 ) );
  nnd2s1 \IDinst/U7720  ( .DIN1(\IDinst/n7684 ), .DIN2(\IDinst/n7683 ), 
        .Q(\IDinst/n7685 ) );
  nnd2s1 \IDinst/U7719  ( .DIN1(\IDinst/n7682 ), .DIN2(n1156), 
        .Q(\IDinst/n7684 ) );
  nnd2s1 \IDinst/U7718  ( .DIN1(\IDinst/n7679 ), .DIN2(n1151), 
        .Q(\IDinst/n7683 ) );
  nnd2s1 \IDinst/U7717  ( .DIN1(\IDinst/n7681 ), .DIN2(\IDinst/n7680 ), 
        .Q(\IDinst/n7682 ) );
  nnd2s1 \IDinst/U7716  ( .DIN1(\IDinst/RegFile[19][18] ), .DIN2(n1074), 
        .Q(\IDinst/n7681 ) );
  nnd2s1 \IDinst/U7715  ( .DIN1(\IDinst/RegFile[18][18] ), .DIN2(n1058), 
        .Q(\IDinst/n7680 ) );
  nnd2s1 \IDinst/U7714  ( .DIN1(\IDinst/n7678 ), .DIN2(\IDinst/n7677 ), 
        .Q(\IDinst/n7679 ) );
  nnd2s1 \IDinst/U7713  ( .DIN1(\IDinst/RegFile[17][18] ), .DIN2(n1074), 
        .Q(\IDinst/n7678 ) );
  nnd2s1 \IDinst/U7712  ( .DIN1(\IDinst/RegFile[16][18] ), .DIN2(n1058), 
        .Q(\IDinst/n7677 ) );
  nnd2s1 \IDinst/U7711  ( .DIN1(\IDinst/n7675 ), .DIN2(\IDinst/n7674 ), 
        .Q(\IDinst/n7676 ) );
  nnd2s1 \IDinst/U7710  ( .DIN1(\IDinst/n7673 ), .DIN2(n644), 
        .Q(\IDinst/n7675 ) );
  nnd2s1 \IDinst/U7709  ( .DIN1(\IDinst/n7652 ), .DIN2(n672), 
        .Q(\IDinst/n7674 ) );
  nnd2s1 \IDinst/U7708  ( .DIN1(\IDinst/n7672 ), .DIN2(\IDinst/n7671 ), 
        .Q(\IDinst/n7673 ) );
  nnd2s1 \IDinst/U7707  ( .DIN1(\IDinst/n7670 ), .DIN2(n1194), 
        .Q(\IDinst/n7672 ) );
  nnd2s1 \IDinst/U7706  ( .DIN1(\IDinst/n7661 ), .DIN2(n1186), 
        .Q(\IDinst/n7671 ) );
  nnd2s1 \IDinst/U7705  ( .DIN1(\IDinst/n7669 ), .DIN2(\IDinst/n7668 ), 
        .Q(\IDinst/n7670 ) );
  nnd2s1 \IDinst/U7704  ( .DIN1(\IDinst/n7667 ), .DIN2(n1156), 
        .Q(\IDinst/n7669 ) );
  nnd2s1 \IDinst/U7703  ( .DIN1(\IDinst/n7664 ), .DIN2(n1151), 
        .Q(\IDinst/n7668 ) );
  nnd2s1 \IDinst/U7702  ( .DIN1(\IDinst/n7666 ), .DIN2(\IDinst/n7665 ), 
        .Q(\IDinst/n7667 ) );
  nnd2s1 \IDinst/U7701  ( .DIN1(\IDinst/RegFile[15][18] ), .DIN2(n1074), 
        .Q(\IDinst/n7666 ) );
  nnd2s1 \IDinst/U7700  ( .DIN1(\IDinst/RegFile[14][18] ), .DIN2(n1058), 
        .Q(\IDinst/n7665 ) );
  nnd2s1 \IDinst/U7699  ( .DIN1(\IDinst/n7663 ), .DIN2(\IDinst/n7662 ), 
        .Q(\IDinst/n7664 ) );
  nnd2s1 \IDinst/U7698  ( .DIN1(\IDinst/RegFile[13][18] ), .DIN2(n1074), 
        .Q(\IDinst/n7663 ) );
  nnd2s1 \IDinst/U7697  ( .DIN1(\IDinst/RegFile[12][18] ), .DIN2(n1058), 
        .Q(\IDinst/n7662 ) );
  nnd2s1 \IDinst/U7696  ( .DIN1(\IDinst/n7660 ), .DIN2(\IDinst/n7659 ), 
        .Q(\IDinst/n7661 ) );
  nnd2s1 \IDinst/U7695  ( .DIN1(\IDinst/n7658 ), .DIN2(n1156), 
        .Q(\IDinst/n7660 ) );
  nnd2s1 \IDinst/U7694  ( .DIN1(\IDinst/n7655 ), .DIN2(n1152), 
        .Q(\IDinst/n7659 ) );
  nnd2s1 \IDinst/U7693  ( .DIN1(\IDinst/n7657 ), .DIN2(\IDinst/n7656 ), 
        .Q(\IDinst/n7658 ) );
  nnd2s1 \IDinst/U7692  ( .DIN1(\IDinst/RegFile[11][18] ), .DIN2(n1074), 
        .Q(\IDinst/n7657 ) );
  nnd2s1 \IDinst/U7691  ( .DIN1(\IDinst/RegFile[10][18] ), .DIN2(n1058), 
        .Q(\IDinst/n7656 ) );
  nnd2s1 \IDinst/U7690  ( .DIN1(\IDinst/n7654 ), .DIN2(\IDinst/n7653 ), 
        .Q(\IDinst/n7655 ) );
  nnd2s1 \IDinst/U7689  ( .DIN1(\IDinst/RegFile[9][18] ), .DIN2(n1074), 
        .Q(\IDinst/n7654 ) );
  nnd2s1 \IDinst/U7688  ( .DIN1(\IDinst/RegFile[8][18] ), .DIN2(n1057), 
        .Q(\IDinst/n7653 ) );
  nnd2s1 \IDinst/U7687  ( .DIN1(\IDinst/n7651 ), .DIN2(\IDinst/n7650 ), 
        .Q(\IDinst/n7652 ) );
  nnd2s1 \IDinst/U7686  ( .DIN1(\IDinst/n7649 ), .DIN2(n1197), 
        .Q(\IDinst/n7651 ) );
  nnd2s1 \IDinst/U7685  ( .DIN1(\IDinst/n7640 ), .DIN2(n1186), 
        .Q(\IDinst/n7650 ) );
  nnd2s1 \IDinst/U7684  ( .DIN1(\IDinst/n7648 ), .DIN2(\IDinst/n7647 ), 
        .Q(\IDinst/n7649 ) );
  nnd2s1 \IDinst/U7683  ( .DIN1(\IDinst/n7646 ), .DIN2(n1156), 
        .Q(\IDinst/n7648 ) );
  nnd2s1 \IDinst/U7682  ( .DIN1(\IDinst/n7643 ), .DIN2(n1152), 
        .Q(\IDinst/n7647 ) );
  nnd2s1 \IDinst/U7681  ( .DIN1(\IDinst/n7645 ), .DIN2(\IDinst/n7644 ), 
        .Q(\IDinst/n7646 ) );
  nnd2s1 \IDinst/U7680  ( .DIN1(\IDinst/RegFile[7][18] ), .DIN2(n1074), 
        .Q(\IDinst/n7645 ) );
  nnd2s1 \IDinst/U7679  ( .DIN1(\IDinst/RegFile[6][18] ), .DIN2(n1057), 
        .Q(\IDinst/n7644 ) );
  nnd2s1 \IDinst/U7678  ( .DIN1(\IDinst/n7642 ), .DIN2(\IDinst/n7641 ), 
        .Q(\IDinst/n7643 ) );
  nnd2s1 \IDinst/U7677  ( .DIN1(\IDinst/RegFile[5][18] ), .DIN2(n1075), 
        .Q(\IDinst/n7642 ) );
  nnd2s1 \IDinst/U7676  ( .DIN1(\IDinst/RegFile[4][18] ), .DIN2(n1057), 
        .Q(\IDinst/n7641 ) );
  nnd2s1 \IDinst/U7675  ( .DIN1(\IDinst/n7639 ), .DIN2(\IDinst/n7638 ), 
        .Q(\IDinst/n7640 ) );
  nnd2s1 \IDinst/U7674  ( .DIN1(\IDinst/n7637 ), .DIN2(n1155), 
        .Q(\IDinst/n7639 ) );
  nnd2s1 \IDinst/U7673  ( .DIN1(\IDinst/n7634 ), .DIN2(n1152), 
        .Q(\IDinst/n7638 ) );
  nnd2s1 \IDinst/U7672  ( .DIN1(\IDinst/n7636 ), .DIN2(\IDinst/n7635 ), 
        .Q(\IDinst/n7637 ) );
  nnd2s1 \IDinst/U7671  ( .DIN1(\IDinst/RegFile[3][18] ), .DIN2(n1075), 
        .Q(\IDinst/n7636 ) );
  nnd2s1 \IDinst/U7670  ( .DIN1(\IDinst/RegFile[2][18] ), .DIN2(n1057), 
        .Q(\IDinst/n7635 ) );
  nnd2s1 \IDinst/U7669  ( .DIN1(\IDinst/n7633 ), .DIN2(\IDinst/n7632 ), 
        .Q(\IDinst/n7634 ) );
  nnd2s1 \IDinst/U7668  ( .DIN1(\IDinst/RegFile[1][18] ), .DIN2(n1075), 
        .Q(\IDinst/n7633 ) );
  nnd2s1 \IDinst/U7667  ( .DIN1(\IDinst/RegFile[0][18] ), .DIN2(n1057), 
        .Q(\IDinst/n7632 ) );
  nnd2s1 \IDinst/U7666  ( .DIN1(\IDinst/n7631 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n5982 ) );
  nnd2s1 \IDinst/U7665  ( .DIN1(\IDinst/n7586 ), .DIN2(n635), 
        .Q(\IDinst/n5983 ) );
  nnd2s1 \IDinst/U7664  ( .DIN1(\IDinst/n7630 ), .DIN2(\IDinst/n7629 ), 
        .Q(\IDinst/n7631 ) );
  nnd2s1 \IDinst/U7663  ( .DIN1(\IDinst/n7628 ), .DIN2(n643), 
        .Q(\IDinst/n7630 ) );
  nnd2s1 \IDinst/U7662  ( .DIN1(\IDinst/n7607 ), .DIN2(n670), 
        .Q(\IDinst/n7629 ) );
  nnd2s1 \IDinst/U7661  ( .DIN1(\IDinst/n7627 ), .DIN2(\IDinst/n7626 ), 
        .Q(\IDinst/n7628 ) );
  nnd2s1 \IDinst/U7660  ( .DIN1(\IDinst/n7625 ), .DIN2(n1192), 
        .Q(\IDinst/n7627 ) );
  nnd2s1 \IDinst/U7659  ( .DIN1(\IDinst/n7616 ), .DIN2(n1186), 
        .Q(\IDinst/n7626 ) );
  nnd2s1 \IDinst/U7658  ( .DIN1(\IDinst/n7624 ), .DIN2(\IDinst/n7623 ), 
        .Q(\IDinst/n7625 ) );
  nnd2s1 \IDinst/U7657  ( .DIN1(\IDinst/n7622 ), .DIN2(n1155), 
        .Q(\IDinst/n7624 ) );
  nnd2s1 \IDinst/U7656  ( .DIN1(\IDinst/n7619 ), .DIN2(n1152), 
        .Q(\IDinst/n7623 ) );
  nnd2s1 \IDinst/U7655  ( .DIN1(\IDinst/n7621 ), .DIN2(\IDinst/n7620 ), 
        .Q(\IDinst/n7622 ) );
  nnd2s1 \IDinst/U7654  ( .DIN1(\IDinst/RegFile[31][17] ), .DIN2(n1075), 
        .Q(\IDinst/n7621 ) );
  nnd2s1 \IDinst/U7653  ( .DIN1(\IDinst/RegFile[30][17] ), .DIN2(n1057), 
        .Q(\IDinst/n7620 ) );
  nnd2s1 \IDinst/U7652  ( .DIN1(\IDinst/n7618 ), .DIN2(\IDinst/n7617 ), 
        .Q(\IDinst/n7619 ) );
  nnd2s1 \IDinst/U7651  ( .DIN1(\IDinst/RegFile[29][17] ), .DIN2(n1075), 
        .Q(\IDinst/n7618 ) );
  nnd2s1 \IDinst/U7650  ( .DIN1(\IDinst/RegFile[28][17] ), .DIN2(n1057), 
        .Q(\IDinst/n7617 ) );
  nnd2s1 \IDinst/U7649  ( .DIN1(\IDinst/n7615 ), .DIN2(\IDinst/n7614 ), 
        .Q(\IDinst/n7616 ) );
  nnd2s1 \IDinst/U7648  ( .DIN1(\IDinst/n7613 ), .DIN2(n1155), 
        .Q(\IDinst/n7615 ) );
  nnd2s1 \IDinst/U7647  ( .DIN1(\IDinst/n7610 ), .DIN2(n1152), 
        .Q(\IDinst/n7614 ) );
  nnd2s1 \IDinst/U7646  ( .DIN1(\IDinst/n7612 ), .DIN2(\IDinst/n7611 ), 
        .Q(\IDinst/n7613 ) );
  nnd2s1 \IDinst/U7645  ( .DIN1(\IDinst/RegFile[27][17] ), .DIN2(n1075), 
        .Q(\IDinst/n7612 ) );
  nnd2s1 \IDinst/U7644  ( .DIN1(\IDinst/RegFile[26][17] ), .DIN2(n1057), 
        .Q(\IDinst/n7611 ) );
  nnd2s1 \IDinst/U7643  ( .DIN1(\IDinst/n7609 ), .DIN2(\IDinst/n7608 ), 
        .Q(\IDinst/n7610 ) );
  nnd2s1 \IDinst/U7642  ( .DIN1(\IDinst/RegFile[25][17] ), .DIN2(n1075), 
        .Q(\IDinst/n7609 ) );
  nnd2s1 \IDinst/U7641  ( .DIN1(\IDinst/RegFile[24][17] ), .DIN2(n1057), 
        .Q(\IDinst/n7608 ) );
  nnd2s1 \IDinst/U7640  ( .DIN1(\IDinst/n7606 ), .DIN2(\IDinst/n7605 ), 
        .Q(\IDinst/n7607 ) );
  nnd2s1 \IDinst/U7639  ( .DIN1(\IDinst/n7604 ), .DIN2(n1192), 
        .Q(\IDinst/n7606 ) );
  nnd2s1 \IDinst/U7638  ( .DIN1(\IDinst/n7595 ), .DIN2(n1186), 
        .Q(\IDinst/n7605 ) );
  nnd2s1 \IDinst/U7637  ( .DIN1(\IDinst/n7603 ), .DIN2(\IDinst/n7602 ), 
        .Q(\IDinst/n7604 ) );
  nnd2s1 \IDinst/U7636  ( .DIN1(\IDinst/n7601 ), .DIN2(n1155), 
        .Q(\IDinst/n7603 ) );
  nnd2s1 \IDinst/U7635  ( .DIN1(\IDinst/n7598 ), .DIN2(n1152), 
        .Q(\IDinst/n7602 ) );
  nnd2s1 \IDinst/U7634  ( .DIN1(\IDinst/n7600 ), .DIN2(\IDinst/n7599 ), 
        .Q(\IDinst/n7601 ) );
  nnd2s1 \IDinst/U7633  ( .DIN1(\IDinst/RegFile[23][17] ), .DIN2(n1075), 
        .Q(\IDinst/n7600 ) );
  nnd2s1 \IDinst/U7632  ( .DIN1(\IDinst/RegFile[22][17] ), .DIN2(n1057), 
        .Q(\IDinst/n7599 ) );
  nnd2s1 \IDinst/U7631  ( .DIN1(\IDinst/n7597 ), .DIN2(\IDinst/n7596 ), 
        .Q(\IDinst/n7598 ) );
  nnd2s1 \IDinst/U7630  ( .DIN1(\IDinst/RegFile[21][17] ), .DIN2(n1075), 
        .Q(\IDinst/n7597 ) );
  nnd2s1 \IDinst/U7629  ( .DIN1(\IDinst/RegFile[20][17] ), .DIN2(n1057), 
        .Q(\IDinst/n7596 ) );
  nnd2s1 \IDinst/U7628  ( .DIN1(\IDinst/n7594 ), .DIN2(\IDinst/n7593 ), 
        .Q(\IDinst/n7595 ) );
  nnd2s1 \IDinst/U7627  ( .DIN1(\IDinst/n7592 ), .DIN2(n1155), 
        .Q(\IDinst/n7594 ) );
  nnd2s1 \IDinst/U7626  ( .DIN1(\IDinst/n7589 ), .DIN2(n1152), 
        .Q(\IDinst/n7593 ) );
  nnd2s1 \IDinst/U7625  ( .DIN1(\IDinst/n7591 ), .DIN2(\IDinst/n7590 ), 
        .Q(\IDinst/n7592 ) );
  nnd2s1 \IDinst/U7624  ( .DIN1(\IDinst/RegFile[19][17] ), .DIN2(n1076), 
        .Q(\IDinst/n7591 ) );
  nnd2s1 \IDinst/U7623  ( .DIN1(\IDinst/RegFile[18][17] ), .DIN2(n1057), 
        .Q(\IDinst/n7590 ) );
  nnd2s1 \IDinst/U7622  ( .DIN1(\IDinst/n7588 ), .DIN2(\IDinst/n7587 ), 
        .Q(\IDinst/n7589 ) );
  nnd2s1 \IDinst/U7621  ( .DIN1(\IDinst/RegFile[17][17] ), .DIN2(n1076), 
        .Q(\IDinst/n7588 ) );
  nnd2s1 \IDinst/U7620  ( .DIN1(\IDinst/RegFile[16][17] ), .DIN2(n1057), 
        .Q(\IDinst/n7587 ) );
  nnd2s1 \IDinst/U7619  ( .DIN1(\IDinst/n7585 ), .DIN2(\IDinst/n7584 ), 
        .Q(\IDinst/n7586 ) );
  nnd2s1 \IDinst/U7618  ( .DIN1(\IDinst/n7583 ), .DIN2(n642), 
        .Q(\IDinst/n7585 ) );
  nnd2s1 \IDinst/U7617  ( .DIN1(\IDinst/n7562 ), .DIN2(n673), 
        .Q(\IDinst/n7584 ) );
  nnd2s1 \IDinst/U7616  ( .DIN1(\IDinst/n7582 ), .DIN2(\IDinst/n7581 ), 
        .Q(\IDinst/n7583 ) );
  nnd2s1 \IDinst/U7615  ( .DIN1(\IDinst/n7580 ), .DIN2(n1192), 
        .Q(\IDinst/n7582 ) );
  nnd2s1 \IDinst/U7614  ( .DIN1(\IDinst/n7571 ), .DIN2(n1185), 
        .Q(\IDinst/n7581 ) );
  nnd2s1 \IDinst/U7613  ( .DIN1(\IDinst/n7579 ), .DIN2(\IDinst/n7578 ), 
        .Q(\IDinst/n7580 ) );
  nnd2s1 \IDinst/U7612  ( .DIN1(\IDinst/n7577 ), .DIN2(n1155), 
        .Q(\IDinst/n7579 ) );
  nnd2s1 \IDinst/U7611  ( .DIN1(\IDinst/n7574 ), .DIN2(n1152), 
        .Q(\IDinst/n7578 ) );
  nnd2s1 \IDinst/U7610  ( .DIN1(\IDinst/n7576 ), .DIN2(\IDinst/n7575 ), 
        .Q(\IDinst/n7577 ) );
  nnd2s1 \IDinst/U7609  ( .DIN1(\IDinst/RegFile[15][17] ), .DIN2(n1076), 
        .Q(\IDinst/n7576 ) );
  nnd2s1 \IDinst/U7608  ( .DIN1(\IDinst/RegFile[14][17] ), .DIN2(n1056), 
        .Q(\IDinst/n7575 ) );
  nnd2s1 \IDinst/U7607  ( .DIN1(\IDinst/n7573 ), .DIN2(\IDinst/n7572 ), 
        .Q(\IDinst/n7574 ) );
  nnd2s1 \IDinst/U7606  ( .DIN1(\IDinst/RegFile[13][17] ), .DIN2(n1076), 
        .Q(\IDinst/n7573 ) );
  nnd2s1 \IDinst/U7605  ( .DIN1(\IDinst/RegFile[12][17] ), .DIN2(n1056), 
        .Q(\IDinst/n7572 ) );
  nnd2s1 \IDinst/U7604  ( .DIN1(\IDinst/n7570 ), .DIN2(\IDinst/n7569 ), 
        .Q(\IDinst/n7571 ) );
  nnd2s1 \IDinst/U7603  ( .DIN1(\IDinst/n7568 ), .DIN2(n1155), 
        .Q(\IDinst/n7570 ) );
  nnd2s1 \IDinst/U7602  ( .DIN1(\IDinst/n7565 ), .DIN2(n1152), 
        .Q(\IDinst/n7569 ) );
  nnd2s1 \IDinst/U7601  ( .DIN1(\IDinst/n7567 ), .DIN2(\IDinst/n7566 ), 
        .Q(\IDinst/n7568 ) );
  nnd2s1 \IDinst/U7600  ( .DIN1(\IDinst/RegFile[11][17] ), .DIN2(n1076), 
        .Q(\IDinst/n7567 ) );
  nnd2s1 \IDinst/U7599  ( .DIN1(\IDinst/RegFile[10][17] ), .DIN2(n1056), 
        .Q(\IDinst/n7566 ) );
  nnd2s1 \IDinst/U7598  ( .DIN1(\IDinst/n7564 ), .DIN2(\IDinst/n7563 ), 
        .Q(\IDinst/n7565 ) );
  nnd2s1 \IDinst/U7597  ( .DIN1(\IDinst/RegFile[9][17] ), .DIN2(n1076), 
        .Q(\IDinst/n7564 ) );
  nnd2s1 \IDinst/U7596  ( .DIN1(\IDinst/RegFile[8][17] ), .DIN2(n1056), 
        .Q(\IDinst/n7563 ) );
  nnd2s1 \IDinst/U7595  ( .DIN1(\IDinst/n7561 ), .DIN2(\IDinst/n7560 ), 
        .Q(\IDinst/n7562 ) );
  nnd2s1 \IDinst/U7594  ( .DIN1(\IDinst/n7559 ), .DIN2(n1192), 
        .Q(\IDinst/n7561 ) );
  nnd2s1 \IDinst/U7593  ( .DIN1(\IDinst/n7550 ), .DIN2(n1185), 
        .Q(\IDinst/n7560 ) );
  nnd2s1 \IDinst/U7592  ( .DIN1(\IDinst/n7558 ), .DIN2(\IDinst/n7557 ), 
        .Q(\IDinst/n7559 ) );
  nnd2s1 \IDinst/U7591  ( .DIN1(\IDinst/n7556 ), .DIN2(n1155), 
        .Q(\IDinst/n7558 ) );
  nnd2s1 \IDinst/U7590  ( .DIN1(\IDinst/n7553 ), .DIN2(n1152), 
        .Q(\IDinst/n7557 ) );
  nnd2s1 \IDinst/U7589  ( .DIN1(\IDinst/n7555 ), .DIN2(\IDinst/n7554 ), 
        .Q(\IDinst/n7556 ) );
  nnd2s1 \IDinst/U7588  ( .DIN1(\IDinst/RegFile[7][17] ), .DIN2(n1076), 
        .Q(\IDinst/n7555 ) );
  nnd2s1 \IDinst/U7587  ( .DIN1(\IDinst/RegFile[6][17] ), .DIN2(n1056), 
        .Q(\IDinst/n7554 ) );
  nnd2s1 \IDinst/U7586  ( .DIN1(\IDinst/n7552 ), .DIN2(\IDinst/n7551 ), 
        .Q(\IDinst/n7553 ) );
  nnd2s1 \IDinst/U7585  ( .DIN1(\IDinst/RegFile[5][17] ), .DIN2(n1076), 
        .Q(\IDinst/n7552 ) );
  nnd2s1 \IDinst/U7584  ( .DIN1(\IDinst/RegFile[4][17] ), .DIN2(n1056), 
        .Q(\IDinst/n7551 ) );
  nnd2s1 \IDinst/U7583  ( .DIN1(\IDinst/n7549 ), .DIN2(\IDinst/n7548 ), 
        .Q(\IDinst/n7550 ) );
  nnd2s1 \IDinst/U7582  ( .DIN1(\IDinst/n7547 ), .DIN2(n1154), 
        .Q(\IDinst/n7549 ) );
  nnd2s1 \IDinst/U7581  ( .DIN1(\IDinst/n7544 ), .DIN2(n1152), 
        .Q(\IDinst/n7548 ) );
  nnd2s1 \IDinst/U7580  ( .DIN1(\IDinst/n7546 ), .DIN2(\IDinst/n7545 ), 
        .Q(\IDinst/n7547 ) );
  nnd2s1 \IDinst/U7579  ( .DIN1(\IDinst/RegFile[3][17] ), .DIN2(n1076), 
        .Q(\IDinst/n7546 ) );
  nnd2s1 \IDinst/U7578  ( .DIN1(\IDinst/RegFile[2][17] ), .DIN2(n1056), 
        .Q(\IDinst/n7545 ) );
  nnd2s1 \IDinst/U7577  ( .DIN1(\IDinst/n7543 ), .DIN2(\IDinst/n7542 ), 
        .Q(\IDinst/n7544 ) );
  nnd2s1 \IDinst/U7576  ( .DIN1(\IDinst/RegFile[1][17] ), .DIN2(n1077), 
        .Q(\IDinst/n7543 ) );
  nnd2s1 \IDinst/U7575  ( .DIN1(\IDinst/RegFile[0][17] ), .DIN2(n1056), 
        .Q(\IDinst/n7542 ) );
  nnd2s1 \IDinst/U7574  ( .DIN1(\IDinst/n7541 ), .DIN2(n539), 
        .Q(\IDinst/n5980 ) );
  nnd2s1 \IDinst/U7573  ( .DIN1(\IDinst/n7496 ), .DIN2(n636), 
        .Q(\IDinst/n5981 ) );
  nnd2s1 \IDinst/U7572  ( .DIN1(\IDinst/n7540 ), .DIN2(\IDinst/n7539 ), 
        .Q(\IDinst/n7541 ) );
  nnd2s1 \IDinst/U7571  ( .DIN1(\IDinst/n7538 ), .DIN2(n641), 
        .Q(\IDinst/n7540 ) );
  nnd2s1 \IDinst/U7570  ( .DIN1(\IDinst/n7517 ), .DIN2(n671), 
        .Q(\IDinst/n7539 ) );
  nnd2s1 \IDinst/U7569  ( .DIN1(\IDinst/n7537 ), .DIN2(\IDinst/n7536 ), 
        .Q(\IDinst/n7538 ) );
  nnd2s1 \IDinst/U7568  ( .DIN1(\IDinst/n7535 ), .DIN2(n1192), 
        .Q(\IDinst/n7537 ) );
  nnd2s1 \IDinst/U7567  ( .DIN1(\IDinst/n7526 ), .DIN2(n1185), 
        .Q(\IDinst/n7536 ) );
  nnd2s1 \IDinst/U7566  ( .DIN1(\IDinst/n7534 ), .DIN2(\IDinst/n7533 ), 
        .Q(\IDinst/n7535 ) );
  nnd2s1 \IDinst/U7565  ( .DIN1(\IDinst/n7532 ), .DIN2(n1155), 
        .Q(\IDinst/n7534 ) );
  nnd2s1 \IDinst/U7564  ( .DIN1(\IDinst/n7529 ), .DIN2(n1152), 
        .Q(\IDinst/n7533 ) );
  nnd2s1 \IDinst/U7563  ( .DIN1(\IDinst/n7531 ), .DIN2(\IDinst/n7530 ), 
        .Q(\IDinst/n7532 ) );
  nnd2s1 \IDinst/U7562  ( .DIN1(\IDinst/RegFile[31][16] ), .DIN2(n1077), 
        .Q(\IDinst/n7531 ) );
  nnd2s1 \IDinst/U7561  ( .DIN1(\IDinst/RegFile[30][16] ), .DIN2(n1056), 
        .Q(\IDinst/n7530 ) );
  nnd2s1 \IDinst/U7560  ( .DIN1(\IDinst/n7528 ), .DIN2(\IDinst/n7527 ), 
        .Q(\IDinst/n7529 ) );
  nnd2s1 \IDinst/U7559  ( .DIN1(\IDinst/RegFile[29][16] ), .DIN2(n1077), 
        .Q(\IDinst/n7528 ) );
  nnd2s1 \IDinst/U7558  ( .DIN1(\IDinst/RegFile[28][16] ), .DIN2(n1056), 
        .Q(\IDinst/n7527 ) );
  nnd2s1 \IDinst/U7557  ( .DIN1(\IDinst/n7525 ), .DIN2(\IDinst/n7524 ), 
        .Q(\IDinst/n7526 ) );
  nnd2s1 \IDinst/U7556  ( .DIN1(\IDinst/n7523 ), .DIN2(n1154), 
        .Q(\IDinst/n7525 ) );
  nnd2s1 \IDinst/U7555  ( .DIN1(\IDinst/n7520 ), .DIN2(n1152), 
        .Q(\IDinst/n7524 ) );
  nnd2s1 \IDinst/U7554  ( .DIN1(\IDinst/n7522 ), .DIN2(\IDinst/n7521 ), 
        .Q(\IDinst/n7523 ) );
  nnd2s1 \IDinst/U7553  ( .DIN1(\IDinst/RegFile[27][16] ), .DIN2(n1077), 
        .Q(\IDinst/n7522 ) );
  nnd2s1 \IDinst/U7552  ( .DIN1(\IDinst/RegFile[26][16] ), .DIN2(n1056), 
        .Q(\IDinst/n7521 ) );
  nnd2s1 \IDinst/U7551  ( .DIN1(\IDinst/n7519 ), .DIN2(\IDinst/n7518 ), 
        .Q(\IDinst/n7520 ) );
  nnd2s1 \IDinst/U7550  ( .DIN1(\IDinst/RegFile[25][16] ), .DIN2(n1077), 
        .Q(\IDinst/n7519 ) );
  nnd2s1 \IDinst/U7549  ( .DIN1(\IDinst/RegFile[24][16] ), .DIN2(n1056), 
        .Q(\IDinst/n7518 ) );
  nnd2s1 \IDinst/U7548  ( .DIN1(\IDinst/n7516 ), .DIN2(\IDinst/n7515 ), 
        .Q(\IDinst/n7517 ) );
  nnd2s1 \IDinst/U7547  ( .DIN1(\IDinst/n7514 ), .DIN2(n1192), 
        .Q(\IDinst/n7516 ) );
  nnd2s1 \IDinst/U7546  ( .DIN1(\IDinst/n7505 ), .DIN2(n1185), 
        .Q(\IDinst/n7515 ) );
  nnd2s1 \IDinst/U7545  ( .DIN1(\IDinst/n7513 ), .DIN2(\IDinst/n7512 ), 
        .Q(\IDinst/n7514 ) );
  nnd2s1 \IDinst/U7544  ( .DIN1(\IDinst/n7511 ), .DIN2(n1154), 
        .Q(\IDinst/n7513 ) );
  nnd2s1 \IDinst/U7543  ( .DIN1(\IDinst/n7508 ), .DIN2(n1152), 
        .Q(\IDinst/n7512 ) );
  nnd2s1 \IDinst/U7542  ( .DIN1(\IDinst/n7510 ), .DIN2(\IDinst/n7509 ), 
        .Q(\IDinst/n7511 ) );
  nnd2s1 \IDinst/U7541  ( .DIN1(\IDinst/RegFile[23][16] ), .DIN2(n1077), 
        .Q(\IDinst/n7510 ) );
  nnd2s1 \IDinst/U7540  ( .DIN1(\IDinst/RegFile[22][16] ), .DIN2(n1056), 
        .Q(\IDinst/n7509 ) );
  nnd2s1 \IDinst/U7539  ( .DIN1(\IDinst/n7507 ), .DIN2(\IDinst/n7506 ), 
        .Q(\IDinst/n7508 ) );
  nnd2s1 \IDinst/U7538  ( .DIN1(\IDinst/RegFile[21][16] ), .DIN2(n1077), 
        .Q(\IDinst/n7507 ) );
  nnd2s1 \IDinst/U7537  ( .DIN1(\IDinst/RegFile[20][16] ), .DIN2(n1055), 
        .Q(\IDinst/n7506 ) );
  nnd2s1 \IDinst/U7536  ( .DIN1(\IDinst/n7504 ), .DIN2(\IDinst/n7503 ), 
        .Q(\IDinst/n7505 ) );
  nnd2s1 \IDinst/U7535  ( .DIN1(\IDinst/n7502 ), .DIN2(n1154), 
        .Q(\IDinst/n7504 ) );
  nnd2s1 \IDinst/U7534  ( .DIN1(\IDinst/n7499 ), .DIN2(n1180), 
        .Q(\IDinst/n7503 ) );
  nnd2s1 \IDinst/U7533  ( .DIN1(\IDinst/n7501 ), .DIN2(\IDinst/n7500 ), 
        .Q(\IDinst/n7502 ) );
  nnd2s1 \IDinst/U7532  ( .DIN1(\IDinst/RegFile[19][16] ), .DIN2(n1077), 
        .Q(\IDinst/n7501 ) );
  nnd2s1 \IDinst/U7531  ( .DIN1(\IDinst/RegFile[18][16] ), .DIN2(n1055), 
        .Q(\IDinst/n7500 ) );
  nnd2s1 \IDinst/U7530  ( .DIN1(\IDinst/n7498 ), .DIN2(\IDinst/n7497 ), 
        .Q(\IDinst/n7499 ) );
  nnd2s1 \IDinst/U7529  ( .DIN1(\IDinst/RegFile[17][16] ), .DIN2(n1077), 
        .Q(\IDinst/n7498 ) );
  nnd2s1 \IDinst/U7528  ( .DIN1(\IDinst/RegFile[16][16] ), .DIN2(n1055), 
        .Q(\IDinst/n7497 ) );
  nnd2s1 \IDinst/U7527  ( .DIN1(\IDinst/n7495 ), .DIN2(\IDinst/n7494 ), 
        .Q(\IDinst/n7496 ) );
  nnd2s1 \IDinst/U7526  ( .DIN1(\IDinst/n7493 ), .DIN2(n644), 
        .Q(\IDinst/n7495 ) );
  nnd2s1 \IDinst/U7525  ( .DIN1(\IDinst/n7472 ), .DIN2(n672), 
        .Q(\IDinst/n7494 ) );
  nnd2s1 \IDinst/U7524  ( .DIN1(\IDinst/n7492 ), .DIN2(\IDinst/n7491 ), 
        .Q(\IDinst/n7493 ) );
  nnd2s1 \IDinst/U7523  ( .DIN1(\IDinst/n7490 ), .DIN2(n1192), 
        .Q(\IDinst/n7492 ) );
  nnd2s1 \IDinst/U7522  ( .DIN1(\IDinst/n7481 ), .DIN2(n1185), 
        .Q(\IDinst/n7491 ) );
  nnd2s1 \IDinst/U7521  ( .DIN1(\IDinst/n7489 ), .DIN2(\IDinst/n7488 ), 
        .Q(\IDinst/n7490 ) );
  nnd2s1 \IDinst/U7520  ( .DIN1(\IDinst/n7487 ), .DIN2(n1154), 
        .Q(\IDinst/n7489 ) );
  nnd2s1 \IDinst/U7519  ( .DIN1(\IDinst/n7484 ), .DIN2(n1151), 
        .Q(\IDinst/n7488 ) );
  nnd2s1 \IDinst/U7518  ( .DIN1(\IDinst/n7486 ), .DIN2(\IDinst/n7485 ), 
        .Q(\IDinst/n7487 ) );
  nnd2s1 \IDinst/U7517  ( .DIN1(\IDinst/RegFile[15][16] ), .DIN2(n1078), 
        .Q(\IDinst/n7486 ) );
  nnd2s1 \IDinst/U7516  ( .DIN1(\IDinst/RegFile[14][16] ), .DIN2(n1055), 
        .Q(\IDinst/n7485 ) );
  nnd2s1 \IDinst/U7515  ( .DIN1(\IDinst/n7483 ), .DIN2(\IDinst/n7482 ), 
        .Q(\IDinst/n7484 ) );
  nnd2s1 \IDinst/U7514  ( .DIN1(\IDinst/RegFile[13][16] ), .DIN2(n1078), 
        .Q(\IDinst/n7483 ) );
  nnd2s1 \IDinst/U7513  ( .DIN1(\IDinst/RegFile[12][16] ), .DIN2(n1055), 
        .Q(\IDinst/n7482 ) );
  nnd2s1 \IDinst/U7512  ( .DIN1(\IDinst/n7480 ), .DIN2(\IDinst/n7479 ), 
        .Q(\IDinst/n7481 ) );
  nnd2s1 \IDinst/U7511  ( .DIN1(\IDinst/n7478 ), .DIN2(n1154), 
        .Q(\IDinst/n7480 ) );
  nnd2s1 \IDinst/U7510  ( .DIN1(\IDinst/n7475 ), .DIN2(n1133), 
        .Q(\IDinst/n7479 ) );
  nnd2s1 \IDinst/U7509  ( .DIN1(\IDinst/n7477 ), .DIN2(\IDinst/n7476 ), 
        .Q(\IDinst/n7478 ) );
  nnd2s1 \IDinst/U7508  ( .DIN1(\IDinst/RegFile[11][16] ), .DIN2(n1078), 
        .Q(\IDinst/n7477 ) );
  nnd2s1 \IDinst/U7507  ( .DIN1(\IDinst/RegFile[10][16] ), .DIN2(n1055), 
        .Q(\IDinst/n7476 ) );
  nnd2s1 \IDinst/U7506  ( .DIN1(\IDinst/n7474 ), .DIN2(\IDinst/n7473 ), 
        .Q(\IDinst/n7475 ) );
  nnd2s1 \IDinst/U7505  ( .DIN1(\IDinst/RegFile[9][16] ), .DIN2(n1078), 
        .Q(\IDinst/n7474 ) );
  nnd2s1 \IDinst/U7504  ( .DIN1(\IDinst/RegFile[8][16] ), .DIN2(n1055), 
        .Q(\IDinst/n7473 ) );
  nnd2s1 \IDinst/U7503  ( .DIN1(\IDinst/n7471 ), .DIN2(\IDinst/n7470 ), 
        .Q(\IDinst/n7472 ) );
  nnd2s1 \IDinst/U7502  ( .DIN1(\IDinst/n7469 ), .DIN2(n1192), 
        .Q(\IDinst/n7471 ) );
  nnd2s1 \IDinst/U7501  ( .DIN1(\IDinst/n7460 ), .DIN2(n1185), 
        .Q(\IDinst/n7470 ) );
  nnd2s1 \IDinst/U7500  ( .DIN1(\IDinst/n7468 ), .DIN2(\IDinst/n7467 ), 
        .Q(\IDinst/n7469 ) );
  nnd2s1 \IDinst/U7499  ( .DIN1(\IDinst/n7466 ), .DIN2(n1154), 
        .Q(\IDinst/n7468 ) );
  nnd2s1 \IDinst/U7498  ( .DIN1(\IDinst/n7463 ), .DIN2(n1180), 
        .Q(\IDinst/n7467 ) );
  nnd2s1 \IDinst/U7497  ( .DIN1(\IDinst/n7465 ), .DIN2(\IDinst/n7464 ), 
        .Q(\IDinst/n7466 ) );
  nnd2s1 \IDinst/U7496  ( .DIN1(\IDinst/RegFile[7][16] ), .DIN2(n1078), 
        .Q(\IDinst/n7465 ) );
  nnd2s1 \IDinst/U7495  ( .DIN1(\IDinst/RegFile[6][16] ), .DIN2(n1055), 
        .Q(\IDinst/n7464 ) );
  nnd2s1 \IDinst/U7494  ( .DIN1(\IDinst/n7462 ), .DIN2(\IDinst/n7461 ), 
        .Q(\IDinst/n7463 ) );
  nnd2s1 \IDinst/U7493  ( .DIN1(\IDinst/RegFile[5][16] ), .DIN2(n1078), 
        .Q(\IDinst/n7462 ) );
  nnd2s1 \IDinst/U7492  ( .DIN1(\IDinst/RegFile[4][16] ), .DIN2(n1055), 
        .Q(\IDinst/n7461 ) );
  nnd2s1 \IDinst/U7491  ( .DIN1(\IDinst/n7459 ), .DIN2(\IDinst/n7458 ), 
        .Q(\IDinst/n7460 ) );
  nnd2s1 \IDinst/U7490  ( .DIN1(\IDinst/n7457 ), .DIN2(n1154), 
        .Q(\IDinst/n7459 ) );
  nnd2s1 \IDinst/U7489  ( .DIN1(\IDinst/n7454 ), .DIN2(n1138), 
        .Q(\IDinst/n7458 ) );
  nnd2s1 \IDinst/U7488  ( .DIN1(\IDinst/n7456 ), .DIN2(\IDinst/n7455 ), 
        .Q(\IDinst/n7457 ) );
  nnd2s1 \IDinst/U7487  ( .DIN1(\IDinst/RegFile[3][16] ), .DIN2(n1078), 
        .Q(\IDinst/n7456 ) );
  nnd2s1 \IDinst/U7486  ( .DIN1(\IDinst/RegFile[2][16] ), .DIN2(n1060), 
        .Q(\IDinst/n7455 ) );
  nnd2s1 \IDinst/U7485  ( .DIN1(\IDinst/n7453 ), .DIN2(\IDinst/n7452 ), 
        .Q(\IDinst/n7454 ) );
  nnd2s1 \IDinst/U7484  ( .DIN1(\IDinst/RegFile[1][16] ), .DIN2(n1078), 
        .Q(\IDinst/n7453 ) );
  nnd2s1 \IDinst/U7483  ( .DIN1(\IDinst/RegFile[0][16] ), .DIN2(n1035), 
        .Q(\IDinst/n7452 ) );
  nnd2s1 \IDinst/U7482  ( .DIN1(\IDinst/n7451 ), .DIN2(n539), 
        .Q(\IDinst/n5978 ) );
  nnd2s1 \IDinst/U7481  ( .DIN1(\IDinst/n7406 ), .DIN2(n635), 
        .Q(\IDinst/n5979 ) );
  nnd2s1 \IDinst/U7480  ( .DIN1(\IDinst/n7450 ), .DIN2(\IDinst/n7449 ), 
        .Q(\IDinst/n7451 ) );
  nnd2s1 \IDinst/U7479  ( .DIN1(\IDinst/n7448 ), .DIN2(n643), 
        .Q(\IDinst/n7450 ) );
  nnd2s1 \IDinst/U7478  ( .DIN1(\IDinst/n7427 ), .DIN2(n670), 
        .Q(\IDinst/n7449 ) );
  nnd2s1 \IDinst/U7477  ( .DIN1(\IDinst/n7447 ), .DIN2(\IDinst/n7446 ), 
        .Q(\IDinst/n7448 ) );
  nnd2s1 \IDinst/U7476  ( .DIN1(\IDinst/n7445 ), .DIN2(n1192), 
        .Q(\IDinst/n7447 ) );
  nnd2s1 \IDinst/U7475  ( .DIN1(\IDinst/n7436 ), .DIN2(n1185), 
        .Q(\IDinst/n7446 ) );
  nnd2s1 \IDinst/U7474  ( .DIN1(\IDinst/n7444 ), .DIN2(\IDinst/n7443 ), 
        .Q(\IDinst/n7445 ) );
  nnd2s1 \IDinst/U7473  ( .DIN1(\IDinst/n7442 ), .DIN2(n1154), 
        .Q(\IDinst/n7444 ) );
  nnd2s1 \IDinst/U7472  ( .DIN1(\IDinst/n7439 ), .DIN2(n1133), 
        .Q(\IDinst/n7443 ) );
  nnd2s1 \IDinst/U7471  ( .DIN1(\IDinst/n7441 ), .DIN2(\IDinst/n7440 ), 
        .Q(\IDinst/n7442 ) );
  nnd2s1 \IDinst/U7470  ( .DIN1(\IDinst/RegFile[31][15] ), .DIN2(n1078), 
        .Q(\IDinst/n7441 ) );
  nnd2s1 \IDinst/U7469  ( .DIN1(\IDinst/RegFile[30][15] ), .DIN2(n1035), 
        .Q(\IDinst/n7440 ) );
  nnd2s1 \IDinst/U7468  ( .DIN1(\IDinst/n7438 ), .DIN2(\IDinst/n7437 ), 
        .Q(\IDinst/n7439 ) );
  nnd2s1 \IDinst/U7467  ( .DIN1(\IDinst/RegFile[29][15] ), .DIN2(n1079), 
        .Q(\IDinst/n7438 ) );
  nnd2s1 \IDinst/U7466  ( .DIN1(\IDinst/RegFile[28][15] ), .DIN2(n1035), 
        .Q(\IDinst/n7437 ) );
  nnd2s1 \IDinst/U7465  ( .DIN1(\IDinst/n7435 ), .DIN2(\IDinst/n7434 ), 
        .Q(\IDinst/n7436 ) );
  nnd2s1 \IDinst/U7464  ( .DIN1(\IDinst/n7433 ), .DIN2(n1168), 
        .Q(\IDinst/n7435 ) );
  nnd2s1 \IDinst/U7463  ( .DIN1(\IDinst/n7430 ), .DIN2(n1133), 
        .Q(\IDinst/n7434 ) );
  nnd2s1 \IDinst/U7462  ( .DIN1(\IDinst/n7432 ), .DIN2(\IDinst/n7431 ), 
        .Q(\IDinst/n7433 ) );
  nnd2s1 \IDinst/U7461  ( .DIN1(\IDinst/RegFile[27][15] ), .DIN2(n1079), 
        .Q(\IDinst/n7432 ) );
  nnd2s1 \IDinst/U7460  ( .DIN1(\IDinst/RegFile[26][15] ), .DIN2(n1035), 
        .Q(\IDinst/n7431 ) );
  nnd2s1 \IDinst/U7459  ( .DIN1(\IDinst/n7429 ), .DIN2(\IDinst/n7428 ), 
        .Q(\IDinst/n7430 ) );
  nnd2s1 \IDinst/U7458  ( .DIN1(\IDinst/RegFile[25][15] ), .DIN2(n1079), 
        .Q(\IDinst/n7429 ) );
  nnd2s1 \IDinst/U7457  ( .DIN1(\IDinst/RegFile[24][15] ), .DIN2(n1035), 
        .Q(\IDinst/n7428 ) );
  nnd2s1 \IDinst/U7456  ( .DIN1(\IDinst/n7426 ), .DIN2(\IDinst/n7425 ), 
        .Q(\IDinst/n7427 ) );
  nnd2s1 \IDinst/U7455  ( .DIN1(\IDinst/n7424 ), .DIN2(n1191), 
        .Q(\IDinst/n7426 ) );
  nnd2s1 \IDinst/U7454  ( .DIN1(\IDinst/n7415 ), .DIN2(n1185), 
        .Q(\IDinst/n7425 ) );
  nnd2s1 \IDinst/U7453  ( .DIN1(\IDinst/n7423 ), .DIN2(\IDinst/n7422 ), 
        .Q(\IDinst/n7424 ) );
  nnd2s1 \IDinst/U7452  ( .DIN1(\IDinst/n7421 ), .DIN2(\IDinst/N40 ), 
        .Q(\IDinst/n7423 ) );
  nnd2s1 \IDinst/U7451  ( .DIN1(\IDinst/n7418 ), .DIN2(n1133), 
        .Q(\IDinst/n7422 ) );
  nnd2s1 \IDinst/U7450  ( .DIN1(\IDinst/n7420 ), .DIN2(\IDinst/n7419 ), 
        .Q(\IDinst/n7421 ) );
  nnd2s1 \IDinst/U7449  ( .DIN1(\IDinst/RegFile[23][15] ), .DIN2(n1079), 
        .Q(\IDinst/n7420 ) );
  nnd2s1 \IDinst/U7448  ( .DIN1(\IDinst/RegFile[22][15] ), .DIN2(n1035), 
        .Q(\IDinst/n7419 ) );
  nnd2s1 \IDinst/U7447  ( .DIN1(\IDinst/n7417 ), .DIN2(\IDinst/n7416 ), 
        .Q(\IDinst/n7418 ) );
  nnd2s1 \IDinst/U7446  ( .DIN1(\IDinst/RegFile[21][15] ), .DIN2(n1079), 
        .Q(\IDinst/n7417 ) );
  nnd2s1 \IDinst/U7445  ( .DIN1(\IDinst/RegFile[20][15] ), .DIN2(n1035), 
        .Q(\IDinst/n7416 ) );
  nnd2s1 \IDinst/U7444  ( .DIN1(\IDinst/n7414 ), .DIN2(\IDinst/n7413 ), 
        .Q(\IDinst/n7415 ) );
  nnd2s1 \IDinst/U7443  ( .DIN1(\IDinst/n7412 ), .DIN2(n1173), 
        .Q(\IDinst/n7414 ) );
  nnd2s1 \IDinst/U7442  ( .DIN1(\IDinst/n7409 ), .DIN2(n1134), 
        .Q(\IDinst/n7413 ) );
  nnd2s1 \IDinst/U7441  ( .DIN1(\IDinst/n7411 ), .DIN2(\IDinst/n7410 ), 
        .Q(\IDinst/n7412 ) );
  nnd2s1 \IDinst/U7440  ( .DIN1(\IDinst/RegFile[19][15] ), .DIN2(n1079), 
        .Q(\IDinst/n7411 ) );
  nnd2s1 \IDinst/U7439  ( .DIN1(\IDinst/RegFile[18][15] ), .DIN2(n1035), 
        .Q(\IDinst/n7410 ) );
  nnd2s1 \IDinst/U7438  ( .DIN1(\IDinst/n7408 ), .DIN2(\IDinst/n7407 ), 
        .Q(\IDinst/n7409 ) );
  nnd2s1 \IDinst/U7437  ( .DIN1(\IDinst/RegFile[17][15] ), .DIN2(n1079), 
        .Q(\IDinst/n7408 ) );
  nnd2s1 \IDinst/U7436  ( .DIN1(\IDinst/RegFile[16][15] ), .DIN2(n1034), 
        .Q(\IDinst/n7407 ) );
  nnd2s1 \IDinst/U7435  ( .DIN1(\IDinst/n7405 ), .DIN2(\IDinst/n7404 ), 
        .Q(\IDinst/n7406 ) );
  nnd2s1 \IDinst/U7434  ( .DIN1(\IDinst/n7403 ), .DIN2(n642), 
        .Q(\IDinst/n7405 ) );
  nnd2s1 \IDinst/U7433  ( .DIN1(\IDinst/n7382 ), .DIN2(n673), 
        .Q(\IDinst/n7404 ) );
  nnd2s1 \IDinst/U7432  ( .DIN1(\IDinst/n7402 ), .DIN2(\IDinst/n7401 ), 
        .Q(\IDinst/n7403 ) );
  nnd2s1 \IDinst/U7431  ( .DIN1(\IDinst/n7400 ), .DIN2(n1197), 
        .Q(\IDinst/n7402 ) );
  nnd2s1 \IDinst/U7430  ( .DIN1(\IDinst/n7391 ), .DIN2(n1185), 
        .Q(\IDinst/n7401 ) );
  nnd2s1 \IDinst/U7429  ( .DIN1(\IDinst/n7399 ), .DIN2(\IDinst/n7398 ), 
        .Q(\IDinst/n7400 ) );
  nnd2s1 \IDinst/U7428  ( .DIN1(\IDinst/n7397 ), .DIN2(n1163), 
        .Q(\IDinst/n7399 ) );
  nnd2s1 \IDinst/U7427  ( .DIN1(\IDinst/n7394 ), .DIN2(n1134), 
        .Q(\IDinst/n7398 ) );
  nnd2s1 \IDinst/U7426  ( .DIN1(\IDinst/n7396 ), .DIN2(\IDinst/n7395 ), 
        .Q(\IDinst/n7397 ) );
  nnd2s1 \IDinst/U7425  ( .DIN1(\IDinst/RegFile[15][15] ), .DIN2(n1079), 
        .Q(\IDinst/n7396 ) );
  nnd2s1 \IDinst/U7424  ( .DIN1(\IDinst/RegFile[14][15] ), .DIN2(n1034), 
        .Q(\IDinst/n7395 ) );
  nnd2s1 \IDinst/U7423  ( .DIN1(\IDinst/n7393 ), .DIN2(\IDinst/n7392 ), 
        .Q(\IDinst/n7394 ) );
  nnd2s1 \IDinst/U7422  ( .DIN1(\IDinst/RegFile[13][15] ), .DIN2(n1079), 
        .Q(\IDinst/n7393 ) );
  nnd2s1 \IDinst/U7421  ( .DIN1(\IDinst/RegFile[12][15] ), .DIN2(n1034), 
        .Q(\IDinst/n7392 ) );
  nnd2s1 \IDinst/U7420  ( .DIN1(\IDinst/n7390 ), .DIN2(\IDinst/n7389 ), 
        .Q(\IDinst/n7391 ) );
  nnd2s1 \IDinst/U7419  ( .DIN1(\IDinst/n7388 ), .DIN2(n1164), 
        .Q(\IDinst/n7390 ) );
  nnd2s1 \IDinst/U7418  ( .DIN1(\IDinst/n7385 ), .DIN2(n1134), 
        .Q(\IDinst/n7389 ) );
  nnd2s1 \IDinst/U7417  ( .DIN1(\IDinst/n7387 ), .DIN2(\IDinst/n7386 ), 
        .Q(\IDinst/n7388 ) );
  nnd2s1 \IDinst/U7416  ( .DIN1(\IDinst/RegFile[11][15] ), .DIN2(n1080), 
        .Q(\IDinst/n7387 ) );
  nnd2s1 \IDinst/U7415  ( .DIN1(\IDinst/RegFile[10][15] ), .DIN2(n1034), 
        .Q(\IDinst/n7386 ) );
  nnd2s1 \IDinst/U7414  ( .DIN1(\IDinst/n7384 ), .DIN2(\IDinst/n7383 ), 
        .Q(\IDinst/n7385 ) );
  nnd2s1 \IDinst/U7413  ( .DIN1(\IDinst/RegFile[9][15] ), .DIN2(n1080), 
        .Q(\IDinst/n7384 ) );
  nnd2s1 \IDinst/U7412  ( .DIN1(\IDinst/RegFile[8][15] ), .DIN2(n1034), 
        .Q(\IDinst/n7383 ) );
  nnd2s1 \IDinst/U7411  ( .DIN1(\IDinst/n7381 ), .DIN2(\IDinst/n7380 ), 
        .Q(\IDinst/n7382 ) );
  nnd2s1 \IDinst/U7410  ( .DIN1(\IDinst/n7379 ), .DIN2(n1196), 
        .Q(\IDinst/n7381 ) );
  nnd2s1 \IDinst/U7409  ( .DIN1(\IDinst/n7370 ), .DIN2(n1185), 
        .Q(\IDinst/n7380 ) );
  nnd2s1 \IDinst/U7408  ( .DIN1(\IDinst/n7378 ), .DIN2(\IDinst/n7377 ), 
        .Q(\IDinst/n7379 ) );
  nnd2s1 \IDinst/U7407  ( .DIN1(\IDinst/n7376 ), .DIN2(n1159), 
        .Q(\IDinst/n7378 ) );
  nnd2s1 \IDinst/U7406  ( .DIN1(\IDinst/n7373 ), .DIN2(n1134), 
        .Q(\IDinst/n7377 ) );
  nnd2s1 \IDinst/U7405  ( .DIN1(\IDinst/n7375 ), .DIN2(\IDinst/n7374 ), 
        .Q(\IDinst/n7376 ) );
  nnd2s1 \IDinst/U7404  ( .DIN1(\IDinst/RegFile[7][15] ), .DIN2(n1080), 
        .Q(\IDinst/n7375 ) );
  nnd2s1 \IDinst/U7403  ( .DIN1(\IDinst/RegFile[6][15] ), .DIN2(n1034), 
        .Q(\IDinst/n7374 ) );
  nnd2s1 \IDinst/U7402  ( .DIN1(\IDinst/n7372 ), .DIN2(\IDinst/n7371 ), 
        .Q(\IDinst/n7373 ) );
  nnd2s1 \IDinst/U7401  ( .DIN1(\IDinst/RegFile[5][15] ), .DIN2(n1080), 
        .Q(\IDinst/n7372 ) );
  nnd2s1 \IDinst/U7400  ( .DIN1(\IDinst/RegFile[4][15] ), .DIN2(n1034), 
        .Q(\IDinst/n7371 ) );
  nnd2s1 \IDinst/U7399  ( .DIN1(\IDinst/n7369 ), .DIN2(\IDinst/n7368 ), 
        .Q(\IDinst/n7370 ) );
  nnd2s1 \IDinst/U7398  ( .DIN1(\IDinst/n7367 ), .DIN2(n1175), 
        .Q(\IDinst/n7369 ) );
  nnd2s1 \IDinst/U7397  ( .DIN1(\IDinst/n7364 ), .DIN2(n1134), 
        .Q(\IDinst/n7368 ) );
  nnd2s1 \IDinst/U7396  ( .DIN1(\IDinst/n7366 ), .DIN2(\IDinst/n7365 ), 
        .Q(\IDinst/n7367 ) );
  nnd2s1 \IDinst/U7395  ( .DIN1(\IDinst/RegFile[3][15] ), .DIN2(n1080), 
        .Q(\IDinst/n7366 ) );
  nnd2s1 \IDinst/U7394  ( .DIN1(\IDinst/RegFile[2][15] ), .DIN2(n1034), 
        .Q(\IDinst/n7365 ) );
  nnd2s1 \IDinst/U7393  ( .DIN1(\IDinst/n7363 ), .DIN2(\IDinst/n7362 ), 
        .Q(\IDinst/n7364 ) );
  nnd2s1 \IDinst/U7392  ( .DIN1(\IDinst/RegFile[1][15] ), .DIN2(n1080), 
        .Q(\IDinst/n7363 ) );
  nnd2s1 \IDinst/U7391  ( .DIN1(\IDinst/RegFile[0][15] ), .DIN2(n1034), 
        .Q(\IDinst/n7362 ) );
  nnd2s1 \IDinst/U7390  ( .DIN1(\IDinst/n7361 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n5976 ) );
  nnd2s1 \IDinst/U7389  ( .DIN1(\IDinst/n7316 ), .DIN2(n636), 
        .Q(\IDinst/n5977 ) );
  nnd2s1 \IDinst/U7388  ( .DIN1(\IDinst/n7360 ), .DIN2(\IDinst/n7359 ), 
        .Q(\IDinst/n7361 ) );
  nnd2s1 \IDinst/U7387  ( .DIN1(\IDinst/n7358 ), .DIN2(n641), 
        .Q(\IDinst/n7360 ) );
  nnd2s1 \IDinst/U7386  ( .DIN1(\IDinst/n7337 ), .DIN2(n671), 
        .Q(\IDinst/n7359 ) );
  nnd2s1 \IDinst/U7385  ( .DIN1(\IDinst/n7357 ), .DIN2(\IDinst/n7356 ), 
        .Q(\IDinst/n7358 ) );
  nnd2s1 \IDinst/U7384  ( .DIN1(\IDinst/n7355 ), .DIN2(n1196), 
        .Q(\IDinst/n7357 ) );
  nnd2s1 \IDinst/U7383  ( .DIN1(\IDinst/n7346 ), .DIN2(n1185), 
        .Q(\IDinst/n7356 ) );
  nnd2s1 \IDinst/U7382  ( .DIN1(\IDinst/n7354 ), .DIN2(\IDinst/n7353 ), 
        .Q(\IDinst/n7355 ) );
  nnd2s1 \IDinst/U7381  ( .DIN1(\IDinst/n7352 ), .DIN2(n1166), 
        .Q(\IDinst/n7354 ) );
  nnd2s1 \IDinst/U7380  ( .DIN1(\IDinst/n7349 ), .DIN2(n1134), 
        .Q(\IDinst/n7353 ) );
  nnd2s1 \IDinst/U7379  ( .DIN1(\IDinst/n7351 ), .DIN2(\IDinst/n7350 ), 
        .Q(\IDinst/n7352 ) );
  nnd2s1 \IDinst/U7378  ( .DIN1(\IDinst/RegFile[31][14] ), .DIN2(n1080), 
        .Q(\IDinst/n7351 ) );
  nnd2s1 \IDinst/U7377  ( .DIN1(\IDinst/RegFile[30][14] ), .DIN2(n1034), 
        .Q(\IDinst/n7350 ) );
  nnd2s1 \IDinst/U7376  ( .DIN1(\IDinst/n7348 ), .DIN2(\IDinst/n7347 ), 
        .Q(\IDinst/n7349 ) );
  nnd2s1 \IDinst/U7375  ( .DIN1(\IDinst/RegFile[29][14] ), .DIN2(n1080), 
        .Q(\IDinst/n7348 ) );
  nnd2s1 \IDinst/U7374  ( .DIN1(\IDinst/RegFile[28][14] ), .DIN2(n1034), 
        .Q(\IDinst/n7347 ) );
  nnd2s1 \IDinst/U7373  ( .DIN1(\IDinst/n7345 ), .DIN2(\IDinst/n7344 ), 
        .Q(\IDinst/n7346 ) );
  nnd2s1 \IDinst/U7372  ( .DIN1(\IDinst/n7343 ), .DIN2(n1153), 
        .Q(\IDinst/n7345 ) );
  nnd2s1 \IDinst/U7371  ( .DIN1(\IDinst/n7340 ), .DIN2(n1134), 
        .Q(\IDinst/n7344 ) );
  nnd2s1 \IDinst/U7370  ( .DIN1(\IDinst/n7342 ), .DIN2(\IDinst/n7341 ), 
        .Q(\IDinst/n7343 ) );
  nnd2s1 \IDinst/U7369  ( .DIN1(\IDinst/RegFile[27][14] ), .DIN2(n1080), 
        .Q(\IDinst/n7342 ) );
  nnd2s1 \IDinst/U7368  ( .DIN1(\IDinst/RegFile[26][14] ), .DIN2(n1034), 
        .Q(\IDinst/n7341 ) );
  nnd2s1 \IDinst/U7367  ( .DIN1(\IDinst/n7339 ), .DIN2(\IDinst/n7338 ), 
        .Q(\IDinst/n7340 ) );
  nnd2s1 \IDinst/U7366  ( .DIN1(\IDinst/RegFile[25][14] ), .DIN2(n1081), 
        .Q(\IDinst/n7339 ) );
  nnd2s1 \IDinst/U7365  ( .DIN1(\IDinst/RegFile[24][14] ), .DIN2(n1034), 
        .Q(\IDinst/n7338 ) );
  nnd2s1 \IDinst/U7364  ( .DIN1(\IDinst/n7336 ), .DIN2(\IDinst/n7335 ), 
        .Q(\IDinst/n7337 ) );
  nnd2s1 \IDinst/U7363  ( .DIN1(\IDinst/n7334 ), .DIN2(n1195), 
        .Q(\IDinst/n7336 ) );
  nnd2s1 \IDinst/U7362  ( .DIN1(\IDinst/n7325 ), .DIN2(n1185), 
        .Q(\IDinst/n7335 ) );
  nnd2s1 \IDinst/U7361  ( .DIN1(\IDinst/n7333 ), .DIN2(\IDinst/n7332 ), 
        .Q(\IDinst/n7334 ) );
  nnd2s1 \IDinst/U7360  ( .DIN1(\IDinst/n7331 ), .DIN2(n1159), 
        .Q(\IDinst/n7333 ) );
  nnd2s1 \IDinst/U7359  ( .DIN1(\IDinst/n7328 ), .DIN2(n1134), 
        .Q(\IDinst/n7332 ) );
  nnd2s1 \IDinst/U7358  ( .DIN1(\IDinst/n7330 ), .DIN2(\IDinst/n7329 ), 
        .Q(\IDinst/n7331 ) );
  nnd2s1 \IDinst/U7357  ( .DIN1(\IDinst/RegFile[23][14] ), .DIN2(n1081), 
        .Q(\IDinst/n7330 ) );
  nnd2s1 \IDinst/U7356  ( .DIN1(\IDinst/RegFile[22][14] ), .DIN2(n1033), 
        .Q(\IDinst/n7329 ) );
  nnd2s1 \IDinst/U7355  ( .DIN1(\IDinst/n7327 ), .DIN2(\IDinst/n7326 ), 
        .Q(\IDinst/n7328 ) );
  nnd2s1 \IDinst/U7354  ( .DIN1(\IDinst/RegFile[21][14] ), .DIN2(n1109), 
        .Q(\IDinst/n7327 ) );
  nnd2s1 \IDinst/U7353  ( .DIN1(\IDinst/RegFile[20][14] ), .DIN2(n1033), 
        .Q(\IDinst/n7326 ) );
  nnd2s1 \IDinst/U7352  ( .DIN1(\IDinst/n7324 ), .DIN2(\IDinst/n7323 ), 
        .Q(\IDinst/n7325 ) );
  nnd2s1 \IDinst/U7351  ( .DIN1(\IDinst/n7322 ), .DIN2(n1178), 
        .Q(\IDinst/n7324 ) );
  nnd2s1 \IDinst/U7350  ( .DIN1(\IDinst/n7319 ), .DIN2(n1134), 
        .Q(\IDinst/n7323 ) );
  nnd2s1 \IDinst/U7349  ( .DIN1(\IDinst/n7321 ), .DIN2(\IDinst/n7320 ), 
        .Q(\IDinst/n7322 ) );
  nnd2s1 \IDinst/U7348  ( .DIN1(\IDinst/RegFile[19][14] ), .DIN2(n1109), 
        .Q(\IDinst/n7321 ) );
  nnd2s1 \IDinst/U7347  ( .DIN1(\IDinst/RegFile[18][14] ), .DIN2(n1033), 
        .Q(\IDinst/n7320 ) );
  nnd2s1 \IDinst/U7346  ( .DIN1(\IDinst/n7318 ), .DIN2(\IDinst/n7317 ), 
        .Q(\IDinst/n7319 ) );
  nnd2s1 \IDinst/U7345  ( .DIN1(\IDinst/RegFile[17][14] ), .DIN2(n1109), 
        .Q(\IDinst/n7318 ) );
  nnd2s1 \IDinst/U7344  ( .DIN1(\IDinst/RegFile[16][14] ), .DIN2(n1033), 
        .Q(\IDinst/n7317 ) );
  nnd2s1 \IDinst/U7343  ( .DIN1(\IDinst/n7315 ), .DIN2(\IDinst/n7314 ), 
        .Q(\IDinst/n7316 ) );
  nnd2s1 \IDinst/U7342  ( .DIN1(\IDinst/n7313 ), .DIN2(n644), 
        .Q(\IDinst/n7315 ) );
  nnd2s1 \IDinst/U7341  ( .DIN1(\IDinst/n7292 ), .DIN2(n672), 
        .Q(\IDinst/n7314 ) );
  nnd2s1 \IDinst/U7340  ( .DIN1(\IDinst/n7312 ), .DIN2(\IDinst/n7311 ), 
        .Q(\IDinst/n7313 ) );
  nnd2s1 \IDinst/U7339  ( .DIN1(\IDinst/n7310 ), .DIN2(n1190), 
        .Q(\IDinst/n7312 ) );
  nnd2s1 \IDinst/U7338  ( .DIN1(\IDinst/n7301 ), .DIN2(n1184), 
        .Q(\IDinst/n7311 ) );
  nnd2s1 \IDinst/U7337  ( .DIN1(\IDinst/n7309 ), .DIN2(\IDinst/n7308 ), 
        .Q(\IDinst/n7310 ) );
  nnd2s1 \IDinst/U7336  ( .DIN1(\IDinst/n7307 ), .DIN2(n1178), 
        .Q(\IDinst/n7309 ) );
  nnd2s1 \IDinst/U7335  ( .DIN1(\IDinst/n7304 ), .DIN2(n1134), 
        .Q(\IDinst/n7308 ) );
  nnd2s1 \IDinst/U7334  ( .DIN1(\IDinst/n7306 ), .DIN2(\IDinst/n7305 ), 
        .Q(\IDinst/n7307 ) );
  nnd2s1 \IDinst/U7333  ( .DIN1(\IDinst/RegFile[15][14] ), .DIN2(n1109), 
        .Q(\IDinst/n7306 ) );
  nnd2s1 \IDinst/U7332  ( .DIN1(\IDinst/RegFile[14][14] ), .DIN2(n1033), 
        .Q(\IDinst/n7305 ) );
  nnd2s1 \IDinst/U7331  ( .DIN1(\IDinst/n7303 ), .DIN2(\IDinst/n7302 ), 
        .Q(\IDinst/n7304 ) );
  nnd2s1 \IDinst/U7330  ( .DIN1(\IDinst/RegFile[13][14] ), .DIN2(n1110), 
        .Q(\IDinst/n7303 ) );
  nnd2s1 \IDinst/U7329  ( .DIN1(\IDinst/RegFile[12][14] ), .DIN2(n1033), 
        .Q(\IDinst/n7302 ) );
  nnd2s1 \IDinst/U7328  ( .DIN1(\IDinst/n7300 ), .DIN2(\IDinst/n7299 ), 
        .Q(\IDinst/n7301 ) );
  nnd2s1 \IDinst/U7327  ( .DIN1(\IDinst/n7298 ), .DIN2(n1177), 
        .Q(\IDinst/n7300 ) );
  nnd2s1 \IDinst/U7326  ( .DIN1(\IDinst/n7295 ), .DIN2(n1134), 
        .Q(\IDinst/n7299 ) );
  nnd2s1 \IDinst/U7325  ( .DIN1(\IDinst/n7297 ), .DIN2(\IDinst/n7296 ), 
        .Q(\IDinst/n7298 ) );
  nnd2s1 \IDinst/U7324  ( .DIN1(\IDinst/RegFile[11][14] ), .DIN2(n1110), 
        .Q(\IDinst/n7297 ) );
  nnd2s1 \IDinst/U7323  ( .DIN1(\IDinst/RegFile[10][14] ), .DIN2(n1033), 
        .Q(\IDinst/n7296 ) );
  nnd2s1 \IDinst/U7322  ( .DIN1(\IDinst/n7294 ), .DIN2(\IDinst/n7293 ), 
        .Q(\IDinst/n7295 ) );
  nnd2s1 \IDinst/U7321  ( .DIN1(\IDinst/RegFile[9][14] ), .DIN2(n1110), 
        .Q(\IDinst/n7294 ) );
  nnd2s1 \IDinst/U7320  ( .DIN1(\IDinst/RegFile[8][14] ), .DIN2(n1033), 
        .Q(\IDinst/n7293 ) );
  nnd2s1 \IDinst/U7319  ( .DIN1(\IDinst/n7291 ), .DIN2(\IDinst/n7290 ), 
        .Q(\IDinst/n7292 ) );
  nnd2s1 \IDinst/U7318  ( .DIN1(\IDinst/n7289 ), .DIN2(n1190), 
        .Q(\IDinst/n7291 ) );
  nnd2s1 \IDinst/U7317  ( .DIN1(\IDinst/n7280 ), .DIN2(n1184), 
        .Q(\IDinst/n7290 ) );
  nnd2s1 \IDinst/U7316  ( .DIN1(\IDinst/n7288 ), .DIN2(\IDinst/n7287 ), 
        .Q(\IDinst/n7289 ) );
  nnd2s1 \IDinst/U7315  ( .DIN1(\IDinst/n7286 ), .DIN2(n1177), 
        .Q(\IDinst/n7288 ) );
  nnd2s1 \IDinst/U7314  ( .DIN1(\IDinst/n7283 ), .DIN2(n1134), 
        .Q(\IDinst/n7287 ) );
  nnd2s1 \IDinst/U7313  ( .DIN1(\IDinst/n7285 ), .DIN2(\IDinst/n7284 ), 
        .Q(\IDinst/n7286 ) );
  nnd2s1 \IDinst/U7312  ( .DIN1(\IDinst/RegFile[7][14] ), .DIN2(n1110), 
        .Q(\IDinst/n7285 ) );
  nnd2s1 \IDinst/U7311  ( .DIN1(\IDinst/RegFile[6][14] ), .DIN2(n1033), 
        .Q(\IDinst/n7284 ) );
  nnd2s1 \IDinst/U7310  ( .DIN1(\IDinst/n7282 ), .DIN2(\IDinst/n7281 ), 
        .Q(\IDinst/n7283 ) );
  nnd2s1 \IDinst/U7309  ( .DIN1(\IDinst/RegFile[5][14] ), .DIN2(n1110), 
        .Q(\IDinst/n7282 ) );
  nnd2s1 \IDinst/U7308  ( .DIN1(\IDinst/RegFile[4][14] ), .DIN2(n1033), 
        .Q(\IDinst/n7281 ) );
  nnd2s1 \IDinst/U7307  ( .DIN1(\IDinst/n7279 ), .DIN2(\IDinst/n7278 ), 
        .Q(\IDinst/n7280 ) );
  nnd2s1 \IDinst/U7306  ( .DIN1(\IDinst/n7277 ), .DIN2(n1177), 
        .Q(\IDinst/n7279 ) );
  nnd2s1 \IDinst/U7305  ( .DIN1(\IDinst/n7274 ), .DIN2(n1134), 
        .Q(\IDinst/n7278 ) );
  nnd2s1 \IDinst/U7304  ( .DIN1(\IDinst/n7276 ), .DIN2(\IDinst/n7275 ), 
        .Q(\IDinst/n7277 ) );
  nnd2s1 \IDinst/U7303  ( .DIN1(\IDinst/RegFile[3][14] ), .DIN2(n1110), 
        .Q(\IDinst/n7276 ) );
  nnd2s1 \IDinst/U7302  ( .DIN1(\IDinst/RegFile[2][14] ), .DIN2(n1033), 
        .Q(\IDinst/n7275 ) );
  nnd2s1 \IDinst/U7301  ( .DIN1(\IDinst/n7273 ), .DIN2(\IDinst/n7272 ), 
        .Q(\IDinst/n7274 ) );
  nnd2s1 \IDinst/U7300  ( .DIN1(\IDinst/RegFile[1][14] ), .DIN2(n1110), 
        .Q(\IDinst/n7273 ) );
  nnd2s1 \IDinst/U7299  ( .DIN1(\IDinst/RegFile[0][14] ), .DIN2(n1033), 
        .Q(\IDinst/n7272 ) );
  nnd2s1 \IDinst/U7298  ( .DIN1(\IDinst/n7271 ), .DIN2(n539), 
        .Q(\IDinst/n5974 ) );
  nnd2s1 \IDinst/U7297  ( .DIN1(\IDinst/n7226 ), .DIN2(n635), 
        .Q(\IDinst/n5975 ) );
  nnd2s1 \IDinst/U7296  ( .DIN1(\IDinst/n7270 ), .DIN2(\IDinst/n7269 ), 
        .Q(\IDinst/n7271 ) );
  nnd2s1 \IDinst/U7295  ( .DIN1(\IDinst/n7268 ), .DIN2(n643), 
        .Q(\IDinst/n7270 ) );
  nnd2s1 \IDinst/U7294  ( .DIN1(\IDinst/n7247 ), .DIN2(n670), 
        .Q(\IDinst/n7269 ) );
  nnd2s1 \IDinst/U7293  ( .DIN1(\IDinst/n7267 ), .DIN2(\IDinst/n7266 ), 
        .Q(\IDinst/n7268 ) );
  nnd2s1 \IDinst/U7292  ( .DIN1(\IDinst/n7265 ), .DIN2(\IDinst/N41 ), 
        .Q(\IDinst/n7267 ) );
  nnd2s1 \IDinst/U7291  ( .DIN1(\IDinst/n7256 ), .DIN2(n1184), 
        .Q(\IDinst/n7266 ) );
  nnd2s1 \IDinst/U7290  ( .DIN1(\IDinst/n7264 ), .DIN2(\IDinst/n7263 ), 
        .Q(\IDinst/n7265 ) );
  nnd2s1 \IDinst/U7289  ( .DIN1(\IDinst/n7262 ), .DIN2(n1177), 
        .Q(\IDinst/n7264 ) );
  nnd2s1 \IDinst/U7288  ( .DIN1(\IDinst/n7259 ), .DIN2(n1135), 
        .Q(\IDinst/n7263 ) );
  nnd2s1 \IDinst/U7287  ( .DIN1(\IDinst/n7261 ), .DIN2(\IDinst/n7260 ), 
        .Q(\IDinst/n7262 ) );
  nnd2s1 \IDinst/U7286  ( .DIN1(\IDinst/RegFile[31][13] ), .DIN2(n1110), 
        .Q(\IDinst/n7261 ) );
  nnd2s1 \IDinst/U7285  ( .DIN1(\IDinst/RegFile[30][13] ), .DIN2(n1033), 
        .Q(\IDinst/n7260 ) );
  nnd2s1 \IDinst/U7284  ( .DIN1(\IDinst/n7258 ), .DIN2(\IDinst/n7257 ), 
        .Q(\IDinst/n7259 ) );
  nnd2s1 \IDinst/U7283  ( .DIN1(\IDinst/RegFile[29][13] ), .DIN2(n1110), 
        .Q(\IDinst/n7258 ) );
  nnd2s1 \IDinst/U7282  ( .DIN1(\IDinst/RegFile[28][13] ), .DIN2(n1032), 
        .Q(\IDinst/n7257 ) );
  nnd2s1 \IDinst/U7281  ( .DIN1(\IDinst/n7255 ), .DIN2(\IDinst/n7254 ), 
        .Q(\IDinst/n7256 ) );
  nnd2s1 \IDinst/U7280  ( .DIN1(\IDinst/n7253 ), .DIN2(n1177), 
        .Q(\IDinst/n7255 ) );
  nnd2s1 \IDinst/U7279  ( .DIN1(\IDinst/n7250 ), .DIN2(n1135), 
        .Q(\IDinst/n7254 ) );
  nnd2s1 \IDinst/U7278  ( .DIN1(\IDinst/n7252 ), .DIN2(\IDinst/n7251 ), 
        .Q(\IDinst/n7253 ) );
  nnd2s1 \IDinst/U7277  ( .DIN1(\IDinst/RegFile[27][13] ), .DIN2(n1111), 
        .Q(\IDinst/n7252 ) );
  nnd2s1 \IDinst/U7276  ( .DIN1(\IDinst/RegFile[26][13] ), .DIN2(n1032), 
        .Q(\IDinst/n7251 ) );
  nnd2s1 \IDinst/U7275  ( .DIN1(\IDinst/n7249 ), .DIN2(\IDinst/n7248 ), 
        .Q(\IDinst/n7250 ) );
  nnd2s1 \IDinst/U7274  ( .DIN1(\IDinst/RegFile[25][13] ), .DIN2(n1111), 
        .Q(\IDinst/n7249 ) );
  nnd2s1 \IDinst/U7273  ( .DIN1(\IDinst/RegFile[24][13] ), .DIN2(n1032), 
        .Q(\IDinst/n7248 ) );
  nnd2s1 \IDinst/U7272  ( .DIN1(\IDinst/n7246 ), .DIN2(\IDinst/n7245 ), 
        .Q(\IDinst/n7247 ) );
  nnd2s1 \IDinst/U7271  ( .DIN1(\IDinst/n7244 ), .DIN2(n1193), 
        .Q(\IDinst/n7246 ) );
  nnd2s1 \IDinst/U7270  ( .DIN1(\IDinst/n7235 ), .DIN2(n1184), 
        .Q(\IDinst/n7245 ) );
  nnd2s1 \IDinst/U7269  ( .DIN1(\IDinst/n7243 ), .DIN2(\IDinst/n7242 ), 
        .Q(\IDinst/n7244 ) );
  nnd2s1 \IDinst/U7268  ( .DIN1(\IDinst/n7241 ), .DIN2(n1177), 
        .Q(\IDinst/n7243 ) );
  nnd2s1 \IDinst/U7267  ( .DIN1(\IDinst/n7238 ), .DIN2(n1135), 
        .Q(\IDinst/n7242 ) );
  nnd2s1 \IDinst/U7266  ( .DIN1(\IDinst/n7240 ), .DIN2(\IDinst/n7239 ), 
        .Q(\IDinst/n7241 ) );
  nnd2s1 \IDinst/U7265  ( .DIN1(\IDinst/RegFile[23][13] ), .DIN2(n1111), 
        .Q(\IDinst/n7240 ) );
  nnd2s1 \IDinst/U7264  ( .DIN1(\IDinst/RegFile[22][13] ), .DIN2(n1032), 
        .Q(\IDinst/n7239 ) );
  nnd2s1 \IDinst/U7263  ( .DIN1(\IDinst/n7237 ), .DIN2(\IDinst/n7236 ), 
        .Q(\IDinst/n7238 ) );
  nnd2s1 \IDinst/U7262  ( .DIN1(\IDinst/RegFile[21][13] ), .DIN2(n1111), 
        .Q(\IDinst/n7237 ) );
  nnd2s1 \IDinst/U7261  ( .DIN1(\IDinst/RegFile[20][13] ), .DIN2(n1032), 
        .Q(\IDinst/n7236 ) );
  nnd2s1 \IDinst/U7260  ( .DIN1(\IDinst/n7234 ), .DIN2(\IDinst/n7233 ), 
        .Q(\IDinst/n7235 ) );
  nnd2s1 \IDinst/U7259  ( .DIN1(\IDinst/n7232 ), .DIN2(n1177), 
        .Q(\IDinst/n7234 ) );
  nnd2s1 \IDinst/U7258  ( .DIN1(\IDinst/n7229 ), .DIN2(n1135), 
        .Q(\IDinst/n7233 ) );
  nnd2s1 \IDinst/U7257  ( .DIN1(\IDinst/n7231 ), .DIN2(\IDinst/n7230 ), 
        .Q(\IDinst/n7232 ) );
  nnd2s1 \IDinst/U7256  ( .DIN1(\IDinst/RegFile[19][13] ), .DIN2(n1111), 
        .Q(\IDinst/n7231 ) );
  nnd2s1 \IDinst/U7255  ( .DIN1(\IDinst/RegFile[18][13] ), .DIN2(n1032), 
        .Q(\IDinst/n7230 ) );
  nnd2s1 \IDinst/U7254  ( .DIN1(\IDinst/n7228 ), .DIN2(\IDinst/n7227 ), 
        .Q(\IDinst/n7229 ) );
  nnd2s1 \IDinst/U7253  ( .DIN1(\IDinst/RegFile[17][13] ), .DIN2(n1111), 
        .Q(\IDinst/n7228 ) );
  nnd2s1 \IDinst/U7252  ( .DIN1(\IDinst/RegFile[16][13] ), .DIN2(n1032), 
        .Q(\IDinst/n7227 ) );
  nnd2s1 \IDinst/U7251  ( .DIN1(\IDinst/n7225 ), .DIN2(\IDinst/n7224 ), 
        .Q(\IDinst/n7226 ) );
  nnd2s1 \IDinst/U7250  ( .DIN1(\IDinst/n7223 ), .DIN2(n642), 
        .Q(\IDinst/n7225 ) );
  nnd2s1 \IDinst/U7249  ( .DIN1(\IDinst/n7202 ), .DIN2(n673), 
        .Q(\IDinst/n7224 ) );
  nnd2s1 \IDinst/U7248  ( .DIN1(\IDinst/n7222 ), .DIN2(\IDinst/n7221 ), 
        .Q(\IDinst/n7223 ) );
  nnd2s1 \IDinst/U7247  ( .DIN1(\IDinst/n7220 ), .DIN2(n1193), 
        .Q(\IDinst/n7222 ) );
  nnd2s1 \IDinst/U7246  ( .DIN1(\IDinst/n7211 ), .DIN2(n1184), 
        .Q(\IDinst/n7221 ) );
  nnd2s1 \IDinst/U7245  ( .DIN1(\IDinst/n7219 ), .DIN2(\IDinst/n7218 ), 
        .Q(\IDinst/n7220 ) );
  nnd2s1 \IDinst/U7244  ( .DIN1(\IDinst/n7217 ), .DIN2(n1177), 
        .Q(\IDinst/n7219 ) );
  nnd2s1 \IDinst/U7243  ( .DIN1(\IDinst/n7214 ), .DIN2(n1135), 
        .Q(\IDinst/n7218 ) );
  nnd2s1 \IDinst/U7242  ( .DIN1(\IDinst/n7216 ), .DIN2(\IDinst/n7215 ), 
        .Q(\IDinst/n7217 ) );
  nnd2s1 \IDinst/U7241  ( .DIN1(\IDinst/RegFile[15][13] ), .DIN2(n1111), 
        .Q(\IDinst/n7216 ) );
  nnd2s1 \IDinst/U7240  ( .DIN1(\IDinst/RegFile[14][13] ), .DIN2(n1032), 
        .Q(\IDinst/n7215 ) );
  nnd2s1 \IDinst/U7239  ( .DIN1(\IDinst/n7213 ), .DIN2(\IDinst/n7212 ), 
        .Q(\IDinst/n7214 ) );
  nnd2s1 \IDinst/U7238  ( .DIN1(\IDinst/RegFile[13][13] ), .DIN2(n1111), 
        .Q(\IDinst/n7213 ) );
  nnd2s1 \IDinst/U7237  ( .DIN1(\IDinst/RegFile[12][13] ), .DIN2(n1032), 
        .Q(\IDinst/n7212 ) );
  nnd2s1 \IDinst/U7236  ( .DIN1(\IDinst/n7210 ), .DIN2(\IDinst/n7209 ), 
        .Q(\IDinst/n7211 ) );
  nnd2s1 \IDinst/U7235  ( .DIN1(\IDinst/n7208 ), .DIN2(n1177), 
        .Q(\IDinst/n7210 ) );
  nnd2s1 \IDinst/U7234  ( .DIN1(\IDinst/n7205 ), .DIN2(n1135), 
        .Q(\IDinst/n7209 ) );
  nnd2s1 \IDinst/U7233  ( .DIN1(\IDinst/n7207 ), .DIN2(\IDinst/n7206 ), 
        .Q(\IDinst/n7208 ) );
  nnd2s1 \IDinst/U7232  ( .DIN1(\IDinst/RegFile[11][13] ), .DIN2(n1111), 
        .Q(\IDinst/n7207 ) );
  nnd2s1 \IDinst/U7231  ( .DIN1(\IDinst/RegFile[10][13] ), .DIN2(n1032), 
        .Q(\IDinst/n7206 ) );
  nnd2s1 \IDinst/U7230  ( .DIN1(\IDinst/n7204 ), .DIN2(\IDinst/n7203 ), 
        .Q(\IDinst/n7205 ) );
  nnd2s1 \IDinst/U7229  ( .DIN1(\IDinst/RegFile[9][13] ), .DIN2(n1112), 
        .Q(\IDinst/n7204 ) );
  nnd2s1 \IDinst/U7228  ( .DIN1(\IDinst/RegFile[8][13] ), .DIN2(n1032), 
        .Q(\IDinst/n7203 ) );
  nnd2s1 \IDinst/U7227  ( .DIN1(\IDinst/n7201 ), .DIN2(\IDinst/n7200 ), 
        .Q(\IDinst/n7202 ) );
  nnd2s1 \IDinst/U7226  ( .DIN1(\IDinst/n7199 ), .DIN2(n1193), 
        .Q(\IDinst/n7201 ) );
  nnd2s1 \IDinst/U7225  ( .DIN1(\IDinst/n7190 ), .DIN2(n1184), 
        .Q(\IDinst/n7200 ) );
  nnd2s1 \IDinst/U7224  ( .DIN1(\IDinst/n7198 ), .DIN2(\IDinst/n7197 ), 
        .Q(\IDinst/n7199 ) );
  nnd2s1 \IDinst/U7223  ( .DIN1(\IDinst/n7196 ), .DIN2(n1176), 
        .Q(\IDinst/n7198 ) );
  nnd2s1 \IDinst/U7222  ( .DIN1(\IDinst/n7193 ), .DIN2(n1135), 
        .Q(\IDinst/n7197 ) );
  nnd2s1 \IDinst/U7221  ( .DIN1(\IDinst/n7195 ), .DIN2(\IDinst/n7194 ), 
        .Q(\IDinst/n7196 ) );
  nnd2s1 \IDinst/U7220  ( .DIN1(\IDinst/RegFile[7][13] ), .DIN2(n1112), 
        .Q(\IDinst/n7195 ) );
  nnd2s1 \IDinst/U7219  ( .DIN1(\IDinst/RegFile[6][13] ), .DIN2(n1032), 
        .Q(\IDinst/n7194 ) );
  nnd2s1 \IDinst/U7218  ( .DIN1(\IDinst/n7192 ), .DIN2(\IDinst/n7191 ), 
        .Q(\IDinst/n7193 ) );
  nnd2s1 \IDinst/U7217  ( .DIN1(\IDinst/RegFile[5][13] ), .DIN2(n1112), 
        .Q(\IDinst/n7192 ) );
  nnd2s1 \IDinst/U7216  ( .DIN1(\IDinst/RegFile[4][13] ), .DIN2(n1032), 
        .Q(\IDinst/n7191 ) );
  nnd2s1 \IDinst/U7215  ( .DIN1(\IDinst/n7189 ), .DIN2(\IDinst/n7188 ), 
        .Q(\IDinst/n7190 ) );
  nnd2s1 \IDinst/U7214  ( .DIN1(\IDinst/n7187 ), .DIN2(n1176), 
        .Q(\IDinst/n7189 ) );
  nnd2s1 \IDinst/U7213  ( .DIN1(\IDinst/n7184 ), .DIN2(n1135), 
        .Q(\IDinst/n7188 ) );
  nnd2s1 \IDinst/U7212  ( .DIN1(\IDinst/n7186 ), .DIN2(\IDinst/n7185 ), 
        .Q(\IDinst/n7187 ) );
  nnd2s1 \IDinst/U7211  ( .DIN1(\IDinst/RegFile[3][13] ), .DIN2(n1112), 
        .Q(\IDinst/n7186 ) );
  nnd2s1 \IDinst/U7210  ( .DIN1(\IDinst/RegFile[2][13] ), .DIN2(n1031), 
        .Q(\IDinst/n7185 ) );
  nnd2s1 \IDinst/U7209  ( .DIN1(\IDinst/n7183 ), .DIN2(\IDinst/n7182 ), 
        .Q(\IDinst/n7184 ) );
  nnd2s1 \IDinst/U7208  ( .DIN1(\IDinst/RegFile[1][13] ), .DIN2(n1112), 
        .Q(\IDinst/n7183 ) );
  nnd2s1 \IDinst/U7207  ( .DIN1(\IDinst/RegFile[0][13] ), .DIN2(n1031), 
        .Q(\IDinst/n7182 ) );
  nnd2s1 \IDinst/U7206  ( .DIN1(\IDinst/n7181 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n5972 ) );
  nnd2s1 \IDinst/U7205  ( .DIN1(\IDinst/n7136 ), .DIN2(n636), 
        .Q(\IDinst/n5973 ) );
  nnd2s1 \IDinst/U7204  ( .DIN1(\IDinst/n7180 ), .DIN2(\IDinst/n7179 ), 
        .Q(\IDinst/n7181 ) );
  nnd2s1 \IDinst/U7203  ( .DIN1(\IDinst/n7178 ), .DIN2(n641), 
        .Q(\IDinst/n7180 ) );
  nnd2s1 \IDinst/U7202  ( .DIN1(\IDinst/n7157 ), .DIN2(n671), 
        .Q(\IDinst/n7179 ) );
  nnd2s1 \IDinst/U7201  ( .DIN1(\IDinst/n7177 ), .DIN2(\IDinst/n7176 ), 
        .Q(\IDinst/n7178 ) );
  nnd2s1 \IDinst/U7200  ( .DIN1(\IDinst/n7175 ), .DIN2(n1193), 
        .Q(\IDinst/n7177 ) );
  nnd2s1 \IDinst/U7199  ( .DIN1(\IDinst/n7166 ), .DIN2(n1184), 
        .Q(\IDinst/n7176 ) );
  nnd2s1 \IDinst/U7198  ( .DIN1(\IDinst/n7174 ), .DIN2(\IDinst/n7173 ), 
        .Q(\IDinst/n7175 ) );
  nnd2s1 \IDinst/U7197  ( .DIN1(\IDinst/n7172 ), .DIN2(n1176), 
        .Q(\IDinst/n7174 ) );
  nnd2s1 \IDinst/U7196  ( .DIN1(\IDinst/n7169 ), .DIN2(n1135), 
        .Q(\IDinst/n7173 ) );
  nnd2s1 \IDinst/U7195  ( .DIN1(\IDinst/n7171 ), .DIN2(\IDinst/n7170 ), 
        .Q(\IDinst/n7172 ) );
  nnd2s1 \IDinst/U7194  ( .DIN1(\IDinst/RegFile[31][12] ), .DIN2(n1112), 
        .Q(\IDinst/n7171 ) );
  nnd2s1 \IDinst/U7193  ( .DIN1(\IDinst/RegFile[30][12] ), .DIN2(n1031), 
        .Q(\IDinst/n7170 ) );
  nnd2s1 \IDinst/U7192  ( .DIN1(\IDinst/n7168 ), .DIN2(\IDinst/n7167 ), 
        .Q(\IDinst/n7169 ) );
  nnd2s1 \IDinst/U7191  ( .DIN1(\IDinst/RegFile[29][12] ), .DIN2(n1112), 
        .Q(\IDinst/n7168 ) );
  nnd2s1 \IDinst/U7190  ( .DIN1(\IDinst/RegFile[28][12] ), .DIN2(n1031), 
        .Q(\IDinst/n7167 ) );
  nnd2s1 \IDinst/U7189  ( .DIN1(\IDinst/n7165 ), .DIN2(\IDinst/n7164 ), 
        .Q(\IDinst/n7166 ) );
  nnd2s1 \IDinst/U7188  ( .DIN1(\IDinst/n7163 ), .DIN2(n1176), 
        .Q(\IDinst/n7165 ) );
  nnd2s1 \IDinst/U7187  ( .DIN1(\IDinst/n7160 ), .DIN2(n1135), 
        .Q(\IDinst/n7164 ) );
  nnd2s1 \IDinst/U7186  ( .DIN1(\IDinst/n7162 ), .DIN2(\IDinst/n7161 ), 
        .Q(\IDinst/n7163 ) );
  nnd2s1 \IDinst/U7185  ( .DIN1(\IDinst/RegFile[27][12] ), .DIN2(n1112), 
        .Q(\IDinst/n7162 ) );
  nnd2s1 \IDinst/U7184  ( .DIN1(\IDinst/RegFile[26][12] ), .DIN2(n1031), 
        .Q(\IDinst/n7161 ) );
  nnd2s1 \IDinst/U7183  ( .DIN1(\IDinst/n7159 ), .DIN2(\IDinst/n7158 ), 
        .Q(\IDinst/n7160 ) );
  nnd2s1 \IDinst/U7182  ( .DIN1(\IDinst/RegFile[25][12] ), .DIN2(n1112), 
        .Q(\IDinst/n7159 ) );
  nnd2s1 \IDinst/U7181  ( .DIN1(\IDinst/RegFile[24][12] ), .DIN2(n1031), 
        .Q(\IDinst/n7158 ) );
  nnd2s1 \IDinst/U7180  ( .DIN1(\IDinst/n7156 ), .DIN2(\IDinst/n7155 ), 
        .Q(\IDinst/n7157 ) );
  nnd2s1 \IDinst/U7179  ( .DIN1(\IDinst/n7154 ), .DIN2(n1193), 
        .Q(\IDinst/n7156 ) );
  nnd2s1 \IDinst/U7178  ( .DIN1(\IDinst/n7145 ), .DIN2(n1184), 
        .Q(\IDinst/n7155 ) );
  nnd2s1 \IDinst/U7177  ( .DIN1(\IDinst/n7153 ), .DIN2(\IDinst/n7152 ), 
        .Q(\IDinst/n7154 ) );
  nnd2s1 \IDinst/U7176  ( .DIN1(\IDinst/n7151 ), .DIN2(n1176), 
        .Q(\IDinst/n7153 ) );
  nnd2s1 \IDinst/U7175  ( .DIN1(\IDinst/n7148 ), .DIN2(n1135), 
        .Q(\IDinst/n7152 ) );
  nnd2s1 \IDinst/U7174  ( .DIN1(\IDinst/n7150 ), .DIN2(\IDinst/n7149 ), 
        .Q(\IDinst/n7151 ) );
  nnd2s1 \IDinst/U7173  ( .DIN1(\IDinst/RegFile[23][12] ), .DIN2(n1113), 
        .Q(\IDinst/n7150 ) );
  nnd2s1 \IDinst/U7172  ( .DIN1(\IDinst/RegFile[22][12] ), .DIN2(n1031), 
        .Q(\IDinst/n7149 ) );
  nnd2s1 \IDinst/U7171  ( .DIN1(\IDinst/n7147 ), .DIN2(\IDinst/n7146 ), 
        .Q(\IDinst/n7148 ) );
  nnd2s1 \IDinst/U7170  ( .DIN1(\IDinst/RegFile[21][12] ), .DIN2(n1113), 
        .Q(\IDinst/n7147 ) );
  nnd2s1 \IDinst/U7169  ( .DIN1(\IDinst/RegFile[20][12] ), .DIN2(n1031), 
        .Q(\IDinst/n7146 ) );
  nnd2s1 \IDinst/U7168  ( .DIN1(\IDinst/n7144 ), .DIN2(\IDinst/n7143 ), 
        .Q(\IDinst/n7145 ) );
  nnd2s1 \IDinst/U7167  ( .DIN1(\IDinst/n7142 ), .DIN2(n1176), 
        .Q(\IDinst/n7144 ) );
  nnd2s1 \IDinst/U7166  ( .DIN1(\IDinst/n7139 ), .DIN2(n1135), 
        .Q(\IDinst/n7143 ) );
  nnd2s1 \IDinst/U7165  ( .DIN1(\IDinst/n7141 ), .DIN2(\IDinst/n7140 ), 
        .Q(\IDinst/n7142 ) );
  nnd2s1 \IDinst/U7164  ( .DIN1(\IDinst/RegFile[19][12] ), .DIN2(n1113), 
        .Q(\IDinst/n7141 ) );
  nnd2s1 \IDinst/U7163  ( .DIN1(\IDinst/RegFile[18][12] ), .DIN2(n1031), 
        .Q(\IDinst/n7140 ) );
  nnd2s1 \IDinst/U7162  ( .DIN1(\IDinst/n7138 ), .DIN2(\IDinst/n7137 ), 
        .Q(\IDinst/n7139 ) );
  nnd2s1 \IDinst/U7161  ( .DIN1(\IDinst/RegFile[17][12] ), .DIN2(n1113), 
        .Q(\IDinst/n7138 ) );
  nnd2s1 \IDinst/U7160  ( .DIN1(\IDinst/RegFile[16][12] ), .DIN2(n1031), 
        .Q(\IDinst/n7137 ) );
  nnd2s1 \IDinst/U7159  ( .DIN1(\IDinst/n7135 ), .DIN2(\IDinst/n7134 ), 
        .Q(\IDinst/n7136 ) );
  nnd2s1 \IDinst/U7158  ( .DIN1(\IDinst/n7133 ), .DIN2(n644), 
        .Q(\IDinst/n7135 ) );
  nnd2s1 \IDinst/U7157  ( .DIN1(\IDinst/n7112 ), .DIN2(n672), 
        .Q(\IDinst/n7134 ) );
  nnd2s1 \IDinst/U7156  ( .DIN1(\IDinst/n7132 ), .DIN2(\IDinst/n7131 ), 
        .Q(\IDinst/n7133 ) );
  nnd2s1 \IDinst/U7155  ( .DIN1(\IDinst/n7130 ), .DIN2(n1193), 
        .Q(\IDinst/n7132 ) );
  nnd2s1 \IDinst/U7154  ( .DIN1(\IDinst/n7121 ), .DIN2(n1184), 
        .Q(\IDinst/n7131 ) );
  nnd2s1 \IDinst/U7153  ( .DIN1(\IDinst/n7129 ), .DIN2(\IDinst/n7128 ), 
        .Q(\IDinst/n7130 ) );
  nnd2s1 \IDinst/U7152  ( .DIN1(\IDinst/n7127 ), .DIN2(n1176), 
        .Q(\IDinst/n7129 ) );
  nnd2s1 \IDinst/U7151  ( .DIN1(\IDinst/n7124 ), .DIN2(n1135), 
        .Q(\IDinst/n7128 ) );
  nnd2s1 \IDinst/U7150  ( .DIN1(\IDinst/n7126 ), .DIN2(\IDinst/n7125 ), 
        .Q(\IDinst/n7127 ) );
  nnd2s1 \IDinst/U7149  ( .DIN1(\IDinst/RegFile[15][12] ), .DIN2(n1113), 
        .Q(\IDinst/n7126 ) );
  nnd2s1 \IDinst/U7148  ( .DIN1(\IDinst/RegFile[14][12] ), .DIN2(n1031), 
        .Q(\IDinst/n7125 ) );
  nnd2s1 \IDinst/U7147  ( .DIN1(\IDinst/n7123 ), .DIN2(\IDinst/n7122 ), 
        .Q(\IDinst/n7124 ) );
  nnd2s1 \IDinst/U7146  ( .DIN1(\IDinst/RegFile[13][12] ), .DIN2(n1113), 
        .Q(\IDinst/n7123 ) );
  nnd2s1 \IDinst/U7145  ( .DIN1(\IDinst/RegFile[12][12] ), .DIN2(n1031), 
        .Q(\IDinst/n7122 ) );
  nnd2s1 \IDinst/U7144  ( .DIN1(\IDinst/n7120 ), .DIN2(\IDinst/n7119 ), 
        .Q(\IDinst/n7121 ) );
  nnd2s1 \IDinst/U7143  ( .DIN1(\IDinst/n7118 ), .DIN2(n1176), 
        .Q(\IDinst/n7120 ) );
  nnd2s1 \IDinst/U7142  ( .DIN1(\IDinst/n7115 ), .DIN2(n1136), 
        .Q(\IDinst/n7119 ) );
  nnd2s1 \IDinst/U7141  ( .DIN1(\IDinst/n7117 ), .DIN2(\IDinst/n7116 ), 
        .Q(\IDinst/n7118 ) );
  nnd2s1 \IDinst/U7140  ( .DIN1(\IDinst/RegFile[11][12] ), .DIN2(n1113), 
        .Q(\IDinst/n7117 ) );
  nnd2s1 \IDinst/U7139  ( .DIN1(\IDinst/RegFile[10][12] ), .DIN2(n1031), 
        .Q(\IDinst/n7116 ) );
  nnd2s1 \IDinst/U7138  ( .DIN1(\IDinst/n7114 ), .DIN2(\IDinst/n7113 ), 
        .Q(\IDinst/n7115 ) );
  nnd2s1 \IDinst/U7137  ( .DIN1(\IDinst/RegFile[9][12] ), .DIN2(n1113), 
        .Q(\IDinst/n7114 ) );
  nnd2s1 \IDinst/U7136  ( .DIN1(\IDinst/RegFile[8][12] ), .DIN2(n1030), 
        .Q(\IDinst/n7113 ) );
  nnd2s1 \IDinst/U7135  ( .DIN1(\IDinst/n7111 ), .DIN2(\IDinst/n7110 ), 
        .Q(\IDinst/n7112 ) );
  nnd2s1 \IDinst/U7134  ( .DIN1(\IDinst/n7109 ), .DIN2(n1193), 
        .Q(\IDinst/n7111 ) );
  nnd2s1 \IDinst/U7133  ( .DIN1(\IDinst/n7100 ), .DIN2(n1184), 
        .Q(\IDinst/n7110 ) );
  nnd2s1 \IDinst/U7132  ( .DIN1(\IDinst/n7108 ), .DIN2(\IDinst/n7107 ), 
        .Q(\IDinst/n7109 ) );
  nnd2s1 \IDinst/U7131  ( .DIN1(\IDinst/n7106 ), .DIN2(n1176), 
        .Q(\IDinst/n7108 ) );
  nnd2s1 \IDinst/U7130  ( .DIN1(\IDinst/n7103 ), .DIN2(n1136), 
        .Q(\IDinst/n7107 ) );
  nnd2s1 \IDinst/U7129  ( .DIN1(\IDinst/n7105 ), .DIN2(\IDinst/n7104 ), 
        .Q(\IDinst/n7106 ) );
  nnd2s1 \IDinst/U7128  ( .DIN1(\IDinst/RegFile[7][12] ), .DIN2(n1113), 
        .Q(\IDinst/n7105 ) );
  nnd2s1 \IDinst/U7127  ( .DIN1(\IDinst/RegFile[6][12] ), .DIN2(n1030), 
        .Q(\IDinst/n7104 ) );
  nnd2s1 \IDinst/U7126  ( .DIN1(\IDinst/n7102 ), .DIN2(\IDinst/n7101 ), 
        .Q(\IDinst/n7103 ) );
  nnd2s1 \IDinst/U7125  ( .DIN1(\IDinst/RegFile[5][12] ), .DIN2(n1114), 
        .Q(\IDinst/n7102 ) );
  nnd2s1 \IDinst/U7124  ( .DIN1(\IDinst/RegFile[4][12] ), .DIN2(n1030), 
        .Q(\IDinst/n7101 ) );
  nnd2s1 \IDinst/U7123  ( .DIN1(\IDinst/n7099 ), .DIN2(\IDinst/n7098 ), 
        .Q(\IDinst/n7100 ) );
  nnd2s1 \IDinst/U7122  ( .DIN1(\IDinst/n7097 ), .DIN2(n1175), 
        .Q(\IDinst/n7099 ) );
  nnd2s1 \IDinst/U7121  ( .DIN1(\IDinst/n7094 ), .DIN2(n1136), 
        .Q(\IDinst/n7098 ) );
  nnd2s1 \IDinst/U7120  ( .DIN1(\IDinst/n7096 ), .DIN2(\IDinst/n7095 ), 
        .Q(\IDinst/n7097 ) );
  nnd2s1 \IDinst/U7119  ( .DIN1(\IDinst/RegFile[3][12] ), .DIN2(n1114), 
        .Q(\IDinst/n7096 ) );
  nnd2s1 \IDinst/U7118  ( .DIN1(\IDinst/RegFile[2][12] ), .DIN2(n1030), 
        .Q(\IDinst/n7095 ) );
  nnd2s1 \IDinst/U7117  ( .DIN1(\IDinst/n7093 ), .DIN2(\IDinst/n7092 ), 
        .Q(\IDinst/n7094 ) );
  nnd2s1 \IDinst/U7116  ( .DIN1(\IDinst/RegFile[1][12] ), .DIN2(n1114), 
        .Q(\IDinst/n7093 ) );
  nnd2s1 \IDinst/U7115  ( .DIN1(\IDinst/RegFile[0][12] ), .DIN2(n1030), 
        .Q(\IDinst/n7092 ) );
  nnd2s1 \IDinst/U7114  ( .DIN1(\IDinst/n7091 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n5970 ) );
  nnd2s1 \IDinst/U7113  ( .DIN1(\IDinst/n7046 ), .DIN2(n635), 
        .Q(\IDinst/n5971 ) );
  nnd2s1 \IDinst/U7112  ( .DIN1(\IDinst/n7090 ), .DIN2(\IDinst/n7089 ), 
        .Q(\IDinst/n7091 ) );
  nnd2s1 \IDinst/U7111  ( .DIN1(\IDinst/n7088 ), .DIN2(n643), 
        .Q(\IDinst/n7090 ) );
  nnd2s1 \IDinst/U7110  ( .DIN1(\IDinst/n7067 ), .DIN2(n670), 
        .Q(\IDinst/n7089 ) );
  nnd2s1 \IDinst/U7109  ( .DIN1(\IDinst/n7087 ), .DIN2(\IDinst/n7086 ), 
        .Q(\IDinst/n7088 ) );
  nnd2s1 \IDinst/U7108  ( .DIN1(\IDinst/n7085 ), .DIN2(n1193), 
        .Q(\IDinst/n7087 ) );
  nnd2s1 \IDinst/U7107  ( .DIN1(\IDinst/n7076 ), .DIN2(n1184), 
        .Q(\IDinst/n7086 ) );
  nnd2s1 \IDinst/U7106  ( .DIN1(\IDinst/n7084 ), .DIN2(\IDinst/n7083 ), 
        .Q(\IDinst/n7085 ) );
  nnd2s1 \IDinst/U7105  ( .DIN1(\IDinst/n7082 ), .DIN2(n1175), 
        .Q(\IDinst/n7084 ) );
  nnd2s1 \IDinst/U7104  ( .DIN1(\IDinst/n7079 ), .DIN2(n1136), 
        .Q(\IDinst/n7083 ) );
  nnd2s1 \IDinst/U7103  ( .DIN1(\IDinst/n7081 ), .DIN2(\IDinst/n7080 ), 
        .Q(\IDinst/n7082 ) );
  nnd2s1 \IDinst/U7102  ( .DIN1(\IDinst/RegFile[31][11] ), .DIN2(n1114), 
        .Q(\IDinst/n7081 ) );
  nnd2s1 \IDinst/U7101  ( .DIN1(\IDinst/RegFile[30][11] ), .DIN2(n1030), 
        .Q(\IDinst/n7080 ) );
  nnd2s1 \IDinst/U7100  ( .DIN1(\IDinst/n7078 ), .DIN2(\IDinst/n7077 ), 
        .Q(\IDinst/n7079 ) );
  nnd2s1 \IDinst/U7099  ( .DIN1(\IDinst/RegFile[29][11] ), .DIN2(n1114), 
        .Q(\IDinst/n7078 ) );
  nnd2s1 \IDinst/U7098  ( .DIN1(\IDinst/RegFile[28][11] ), .DIN2(n1030), 
        .Q(\IDinst/n7077 ) );
  nnd2s1 \IDinst/U7097  ( .DIN1(\IDinst/n7075 ), .DIN2(\IDinst/n7074 ), 
        .Q(\IDinst/n7076 ) );
  nnd2s1 \IDinst/U7096  ( .DIN1(\IDinst/n7073 ), .DIN2(n1175), 
        .Q(\IDinst/n7075 ) );
  nnd2s1 \IDinst/U7095  ( .DIN1(\IDinst/n7070 ), .DIN2(n1136), 
        .Q(\IDinst/n7074 ) );
  nnd2s1 \IDinst/U7094  ( .DIN1(\IDinst/n7072 ), .DIN2(\IDinst/n7071 ), 
        .Q(\IDinst/n7073 ) );
  nnd2s1 \IDinst/U7093  ( .DIN1(\IDinst/RegFile[27][11] ), .DIN2(n1114), 
        .Q(\IDinst/n7072 ) );
  nnd2s1 \IDinst/U7092  ( .DIN1(\IDinst/RegFile[26][11] ), .DIN2(n1030), 
        .Q(\IDinst/n7071 ) );
  nnd2s1 \IDinst/U7091  ( .DIN1(\IDinst/n7069 ), .DIN2(\IDinst/n7068 ), 
        .Q(\IDinst/n7070 ) );
  nnd2s1 \IDinst/U7090  ( .DIN1(\IDinst/RegFile[25][11] ), .DIN2(n1114), 
        .Q(\IDinst/n7069 ) );
  nnd2s1 \IDinst/U7089  ( .DIN1(\IDinst/RegFile[24][11] ), .DIN2(n1030), 
        .Q(\IDinst/n7068 ) );
  nnd2s1 \IDinst/U7088  ( .DIN1(\IDinst/n7066 ), .DIN2(\IDinst/n7065 ), 
        .Q(\IDinst/n7067 ) );
  nnd2s1 \IDinst/U7087  ( .DIN1(\IDinst/n7064 ), .DIN2(n1193), 
        .Q(\IDinst/n7066 ) );
  nnd2s1 \IDinst/U7086  ( .DIN1(\IDinst/n7055 ), .DIN2(n1184), 
        .Q(\IDinst/n7065 ) );
  nnd2s1 \IDinst/U7085  ( .DIN1(\IDinst/n7063 ), .DIN2(\IDinst/n7062 ), 
        .Q(\IDinst/n7064 ) );
  nnd2s1 \IDinst/U7084  ( .DIN1(\IDinst/n7061 ), .DIN2(n1175), 
        .Q(\IDinst/n7063 ) );
  nnd2s1 \IDinst/U7083  ( .DIN1(\IDinst/n7058 ), .DIN2(n1136), 
        .Q(\IDinst/n7062 ) );
  nnd2s1 \IDinst/U7082  ( .DIN1(\IDinst/n7060 ), .DIN2(\IDinst/n7059 ), 
        .Q(\IDinst/n7061 ) );
  nnd2s1 \IDinst/U7081  ( .DIN1(\IDinst/RegFile[23][11] ), .DIN2(n1114), 
        .Q(\IDinst/n7060 ) );
  nnd2s1 \IDinst/U7080  ( .DIN1(\IDinst/RegFile[22][11] ), .DIN2(n1030), 
        .Q(\IDinst/n7059 ) );
  nnd2s1 \IDinst/U7079  ( .DIN1(\IDinst/n7057 ), .DIN2(\IDinst/n7056 ), 
        .Q(\IDinst/n7058 ) );
  nnd2s1 \IDinst/U7078  ( .DIN1(\IDinst/RegFile[21][11] ), .DIN2(n1114), 
        .Q(\IDinst/n7057 ) );
  nnd2s1 \IDinst/U7077  ( .DIN1(\IDinst/RegFile[20][11] ), .DIN2(n1030), 
        .Q(\IDinst/n7056 ) );
  nnd2s1 \IDinst/U7076  ( .DIN1(\IDinst/n7054 ), .DIN2(\IDinst/n7053 ), 
        .Q(\IDinst/n7055 ) );
  nnd2s1 \IDinst/U7075  ( .DIN1(\IDinst/n7052 ), .DIN2(n1175), 
        .Q(\IDinst/n7054 ) );
  nnd2s1 \IDinst/U7074  ( .DIN1(\IDinst/n7049 ), .DIN2(n1136), 
        .Q(\IDinst/n7053 ) );
  nnd2s1 \IDinst/U7073  ( .DIN1(\IDinst/n7051 ), .DIN2(\IDinst/n7050 ), 
        .Q(\IDinst/n7052 ) );
  nnd2s1 \IDinst/U7072  ( .DIN1(\IDinst/RegFile[19][11] ), .DIN2(n1115), 
        .Q(\IDinst/n7051 ) );
  nnd2s1 \IDinst/U7071  ( .DIN1(\IDinst/RegFile[18][11] ), .DIN2(n1030), 
        .Q(\IDinst/n7050 ) );
  nnd2s1 \IDinst/U7070  ( .DIN1(\IDinst/n7048 ), .DIN2(\IDinst/n7047 ), 
        .Q(\IDinst/n7049 ) );
  nnd2s1 \IDinst/U7069  ( .DIN1(\IDinst/RegFile[17][11] ), .DIN2(n1115), 
        .Q(\IDinst/n7048 ) );
  nnd2s1 \IDinst/U7068  ( .DIN1(\IDinst/RegFile[16][11] ), .DIN2(n1029), 
        .Q(\IDinst/n7047 ) );
  nnd2s1 \IDinst/U7067  ( .DIN1(\IDinst/n7045 ), .DIN2(\IDinst/n7044 ), 
        .Q(\IDinst/n7046 ) );
  nnd2s1 \IDinst/U7066  ( .DIN1(\IDinst/n7043 ), .DIN2(n642), 
        .Q(\IDinst/n7045 ) );
  nnd2s1 \IDinst/U7065  ( .DIN1(\IDinst/n7022 ), .DIN2(n673), 
        .Q(\IDinst/n7044 ) );
  nnd2s1 \IDinst/U7064  ( .DIN1(\IDinst/n7042 ), .DIN2(\IDinst/n7041 ), 
        .Q(\IDinst/n7043 ) );
  nnd2s1 \IDinst/U7063  ( .DIN1(\IDinst/n7040 ), .DIN2(n1190), 
        .Q(\IDinst/n7042 ) );
  nnd2s1 \IDinst/U7062  ( .DIN1(\IDinst/n7031 ), .DIN2(n1184), 
        .Q(\IDinst/n7041 ) );
  nnd2s1 \IDinst/U7061  ( .DIN1(\IDinst/n7039 ), .DIN2(\IDinst/n7038 ), 
        .Q(\IDinst/n7040 ) );
  nnd2s1 \IDinst/U7060  ( .DIN1(\IDinst/n7037 ), .DIN2(n1175), 
        .Q(\IDinst/n7039 ) );
  nnd2s1 \IDinst/U7059  ( .DIN1(\IDinst/n7034 ), .DIN2(n1136), 
        .Q(\IDinst/n7038 ) );
  nnd2s1 \IDinst/U7058  ( .DIN1(\IDinst/n7036 ), .DIN2(\IDinst/n7035 ), 
        .Q(\IDinst/n7037 ) );
  nnd2s1 \IDinst/U7057  ( .DIN1(\IDinst/RegFile[15][11] ), .DIN2(n1115), 
        .Q(\IDinst/n7036 ) );
  nnd2s1 \IDinst/U7056  ( .DIN1(\IDinst/RegFile[14][11] ), .DIN2(n1029), 
        .Q(\IDinst/n7035 ) );
  nnd2s1 \IDinst/U7055  ( .DIN1(\IDinst/n7033 ), .DIN2(\IDinst/n7032 ), 
        .Q(\IDinst/n7034 ) );
  nnd2s1 \IDinst/U7054  ( .DIN1(\IDinst/RegFile[13][11] ), .DIN2(n1115), 
        .Q(\IDinst/n7033 ) );
  nnd2s1 \IDinst/U7053  ( .DIN1(\IDinst/RegFile[12][11] ), .DIN2(n1029), 
        .Q(\IDinst/n7032 ) );
  nnd2s1 \IDinst/U7052  ( .DIN1(\IDinst/n7030 ), .DIN2(\IDinst/n7029 ), 
        .Q(\IDinst/n7031 ) );
  nnd2s1 \IDinst/U7051  ( .DIN1(\IDinst/n7028 ), .DIN2(n1175), 
        .Q(\IDinst/n7030 ) );
  nnd2s1 \IDinst/U7050  ( .DIN1(\IDinst/n7025 ), .DIN2(n1136), 
        .Q(\IDinst/n7029 ) );
  nnd2s1 \IDinst/U7049  ( .DIN1(\IDinst/n7027 ), .DIN2(\IDinst/n7026 ), 
        .Q(\IDinst/n7028 ) );
  nnd2s1 \IDinst/U7048  ( .DIN1(\IDinst/RegFile[11][11] ), .DIN2(n1115), 
        .Q(\IDinst/n7027 ) );
  nnd2s1 \IDinst/U7047  ( .DIN1(\IDinst/RegFile[10][11] ), .DIN2(n1029), 
        .Q(\IDinst/n7026 ) );
  nnd2s1 \IDinst/U7046  ( .DIN1(\IDinst/n7024 ), .DIN2(\IDinst/n7023 ), 
        .Q(\IDinst/n7025 ) );
  nnd2s1 \IDinst/U7045  ( .DIN1(\IDinst/RegFile[9][11] ), .DIN2(n1115), 
        .Q(\IDinst/n7024 ) );
  nnd2s1 \IDinst/U7044  ( .DIN1(\IDinst/RegFile[8][11] ), .DIN2(n1029), 
        .Q(\IDinst/n7023 ) );
  nnd2s1 \IDinst/U7043  ( .DIN1(\IDinst/n7021 ), .DIN2(\IDinst/n7020 ), 
        .Q(\IDinst/n7022 ) );
  nnd2s1 \IDinst/U7042  ( .DIN1(\IDinst/n7019 ), .DIN2(n1194), 
        .Q(\IDinst/n7021 ) );
  nnd2s1 \IDinst/U7041  ( .DIN1(\IDinst/n7010 ), .DIN2(n1183), 
        .Q(\IDinst/n7020 ) );
  nnd2s1 \IDinst/U7040  ( .DIN1(\IDinst/n7018 ), .DIN2(\IDinst/n7017 ), 
        .Q(\IDinst/n7019 ) );
  nnd2s1 \IDinst/U7039  ( .DIN1(\IDinst/n7016 ), .DIN2(n1175), 
        .Q(\IDinst/n7018 ) );
  nnd2s1 \IDinst/U7038  ( .DIN1(\IDinst/n7013 ), .DIN2(n1136), 
        .Q(\IDinst/n7017 ) );
  nnd2s1 \IDinst/U7037  ( .DIN1(\IDinst/n7015 ), .DIN2(\IDinst/n7014 ), 
        .Q(\IDinst/n7016 ) );
  nnd2s1 \IDinst/U7036  ( .DIN1(\IDinst/RegFile[7][11] ), .DIN2(n1115), 
        .Q(\IDinst/n7015 ) );
  nnd2s1 \IDinst/U7035  ( .DIN1(\IDinst/RegFile[6][11] ), .DIN2(n1029), 
        .Q(\IDinst/n7014 ) );
  nnd2s1 \IDinst/U7034  ( .DIN1(\IDinst/n7012 ), .DIN2(\IDinst/n7011 ), 
        .Q(\IDinst/n7013 ) );
  nnd2s1 \IDinst/U7033  ( .DIN1(\IDinst/RegFile[5][11] ), .DIN2(n1115), 
        .Q(\IDinst/n7012 ) );
  nnd2s1 \IDinst/U7032  ( .DIN1(\IDinst/RegFile[4][11] ), .DIN2(n1029), 
        .Q(\IDinst/n7011 ) );
  nnd2s1 \IDinst/U7031  ( .DIN1(\IDinst/n7009 ), .DIN2(\IDinst/n7008 ), 
        .Q(\IDinst/n7010 ) );
  nnd2s1 \IDinst/U7030  ( .DIN1(\IDinst/n7007 ), .DIN2(n1175), 
        .Q(\IDinst/n7009 ) );
  nnd2s1 \IDinst/U7029  ( .DIN1(\IDinst/n7004 ), .DIN2(n1136), 
        .Q(\IDinst/n7008 ) );
  nnd2s1 \IDinst/U7028  ( .DIN1(\IDinst/n7006 ), .DIN2(\IDinst/n7005 ), 
        .Q(\IDinst/n7007 ) );
  nnd2s1 \IDinst/U7027  ( .DIN1(\IDinst/RegFile[3][11] ), .DIN2(n1115), 
        .Q(\IDinst/n7006 ) );
  nnd2s1 \IDinst/U7026  ( .DIN1(\IDinst/RegFile[2][11] ), .DIN2(n1029), 
        .Q(\IDinst/n7005 ) );
  nnd2s1 \IDinst/U7025  ( .DIN1(\IDinst/n7003 ), .DIN2(\IDinst/n7002 ), 
        .Q(\IDinst/n7004 ) );
  nnd2s1 \IDinst/U7024  ( .DIN1(\IDinst/RegFile[1][11] ), .DIN2(n1116), 
        .Q(\IDinst/n7003 ) );
  nnd2s1 \IDinst/U7023  ( .DIN1(\IDinst/RegFile[0][11] ), .DIN2(n1029), 
        .Q(\IDinst/n7002 ) );
  nnd2s1 \IDinst/U7022  ( .DIN1(\IDinst/n7001 ), .DIN2(n539), 
        .Q(\IDinst/n5968 ) );
  nnd2s1 \IDinst/U7021  ( .DIN1(\IDinst/n6956 ), .DIN2(n636), 
        .Q(\IDinst/n5969 ) );
  nnd2s1 \IDinst/U7020  ( .DIN1(\IDinst/n7000 ), .DIN2(\IDinst/n6999 ), 
        .Q(\IDinst/n7001 ) );
  nnd2s1 \IDinst/U7019  ( .DIN1(\IDinst/n6998 ), .DIN2(n641), 
        .Q(\IDinst/n7000 ) );
  nnd2s1 \IDinst/U7018  ( .DIN1(\IDinst/n6977 ), .DIN2(n671), 
        .Q(\IDinst/n6999 ) );
  nnd2s1 \IDinst/U7017  ( .DIN1(\IDinst/n6997 ), .DIN2(\IDinst/n6996 ), 
        .Q(\IDinst/n6998 ) );
  nnd2s1 \IDinst/U7016  ( .DIN1(\IDinst/n6995 ), .DIN2(n1197), 
        .Q(\IDinst/n6997 ) );
  nnd2s1 \IDinst/U7015  ( .DIN1(\IDinst/n6986 ), .DIN2(n1183), 
        .Q(\IDinst/n6996 ) );
  nnd2s1 \IDinst/U7014  ( .DIN1(\IDinst/n6994 ), .DIN2(\IDinst/n6993 ), 
        .Q(\IDinst/n6995 ) );
  nnd2s1 \IDinst/U7013  ( .DIN1(\IDinst/n6992 ), .DIN2(n1174), 
        .Q(\IDinst/n6994 ) );
  nnd2s1 \IDinst/U7012  ( .DIN1(\IDinst/n6989 ), .DIN2(n1136), 
        .Q(\IDinst/n6993 ) );
  nnd2s1 \IDinst/U7011  ( .DIN1(\IDinst/n6991 ), .DIN2(\IDinst/n6990 ), 
        .Q(\IDinst/n6992 ) );
  nnd2s1 \IDinst/U7010  ( .DIN1(\IDinst/RegFile[31][10] ), .DIN2(n1122), 
        .Q(\IDinst/n6991 ) );
  nnd2s1 \IDinst/U7009  ( .DIN1(\IDinst/RegFile[30][10] ), .DIN2(n1029), 
        .Q(\IDinst/n6990 ) );
  nnd2s1 \IDinst/U7008  ( .DIN1(\IDinst/n6988 ), .DIN2(\IDinst/n6987 ), 
        .Q(\IDinst/n6989 ) );
  nnd2s1 \IDinst/U7007  ( .DIN1(\IDinst/RegFile[29][10] ), .DIN2(n1122), 
        .Q(\IDinst/n6988 ) );
  nnd2s1 \IDinst/U7006  ( .DIN1(\IDinst/RegFile[28][10] ), .DIN2(n1029), 
        .Q(\IDinst/n6987 ) );
  nnd2s1 \IDinst/U7005  ( .DIN1(\IDinst/n6985 ), .DIN2(\IDinst/n6984 ), 
        .Q(\IDinst/n6986 ) );
  nnd2s1 \IDinst/U7004  ( .DIN1(\IDinst/n6983 ), .DIN2(n1174), 
        .Q(\IDinst/n6985 ) );
  nnd2s1 \IDinst/U7003  ( .DIN1(\IDinst/n6980 ), .DIN2(n1136), 
        .Q(\IDinst/n6984 ) );
  nnd2s1 \IDinst/U7002  ( .DIN1(\IDinst/n6982 ), .DIN2(\IDinst/n6981 ), 
        .Q(\IDinst/n6983 ) );
  nnd2s1 \IDinst/U7001  ( .DIN1(\IDinst/RegFile[27][10] ), .DIN2(n1122), 
        .Q(\IDinst/n6982 ) );
  nnd2s1 \IDinst/U7000  ( .DIN1(\IDinst/RegFile[26][10] ), .DIN2(n1029), 
        .Q(\IDinst/n6981 ) );
  nnd2s1 \IDinst/U6999  ( .DIN1(\IDinst/n6979 ), .DIN2(\IDinst/n6978 ), 
        .Q(\IDinst/n6980 ) );
  nnd2s1 \IDinst/U6998  ( .DIN1(\IDinst/RegFile[25][10] ), .DIN2(n1122), 
        .Q(\IDinst/n6979 ) );
  nnd2s1 \IDinst/U6997  ( .DIN1(\IDinst/RegFile[24][10] ), .DIN2(n1029), 
        .Q(\IDinst/n6978 ) );
  nnd2s1 \IDinst/U6996  ( .DIN1(\IDinst/n6976 ), .DIN2(\IDinst/n6975 ), 
        .Q(\IDinst/n6977 ) );
  nnd2s1 \IDinst/U6995  ( .DIN1(\IDinst/n6974 ), .DIN2(n1196), 
        .Q(\IDinst/n6976 ) );
  nnd2s1 \IDinst/U6994  ( .DIN1(\IDinst/n6965 ), .DIN2(n1183), 
        .Q(\IDinst/n6975 ) );
  nnd2s1 \IDinst/U6993  ( .DIN1(\IDinst/n6973 ), .DIN2(\IDinst/n6972 ), 
        .Q(\IDinst/n6974 ) );
  nnd2s1 \IDinst/U6992  ( .DIN1(\IDinst/n6971 ), .DIN2(n1174), 
        .Q(\IDinst/n6973 ) );
  nnd2s1 \IDinst/U6991  ( .DIN1(\IDinst/n6968 ), .DIN2(n1137), 
        .Q(\IDinst/n6972 ) );
  nnd2s1 \IDinst/U6990  ( .DIN1(\IDinst/n6970 ), .DIN2(\IDinst/n6969 ), 
        .Q(\IDinst/n6971 ) );
  nnd2s1 \IDinst/U6989  ( .DIN1(\IDinst/RegFile[23][10] ), .DIN2(n1122), 
        .Q(\IDinst/n6970 ) );
  nnd2s1 \IDinst/U6988  ( .DIN1(\IDinst/RegFile[22][10] ), .DIN2(n1028), 
        .Q(\IDinst/n6969 ) );
  nnd2s1 \IDinst/U6987  ( .DIN1(\IDinst/n6967 ), .DIN2(\IDinst/n6966 ), 
        .Q(\IDinst/n6968 ) );
  nnd2s1 \IDinst/U6986  ( .DIN1(\IDinst/RegFile[21][10] ), .DIN2(n1122), 
        .Q(\IDinst/n6967 ) );
  nnd2s1 \IDinst/U6985  ( .DIN1(\IDinst/RegFile[20][10] ), .DIN2(n1028), 
        .Q(\IDinst/n6966 ) );
  nnd2s1 \IDinst/U6984  ( .DIN1(\IDinst/n6964 ), .DIN2(\IDinst/n6963 ), 
        .Q(\IDinst/n6965 ) );
  nnd2s1 \IDinst/U6983  ( .DIN1(\IDinst/n6962 ), .DIN2(n1174), 
        .Q(\IDinst/n6964 ) );
  nnd2s1 \IDinst/U6982  ( .DIN1(\IDinst/n6959 ), .DIN2(n1137), 
        .Q(\IDinst/n6963 ) );
  nnd2s1 \IDinst/U6981  ( .DIN1(\IDinst/n6961 ), .DIN2(\IDinst/n6960 ), 
        .Q(\IDinst/n6962 ) );
  nnd2s1 \IDinst/U6980  ( .DIN1(\IDinst/RegFile[19][10] ), .DIN2(n1121), 
        .Q(\IDinst/n6961 ) );
  nnd2s1 \IDinst/U6979  ( .DIN1(\IDinst/RegFile[18][10] ), .DIN2(n1028), 
        .Q(\IDinst/n6960 ) );
  nnd2s1 \IDinst/U6978  ( .DIN1(\IDinst/n6958 ), .DIN2(\IDinst/n6957 ), 
        .Q(\IDinst/n6959 ) );
  nnd2s1 \IDinst/U6977  ( .DIN1(\IDinst/RegFile[17][10] ), .DIN2(n1121), 
        .Q(\IDinst/n6958 ) );
  nnd2s1 \IDinst/U6976  ( .DIN1(\IDinst/RegFile[16][10] ), .DIN2(n1028), 
        .Q(\IDinst/n6957 ) );
  nnd2s1 \IDinst/U6975  ( .DIN1(\IDinst/n6955 ), .DIN2(\IDinst/n6954 ), 
        .Q(\IDinst/n6956 ) );
  nnd2s1 \IDinst/U6974  ( .DIN1(\IDinst/n6953 ), .DIN2(n644), 
        .Q(\IDinst/n6955 ) );
  nnd2s1 \IDinst/U6973  ( .DIN1(\IDinst/n6932 ), .DIN2(n672), 
        .Q(\IDinst/n6954 ) );
  nnd2s1 \IDinst/U6972  ( .DIN1(\IDinst/n6952 ), .DIN2(\IDinst/n6951 ), 
        .Q(\IDinst/n6953 ) );
  nnd2s1 \IDinst/U6971  ( .DIN1(\IDinst/n6950 ), .DIN2(n1191), 
        .Q(\IDinst/n6952 ) );
  nnd2s1 \IDinst/U6970  ( .DIN1(\IDinst/n6941 ), .DIN2(n1183), 
        .Q(\IDinst/n6951 ) );
  nnd2s1 \IDinst/U6969  ( .DIN1(\IDinst/n6949 ), .DIN2(\IDinst/n6948 ), 
        .Q(\IDinst/n6950 ) );
  nnd2s1 \IDinst/U6968  ( .DIN1(\IDinst/n6947 ), .DIN2(n1174), 
        .Q(\IDinst/n6949 ) );
  nnd2s1 \IDinst/U6967  ( .DIN1(\IDinst/n6944 ), .DIN2(n1137), 
        .Q(\IDinst/n6948 ) );
  nnd2s1 \IDinst/U6966  ( .DIN1(\IDinst/n6946 ), .DIN2(\IDinst/n6945 ), 
        .Q(\IDinst/n6947 ) );
  nnd2s1 \IDinst/U6965  ( .DIN1(\IDinst/RegFile[15][10] ), .DIN2(n1121), 
        .Q(\IDinst/n6946 ) );
  nnd2s1 \IDinst/U6964  ( .DIN1(\IDinst/RegFile[14][10] ), .DIN2(n1028), 
        .Q(\IDinst/n6945 ) );
  nnd2s1 \IDinst/U6963  ( .DIN1(\IDinst/n6943 ), .DIN2(\IDinst/n6942 ), 
        .Q(\IDinst/n6944 ) );
  nnd2s1 \IDinst/U6962  ( .DIN1(\IDinst/RegFile[13][10] ), .DIN2(n1121), 
        .Q(\IDinst/n6943 ) );
  nnd2s1 \IDinst/U6961  ( .DIN1(\IDinst/RegFile[12][10] ), .DIN2(n1028), 
        .Q(\IDinst/n6942 ) );
  nnd2s1 \IDinst/U6960  ( .DIN1(\IDinst/n6940 ), .DIN2(\IDinst/n6939 ), 
        .Q(\IDinst/n6941 ) );
  nnd2s1 \IDinst/U6959  ( .DIN1(\IDinst/n6938 ), .DIN2(n1174), 
        .Q(\IDinst/n6940 ) );
  nnd2s1 \IDinst/U6958  ( .DIN1(\IDinst/n6935 ), .DIN2(n1137), 
        .Q(\IDinst/n6939 ) );
  nnd2s1 \IDinst/U6957  ( .DIN1(\IDinst/n6937 ), .DIN2(\IDinst/n6936 ), 
        .Q(\IDinst/n6938 ) );
  nnd2s1 \IDinst/U6956  ( .DIN1(\IDinst/RegFile[11][10] ), .DIN2(n1121), 
        .Q(\IDinst/n6937 ) );
  nnd2s1 \IDinst/U6955  ( .DIN1(\IDinst/RegFile[10][10] ), .DIN2(n1028), 
        .Q(\IDinst/n6936 ) );
  nnd2s1 \IDinst/U6954  ( .DIN1(\IDinst/n6934 ), .DIN2(\IDinst/n6933 ), 
        .Q(\IDinst/n6935 ) );
  nnd2s1 \IDinst/U6953  ( .DIN1(\IDinst/RegFile[9][10] ), .DIN2(n1121), 
        .Q(\IDinst/n6934 ) );
  nnd2s1 \IDinst/U6952  ( .DIN1(\IDinst/RegFile[8][10] ), .DIN2(n1028), 
        .Q(\IDinst/n6933 ) );
  nnd2s1 \IDinst/U6951  ( .DIN1(\IDinst/n6931 ), .DIN2(\IDinst/n6930 ), 
        .Q(\IDinst/n6932 ) );
  nnd2s1 \IDinst/U6950  ( .DIN1(\IDinst/n6929 ), .DIN2(n1195), 
        .Q(\IDinst/n6931 ) );
  nnd2s1 \IDinst/U6949  ( .DIN1(\IDinst/n6920 ), .DIN2(n1183), 
        .Q(\IDinst/n6930 ) );
  nnd2s1 \IDinst/U6948  ( .DIN1(\IDinst/n6928 ), .DIN2(\IDinst/n6927 ), 
        .Q(\IDinst/n6929 ) );
  nnd2s1 \IDinst/U6947  ( .DIN1(\IDinst/n6926 ), .DIN2(n1174), 
        .Q(\IDinst/n6928 ) );
  nnd2s1 \IDinst/U6946  ( .DIN1(\IDinst/n6923 ), .DIN2(n1137), 
        .Q(\IDinst/n6927 ) );
  nnd2s1 \IDinst/U6945  ( .DIN1(\IDinst/n6925 ), .DIN2(\IDinst/n6924 ), 
        .Q(\IDinst/n6926 ) );
  nnd2s1 \IDinst/U6944  ( .DIN1(\IDinst/RegFile[7][10] ), .DIN2(n1121), 
        .Q(\IDinst/n6925 ) );
  nnd2s1 \IDinst/U6943  ( .DIN1(\IDinst/RegFile[6][10] ), .DIN2(n1028), 
        .Q(\IDinst/n6924 ) );
  nnd2s1 \IDinst/U6942  ( .DIN1(\IDinst/n6922 ), .DIN2(\IDinst/n6921 ), 
        .Q(\IDinst/n6923 ) );
  nnd2s1 \IDinst/U6941  ( .DIN1(\IDinst/RegFile[5][10] ), .DIN2(n1121), 
        .Q(\IDinst/n6922 ) );
  nnd2s1 \IDinst/U6940  ( .DIN1(\IDinst/RegFile[4][10] ), .DIN2(n1028), 
        .Q(\IDinst/n6921 ) );
  nnd2s1 \IDinst/U6939  ( .DIN1(\IDinst/n6919 ), .DIN2(\IDinst/n6918 ), 
        .Q(\IDinst/n6920 ) );
  nnd2s1 \IDinst/U6938  ( .DIN1(\IDinst/n6917 ), .DIN2(n1174), 
        .Q(\IDinst/n6919 ) );
  nnd2s1 \IDinst/U6937  ( .DIN1(\IDinst/n6914 ), .DIN2(n1137), 
        .Q(\IDinst/n6918 ) );
  nnd2s1 \IDinst/U6936  ( .DIN1(\IDinst/n6916 ), .DIN2(\IDinst/n6915 ), 
        .Q(\IDinst/n6917 ) );
  nnd2s1 \IDinst/U6935  ( .DIN1(\IDinst/RegFile[3][10] ), .DIN2(n1121), 
        .Q(\IDinst/n6916 ) );
  nnd2s1 \IDinst/U6934  ( .DIN1(\IDinst/RegFile[2][10] ), .DIN2(n1028), 
        .Q(\IDinst/n6915 ) );
  nnd2s1 \IDinst/U6933  ( .DIN1(\IDinst/n6913 ), .DIN2(\IDinst/n6912 ), 
        .Q(\IDinst/n6914 ) );
  nnd2s1 \IDinst/U6932  ( .DIN1(\IDinst/RegFile[1][10] ), .DIN2(n1120), 
        .Q(\IDinst/n6913 ) );
  nnd2s1 \IDinst/U6931  ( .DIN1(\IDinst/RegFile[0][10] ), .DIN2(n1028), 
        .Q(\IDinst/n6912 ) );
  nnd2s1 \IDinst/U6930  ( .DIN1(\IDinst/n6911 ), .DIN2(n539), 
        .Q(\IDinst/n5966 ) );
  nnd2s1 \IDinst/U6929  ( .DIN1(\IDinst/n6866 ), .DIN2(n635), 
        .Q(\IDinst/n5967 ) );
  nnd2s1 \IDinst/U6928  ( .DIN1(\IDinst/n6910 ), .DIN2(\IDinst/n6909 ), 
        .Q(\IDinst/n6911 ) );
  nnd2s1 \IDinst/U6927  ( .DIN1(\IDinst/n6908 ), .DIN2(n643), 
        .Q(\IDinst/n6910 ) );
  nnd2s1 \IDinst/U6926  ( .DIN1(\IDinst/n6887 ), .DIN2(n670), 
        .Q(\IDinst/n6909 ) );
  nnd2s1 \IDinst/U6925  ( .DIN1(\IDinst/n6907 ), .DIN2(\IDinst/n6906 ), 
        .Q(\IDinst/n6908 ) );
  nnd2s1 \IDinst/U6924  ( .DIN1(\IDinst/n6905 ), .DIN2(n1193), 
        .Q(\IDinst/n6907 ) );
  nnd2s1 \IDinst/U6923  ( .DIN1(\IDinst/n6896 ), .DIN2(n1183), 
        .Q(\IDinst/n6906 ) );
  nnd2s1 \IDinst/U6922  ( .DIN1(\IDinst/n6904 ), .DIN2(\IDinst/n6903 ), 
        .Q(\IDinst/n6905 ) );
  nnd2s1 \IDinst/U6921  ( .DIN1(\IDinst/n6902 ), .DIN2(n1174), 
        .Q(\IDinst/n6904 ) );
  nnd2s1 \IDinst/U6920  ( .DIN1(\IDinst/n6899 ), .DIN2(n1137), 
        .Q(\IDinst/n6903 ) );
  nnd2s1 \IDinst/U6919  ( .DIN1(\IDinst/n6901 ), .DIN2(\IDinst/n6900 ), 
        .Q(\IDinst/n6902 ) );
  nnd2s1 \IDinst/U6918  ( .DIN1(\IDinst/RegFile[31][9] ), .DIN2(n1120), 
        .Q(\IDinst/n6901 ) );
  nnd2s1 \IDinst/U6917  ( .DIN1(\IDinst/RegFile[30][9] ), .DIN2(n1028), 
        .Q(\IDinst/n6900 ) );
  nnd2s1 \IDinst/U6916  ( .DIN1(\IDinst/n6898 ), .DIN2(\IDinst/n6897 ), 
        .Q(\IDinst/n6899 ) );
  nnd2s1 \IDinst/U6915  ( .DIN1(\IDinst/RegFile[29][9] ), .DIN2(n1120), 
        .Q(\IDinst/n6898 ) );
  nnd2s1 \IDinst/U6914  ( .DIN1(\IDinst/RegFile[28][9] ), .DIN2(n1027), 
        .Q(\IDinst/n6897 ) );
  nnd2s1 \IDinst/U6913  ( .DIN1(\IDinst/n6895 ), .DIN2(\IDinst/n6894 ), 
        .Q(\IDinst/n6896 ) );
  nnd2s1 \IDinst/U6912  ( .DIN1(\IDinst/n6893 ), .DIN2(n1173), 
        .Q(\IDinst/n6895 ) );
  nnd2s1 \IDinst/U6911  ( .DIN1(\IDinst/n6890 ), .DIN2(n1137), 
        .Q(\IDinst/n6894 ) );
  nnd2s1 \IDinst/U6910  ( .DIN1(\IDinst/n6892 ), .DIN2(\IDinst/n6891 ), 
        .Q(\IDinst/n6893 ) );
  nnd2s1 \IDinst/U6909  ( .DIN1(\IDinst/RegFile[27][9] ), .DIN2(n1120), 
        .Q(\IDinst/n6892 ) );
  nnd2s1 \IDinst/U6908  ( .DIN1(\IDinst/RegFile[26][9] ), .DIN2(n1027), 
        .Q(\IDinst/n6891 ) );
  nnd2s1 \IDinst/U6907  ( .DIN1(\IDinst/n6889 ), .DIN2(\IDinst/n6888 ), 
        .Q(\IDinst/n6890 ) );
  nnd2s1 \IDinst/U6906  ( .DIN1(\IDinst/RegFile[25][9] ), .DIN2(n1120), 
        .Q(\IDinst/n6889 ) );
  nnd2s1 \IDinst/U6905  ( .DIN1(\IDinst/RegFile[24][9] ), .DIN2(n1027), 
        .Q(\IDinst/n6888 ) );
  nnd2s1 \IDinst/U6904  ( .DIN1(\IDinst/n6886 ), .DIN2(\IDinst/n6885 ), 
        .Q(\IDinst/n6887 ) );
  nnd2s1 \IDinst/U6903  ( .DIN1(\IDinst/n6884 ), .DIN2(n1192), 
        .Q(\IDinst/n6886 ) );
  nnd2s1 \IDinst/U6902  ( .DIN1(\IDinst/n6875 ), .DIN2(n1183), 
        .Q(\IDinst/n6885 ) );
  nnd2s1 \IDinst/U6901  ( .DIN1(\IDinst/n6883 ), .DIN2(\IDinst/n6882 ), 
        .Q(\IDinst/n6884 ) );
  nnd2s1 \IDinst/U6900  ( .DIN1(\IDinst/n6881 ), .DIN2(n1173), 
        .Q(\IDinst/n6883 ) );
  nnd2s1 \IDinst/U6899  ( .DIN1(\IDinst/n6878 ), .DIN2(n1137), 
        .Q(\IDinst/n6882 ) );
  nnd2s1 \IDinst/U6898  ( .DIN1(\IDinst/n6880 ), .DIN2(\IDinst/n6879 ), 
        .Q(\IDinst/n6881 ) );
  nnd2s1 \IDinst/U6897  ( .DIN1(\IDinst/RegFile[23][9] ), .DIN2(n1120), 
        .Q(\IDinst/n6880 ) );
  nnd2s1 \IDinst/U6896  ( .DIN1(\IDinst/RegFile[22][9] ), .DIN2(n1027), 
        .Q(\IDinst/n6879 ) );
  nnd2s1 \IDinst/U6895  ( .DIN1(\IDinst/n6877 ), .DIN2(\IDinst/n6876 ), 
        .Q(\IDinst/n6878 ) );
  nnd2s1 \IDinst/U6894  ( .DIN1(\IDinst/RegFile[21][9] ), .DIN2(n1120), 
        .Q(\IDinst/n6877 ) );
  nnd2s1 \IDinst/U6893  ( .DIN1(\IDinst/RegFile[20][9] ), .DIN2(n1027), 
        .Q(\IDinst/n6876 ) );
  nnd2s1 \IDinst/U6892  ( .DIN1(\IDinst/n6874 ), .DIN2(\IDinst/n6873 ), 
        .Q(\IDinst/n6875 ) );
  nnd2s1 \IDinst/U6891  ( .DIN1(\IDinst/n6872 ), .DIN2(n1173), 
        .Q(\IDinst/n6874 ) );
  nnd2s1 \IDinst/U6890  ( .DIN1(\IDinst/n6869 ), .DIN2(n1137), 
        .Q(\IDinst/n6873 ) );
  nnd2s1 \IDinst/U6889  ( .DIN1(\IDinst/n6871 ), .DIN2(\IDinst/n6870 ), 
        .Q(\IDinst/n6872 ) );
  nnd2s1 \IDinst/U6888  ( .DIN1(\IDinst/RegFile[19][9] ), .DIN2(n1120), 
        .Q(\IDinst/n6871 ) );
  nnd2s1 \IDinst/U6887  ( .DIN1(\IDinst/RegFile[18][9] ), .DIN2(n1027), 
        .Q(\IDinst/n6870 ) );
  nnd2s1 \IDinst/U6886  ( .DIN1(\IDinst/n6868 ), .DIN2(\IDinst/n6867 ), 
        .Q(\IDinst/n6869 ) );
  nnd2s1 \IDinst/U6885  ( .DIN1(\IDinst/RegFile[17][9] ), .DIN2(n1120), 
        .Q(\IDinst/n6868 ) );
  nnd2s1 \IDinst/U6884  ( .DIN1(\IDinst/RegFile[16][9] ), .DIN2(n1027), 
        .Q(\IDinst/n6867 ) );
  nnd2s1 \IDinst/U6883  ( .DIN1(\IDinst/n6865 ), .DIN2(\IDinst/n6864 ), 
        .Q(\IDinst/n6866 ) );
  nnd2s1 \IDinst/U6882  ( .DIN1(\IDinst/n6863 ), .DIN2(n642), 
        .Q(\IDinst/n6865 ) );
  nnd2s1 \IDinst/U6881  ( .DIN1(\IDinst/n6842 ), .DIN2(n673), 
        .Q(\IDinst/n6864 ) );
  nnd2s1 \IDinst/U6880  ( .DIN1(\IDinst/n6862 ), .DIN2(\IDinst/n6861 ), 
        .Q(\IDinst/n6863 ) );
  nnd2s1 \IDinst/U6879  ( .DIN1(\IDinst/n6860 ), .DIN2(n1192), 
        .Q(\IDinst/n6862 ) );
  nnd2s1 \IDinst/U6878  ( .DIN1(\IDinst/n6851 ), .DIN2(n1183), 
        .Q(\IDinst/n6861 ) );
  nnd2s1 \IDinst/U6877  ( .DIN1(\IDinst/n6859 ), .DIN2(\IDinst/n6858 ), 
        .Q(\IDinst/n6860 ) );
  nnd2s1 \IDinst/U6876  ( .DIN1(\IDinst/n6857 ), .DIN2(n1173), 
        .Q(\IDinst/n6859 ) );
  nnd2s1 \IDinst/U6875  ( .DIN1(\IDinst/n6854 ), .DIN2(n1137), 
        .Q(\IDinst/n6858 ) );
  nnd2s1 \IDinst/U6874  ( .DIN1(\IDinst/n6856 ), .DIN2(\IDinst/n6855 ), 
        .Q(\IDinst/n6857 ) );
  nnd2s1 \IDinst/U6873  ( .DIN1(\IDinst/RegFile[15][9] ), .DIN2(n1119), 
        .Q(\IDinst/n6856 ) );
  nnd2s1 \IDinst/U6872  ( .DIN1(\IDinst/RegFile[14][9] ), .DIN2(n1027), 
        .Q(\IDinst/n6855 ) );
  nnd2s1 \IDinst/U6871  ( .DIN1(\IDinst/n6853 ), .DIN2(\IDinst/n6852 ), 
        .Q(\IDinst/n6854 ) );
  nnd2s1 \IDinst/U6870  ( .DIN1(\IDinst/RegFile[13][9] ), .DIN2(n1119), 
        .Q(\IDinst/n6853 ) );
  nnd2s1 \IDinst/U6869  ( .DIN1(\IDinst/RegFile[12][9] ), .DIN2(n1027), 
        .Q(\IDinst/n6852 ) );
  nnd2s1 \IDinst/U6868  ( .DIN1(\IDinst/n6850 ), .DIN2(\IDinst/n6849 ), 
        .Q(\IDinst/n6851 ) );
  nnd2s1 \IDinst/U6867  ( .DIN1(\IDinst/n6848 ), .DIN2(n1173), 
        .Q(\IDinst/n6850 ) );
  nnd2s1 \IDinst/U6866  ( .DIN1(\IDinst/n6845 ), .DIN2(n1137), 
        .Q(\IDinst/n6849 ) );
  nnd2s1 \IDinst/U6865  ( .DIN1(\IDinst/n6847 ), .DIN2(\IDinst/n6846 ), 
        .Q(\IDinst/n6848 ) );
  nnd2s1 \IDinst/U6864  ( .DIN1(\IDinst/RegFile[11][9] ), .DIN2(n1119), 
        .Q(\IDinst/n6847 ) );
  nnd2s1 \IDinst/U6863  ( .DIN1(\IDinst/RegFile[10][9] ), .DIN2(n1027), 
        .Q(\IDinst/n6846 ) );
  nnd2s1 \IDinst/U6862  ( .DIN1(\IDinst/n6844 ), .DIN2(\IDinst/n6843 ), 
        .Q(\IDinst/n6845 ) );
  nnd2s1 \IDinst/U6861  ( .DIN1(\IDinst/RegFile[9][9] ), .DIN2(n1119), 
        .Q(\IDinst/n6844 ) );
  nnd2s1 \IDinst/U6860  ( .DIN1(\IDinst/RegFile[8][9] ), .DIN2(n1027), 
        .Q(\IDinst/n6843 ) );
  nnd2s1 \IDinst/U6859  ( .DIN1(\IDinst/n6841 ), .DIN2(\IDinst/n6840 ), 
        .Q(\IDinst/n6842 ) );
  nnd2s1 \IDinst/U6858  ( .DIN1(\IDinst/n6839 ), .DIN2(n1194), 
        .Q(\IDinst/n6841 ) );
  nnd2s1 \IDinst/U6857  ( .DIN1(\IDinst/n6830 ), .DIN2(n1183), 
        .Q(\IDinst/n6840 ) );
  nnd2s1 \IDinst/U6856  ( .DIN1(\IDinst/n6838 ), .DIN2(\IDinst/n6837 ), 
        .Q(\IDinst/n6839 ) );
  nnd2s1 \IDinst/U6855  ( .DIN1(\IDinst/n6836 ), .DIN2(n1173), 
        .Q(\IDinst/n6838 ) );
  nnd2s1 \IDinst/U6854  ( .DIN1(\IDinst/n6833 ), .DIN2(n1137), 
        .Q(\IDinst/n6837 ) );
  nnd2s1 \IDinst/U6853  ( .DIN1(\IDinst/n6835 ), .DIN2(\IDinst/n6834 ), 
        .Q(\IDinst/n6836 ) );
  nnd2s1 \IDinst/U6852  ( .DIN1(\IDinst/RegFile[7][9] ), .DIN2(n1119), 
        .Q(\IDinst/n6835 ) );
  nnd2s1 \IDinst/U6851  ( .DIN1(\IDinst/RegFile[6][9] ), .DIN2(n1027), 
        .Q(\IDinst/n6834 ) );
  nnd2s1 \IDinst/U6850  ( .DIN1(\IDinst/n6832 ), .DIN2(\IDinst/n6831 ), 
        .Q(\IDinst/n6833 ) );
  nnd2s1 \IDinst/U6849  ( .DIN1(\IDinst/RegFile[5][9] ), .DIN2(n1119), 
        .Q(\IDinst/n6832 ) );
  nnd2s1 \IDinst/U6848  ( .DIN1(\IDinst/RegFile[4][9] ), .DIN2(n1027), 
        .Q(\IDinst/n6831 ) );
  nnd2s1 \IDinst/U6847  ( .DIN1(\IDinst/n6829 ), .DIN2(\IDinst/n6828 ), 
        .Q(\IDinst/n6830 ) );
  nnd2s1 \IDinst/U6846  ( .DIN1(\IDinst/n6827 ), .DIN2(n1173), 
        .Q(\IDinst/n6829 ) );
  nnd2s1 \IDinst/U6845  ( .DIN1(\IDinst/n6824 ), .DIN2(n1138), 
        .Q(\IDinst/n6828 ) );
  nnd2s1 \IDinst/U6844  ( .DIN1(\IDinst/n6826 ), .DIN2(\IDinst/n6825 ), 
        .Q(\IDinst/n6827 ) );
  nnd2s1 \IDinst/U6843  ( .DIN1(\IDinst/RegFile[3][9] ), .DIN2(n1119), 
        .Q(\IDinst/n6826 ) );
  nnd2s1 \IDinst/U6842  ( .DIN1(\IDinst/RegFile[2][9] ), .DIN2(n1026), 
        .Q(\IDinst/n6825 ) );
  nnd2s1 \IDinst/U6841  ( .DIN1(\IDinst/n6823 ), .DIN2(\IDinst/n6822 ), 
        .Q(\IDinst/n6824 ) );
  nnd2s1 \IDinst/U6840  ( .DIN1(\IDinst/RegFile[1][9] ), .DIN2(n1119), 
        .Q(\IDinst/n6823 ) );
  nnd2s1 \IDinst/U6839  ( .DIN1(\IDinst/RegFile[0][9] ), .DIN2(n1026), 
        .Q(\IDinst/n6822 ) );
  nnd2s1 \IDinst/U6838  ( .DIN1(\IDinst/n6821 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n5964 ) );
  nnd2s1 \IDinst/U6837  ( .DIN1(\IDinst/n6776 ), .DIN2(n636), 
        .Q(\IDinst/n5965 ) );
  nnd2s1 \IDinst/U6836  ( .DIN1(\IDinst/n6820 ), .DIN2(\IDinst/n6819 ), 
        .Q(\IDinst/n6821 ) );
  nnd2s1 \IDinst/U6835  ( .DIN1(\IDinst/n6818 ), .DIN2(n641), 
        .Q(\IDinst/n6820 ) );
  nnd2s1 \IDinst/U6834  ( .DIN1(\IDinst/n6797 ), .DIN2(n671), 
        .Q(\IDinst/n6819 ) );
  nnd2s1 \IDinst/U6833  ( .DIN1(\IDinst/n6817 ), .DIN2(\IDinst/n6816 ), 
        .Q(\IDinst/n6818 ) );
  nnd2s1 \IDinst/U6832  ( .DIN1(\IDinst/n6815 ), .DIN2(n1194), 
        .Q(\IDinst/n6817 ) );
  nnd2s1 \IDinst/U6831  ( .DIN1(\IDinst/n6806 ), .DIN2(n1183), 
        .Q(\IDinst/n6816 ) );
  nnd2s1 \IDinst/U6830  ( .DIN1(\IDinst/n6814 ), .DIN2(\IDinst/n6813 ), 
        .Q(\IDinst/n6815 ) );
  nnd2s1 \IDinst/U6829  ( .DIN1(\IDinst/n6812 ), .DIN2(n1173), 
        .Q(\IDinst/n6814 ) );
  nnd2s1 \IDinst/U6828  ( .DIN1(\IDinst/n6809 ), .DIN2(n1138), 
        .Q(\IDinst/n6813 ) );
  nnd2s1 \IDinst/U6827  ( .DIN1(\IDinst/n6811 ), .DIN2(\IDinst/n6810 ), 
        .Q(\IDinst/n6812 ) );
  nnd2s1 \IDinst/U6826  ( .DIN1(\IDinst/RegFile[31][8] ), .DIN2(n1118), 
        .Q(\IDinst/n6811 ) );
  nnd2s1 \IDinst/U6825  ( .DIN1(\IDinst/RegFile[30][8] ), .DIN2(n1026), 
        .Q(\IDinst/n6810 ) );
  nnd2s1 \IDinst/U6824  ( .DIN1(\IDinst/n6808 ), .DIN2(\IDinst/n6807 ), 
        .Q(\IDinst/n6809 ) );
  nnd2s1 \IDinst/U6823  ( .DIN1(\IDinst/RegFile[29][8] ), .DIN2(n1118), 
        .Q(\IDinst/n6808 ) );
  nnd2s1 \IDinst/U6822  ( .DIN1(\IDinst/RegFile[28][8] ), .DIN2(n1026), 
        .Q(\IDinst/n6807 ) );
  nnd2s1 \IDinst/U6821  ( .DIN1(\IDinst/n6805 ), .DIN2(\IDinst/n6804 ), 
        .Q(\IDinst/n6806 ) );
  nnd2s1 \IDinst/U6820  ( .DIN1(\IDinst/n6803 ), .DIN2(n1173), 
        .Q(\IDinst/n6805 ) );
  nnd2s1 \IDinst/U6819  ( .DIN1(\IDinst/n6800 ), .DIN2(n1138), 
        .Q(\IDinst/n6804 ) );
  nnd2s1 \IDinst/U6818  ( .DIN1(\IDinst/n6802 ), .DIN2(\IDinst/n6801 ), 
        .Q(\IDinst/n6803 ) );
  nnd2s1 \IDinst/U6817  ( .DIN1(\IDinst/RegFile[27][8] ), .DIN2(n1118), 
        .Q(\IDinst/n6802 ) );
  nnd2s1 \IDinst/U6816  ( .DIN1(\IDinst/RegFile[26][8] ), .DIN2(n1026), 
        .Q(\IDinst/n6801 ) );
  nnd2s1 \IDinst/U6815  ( .DIN1(\IDinst/n6799 ), .DIN2(\IDinst/n6798 ), 
        .Q(\IDinst/n6800 ) );
  nnd2s1 \IDinst/U6814  ( .DIN1(\IDinst/RegFile[25][8] ), .DIN2(n1118), 
        .Q(\IDinst/n6799 ) );
  nnd2s1 \IDinst/U6813  ( .DIN1(\IDinst/RegFile[24][8] ), .DIN2(n1026), 
        .Q(\IDinst/n6798 ) );
  nnd2s1 \IDinst/U6812  ( .DIN1(\IDinst/n6796 ), .DIN2(\IDinst/n6795 ), 
        .Q(\IDinst/n6797 ) );
  nnd2s1 \IDinst/U6811  ( .DIN1(\IDinst/n6794 ), .DIN2(n1194), 
        .Q(\IDinst/n6796 ) );
  nnd2s1 \IDinst/U6810  ( .DIN1(\IDinst/n6785 ), .DIN2(n1183), 
        .Q(\IDinst/n6795 ) );
  nnd2s1 \IDinst/U6809  ( .DIN1(\IDinst/n6793 ), .DIN2(\IDinst/n6792 ), 
        .Q(\IDinst/n6794 ) );
  nnd2s1 \IDinst/U6808  ( .DIN1(\IDinst/n6791 ), .DIN2(n1172), 
        .Q(\IDinst/n6793 ) );
  nnd2s1 \IDinst/U6807  ( .DIN1(\IDinst/n6788 ), .DIN2(n1138), 
        .Q(\IDinst/n6792 ) );
  nnd2s1 \IDinst/U6806  ( .DIN1(\IDinst/n6790 ), .DIN2(\IDinst/n6789 ), 
        .Q(\IDinst/n6791 ) );
  nnd2s1 \IDinst/U6805  ( .DIN1(\IDinst/RegFile[23][8] ), .DIN2(n1118), 
        .Q(\IDinst/n6790 ) );
  nnd2s1 \IDinst/U6804  ( .DIN1(\IDinst/RegFile[22][8] ), .DIN2(n1026), 
        .Q(\IDinst/n6789 ) );
  nnd2s1 \IDinst/U6803  ( .DIN1(\IDinst/n6787 ), .DIN2(\IDinst/n6786 ), 
        .Q(\IDinst/n6788 ) );
  nnd2s1 \IDinst/U6802  ( .DIN1(\IDinst/RegFile[21][8] ), .DIN2(n1118), 
        .Q(\IDinst/n6787 ) );
  nnd2s1 \IDinst/U6801  ( .DIN1(\IDinst/RegFile[20][8] ), .DIN2(n1026), 
        .Q(\IDinst/n6786 ) );
  nnd2s1 \IDinst/U6800  ( .DIN1(\IDinst/n6784 ), .DIN2(\IDinst/n6783 ), 
        .Q(\IDinst/n6785 ) );
  nnd2s1 \IDinst/U6799  ( .DIN1(\IDinst/n6782 ), .DIN2(n1172), 
        .Q(\IDinst/n6784 ) );
  nnd2s1 \IDinst/U6798  ( .DIN1(\IDinst/n6779 ), .DIN2(n1138), 
        .Q(\IDinst/n6783 ) );
  nnd2s1 \IDinst/U6797  ( .DIN1(\IDinst/n6781 ), .DIN2(\IDinst/n6780 ), 
        .Q(\IDinst/n6782 ) );
  nnd2s1 \IDinst/U6796  ( .DIN1(\IDinst/RegFile[19][8] ), .DIN2(n1118), 
        .Q(\IDinst/n6781 ) );
  nnd2s1 \IDinst/U6795  ( .DIN1(\IDinst/RegFile[18][8] ), .DIN2(n1026), 
        .Q(\IDinst/n6780 ) );
  nnd2s1 \IDinst/U6794  ( .DIN1(\IDinst/n6778 ), .DIN2(\IDinst/n6777 ), 
        .Q(\IDinst/n6779 ) );
  nnd2s1 \IDinst/U6793  ( .DIN1(\IDinst/RegFile[17][8] ), .DIN2(n1118), 
        .Q(\IDinst/n6778 ) );
  nnd2s1 \IDinst/U6792  ( .DIN1(\IDinst/RegFile[16][8] ), .DIN2(n1026), 
        .Q(\IDinst/n6777 ) );
  nnd2s1 \IDinst/U6791  ( .DIN1(\IDinst/n6775 ), .DIN2(\IDinst/n6774 ), 
        .Q(\IDinst/n6776 ) );
  nnd2s1 \IDinst/U6790  ( .DIN1(\IDinst/n6773 ), .DIN2(n644), 
        .Q(\IDinst/n6775 ) );
  nnd2s1 \IDinst/U6789  ( .DIN1(\IDinst/n6752 ), .DIN2(n672), 
        .Q(\IDinst/n6774 ) );
  nnd2s1 \IDinst/U6788  ( .DIN1(\IDinst/n6772 ), .DIN2(\IDinst/n6771 ), 
        .Q(\IDinst/n6773 ) );
  nnd2s1 \IDinst/U6787  ( .DIN1(\IDinst/n6770 ), .DIN2(n1194), 
        .Q(\IDinst/n6772 ) );
  nnd2s1 \IDinst/U6786  ( .DIN1(\IDinst/n6761 ), .DIN2(n1183), 
        .Q(\IDinst/n6771 ) );
  nnd2s1 \IDinst/U6785  ( .DIN1(\IDinst/n6769 ), .DIN2(\IDinst/n6768 ), 
        .Q(\IDinst/n6770 ) );
  nnd2s1 \IDinst/U6784  ( .DIN1(\IDinst/n6767 ), .DIN2(n1172), 
        .Q(\IDinst/n6769 ) );
  nnd2s1 \IDinst/U6783  ( .DIN1(\IDinst/n6764 ), .DIN2(n1138), 
        .Q(\IDinst/n6768 ) );
  nnd2s1 \IDinst/U6782  ( .DIN1(\IDinst/n6766 ), .DIN2(\IDinst/n6765 ), 
        .Q(\IDinst/n6767 ) );
  nnd2s1 \IDinst/U6781  ( .DIN1(\IDinst/RegFile[15][8] ), .DIN2(n1118), 
        .Q(\IDinst/n6766 ) );
  nnd2s1 \IDinst/U6780  ( .DIN1(\IDinst/RegFile[14][8] ), .DIN2(n1026), 
        .Q(\IDinst/n6765 ) );
  nnd2s1 \IDinst/U6779  ( .DIN1(\IDinst/n6763 ), .DIN2(\IDinst/n6762 ), 
        .Q(\IDinst/n6764 ) );
  nnd2s1 \IDinst/U6778  ( .DIN1(\IDinst/RegFile[13][8] ), .DIN2(n1117), 
        .Q(\IDinst/n6763 ) );
  nnd2s1 \IDinst/U6777  ( .DIN1(\IDinst/RegFile[12][8] ), .DIN2(n1026), 
        .Q(\IDinst/n6762 ) );
  nnd2s1 \IDinst/U6776  ( .DIN1(\IDinst/n6760 ), .DIN2(\IDinst/n6759 ), 
        .Q(\IDinst/n6761 ) );
  nnd2s1 \IDinst/U6775  ( .DIN1(\IDinst/n6758 ), .DIN2(n1172), 
        .Q(\IDinst/n6760 ) );
  nnd2s1 \IDinst/U6774  ( .DIN1(\IDinst/n6755 ), .DIN2(n1138), 
        .Q(\IDinst/n6759 ) );
  nnd2s1 \IDinst/U6773  ( .DIN1(\IDinst/n6757 ), .DIN2(\IDinst/n6756 ), 
        .Q(\IDinst/n6758 ) );
  nnd2s1 \IDinst/U6772  ( .DIN1(\IDinst/RegFile[11][8] ), .DIN2(n1117), 
        .Q(\IDinst/n6757 ) );
  nnd2s1 \IDinst/U6771  ( .DIN1(\IDinst/RegFile[10][8] ), .DIN2(n1026), 
        .Q(\IDinst/n6756 ) );
  nnd2s1 \IDinst/U6770  ( .DIN1(\IDinst/n6754 ), .DIN2(\IDinst/n6753 ), 
        .Q(\IDinst/n6755 ) );
  nnd2s1 \IDinst/U6769  ( .DIN1(\IDinst/RegFile[9][8] ), .DIN2(n1117), 
        .Q(\IDinst/n6754 ) );
  nnd2s1 \IDinst/U6768  ( .DIN1(\IDinst/RegFile[8][8] ), .DIN2(n1025), 
        .Q(\IDinst/n6753 ) );
  nnd2s1 \IDinst/U6767  ( .DIN1(\IDinst/n6751 ), .DIN2(\IDinst/n6750 ), 
        .Q(\IDinst/n6752 ) );
  nnd2s1 \IDinst/U6766  ( .DIN1(\IDinst/n6749 ), .DIN2(n1194), 
        .Q(\IDinst/n6751 ) );
  nnd2s1 \IDinst/U6765  ( .DIN1(\IDinst/n6740 ), .DIN2(n1183), 
        .Q(\IDinst/n6750 ) );
  nnd2s1 \IDinst/U6764  ( .DIN1(\IDinst/n6748 ), .DIN2(\IDinst/n6747 ), 
        .Q(\IDinst/n6749 ) );
  nnd2s1 \IDinst/U6763  ( .DIN1(\IDinst/n6746 ), .DIN2(n1172), 
        .Q(\IDinst/n6748 ) );
  nnd2s1 \IDinst/U6762  ( .DIN1(\IDinst/n6743 ), .DIN2(n1138), 
        .Q(\IDinst/n6747 ) );
  nnd2s1 \IDinst/U6761  ( .DIN1(\IDinst/n6745 ), .DIN2(\IDinst/n6744 ), 
        .Q(\IDinst/n6746 ) );
  nnd2s1 \IDinst/U6760  ( .DIN1(\IDinst/RegFile[7][8] ), .DIN2(n1117), 
        .Q(\IDinst/n6745 ) );
  nnd2s1 \IDinst/U6759  ( .DIN1(\IDinst/RegFile[6][8] ), .DIN2(n1025), 
        .Q(\IDinst/n6744 ) );
  nnd2s1 \IDinst/U6758  ( .DIN1(\IDinst/n6742 ), .DIN2(\IDinst/n6741 ), 
        .Q(\IDinst/n6743 ) );
  nnd2s1 \IDinst/U6757  ( .DIN1(\IDinst/RegFile[5][8] ), .DIN2(n1117), 
        .Q(\IDinst/n6742 ) );
  nnd2s1 \IDinst/U6756  ( .DIN1(\IDinst/RegFile[4][8] ), .DIN2(n1025), 
        .Q(\IDinst/n6741 ) );
  nnd2s1 \IDinst/U6755  ( .DIN1(\IDinst/n6739 ), .DIN2(\IDinst/n6738 ), 
        .Q(\IDinst/n6740 ) );
  nnd2s1 \IDinst/U6754  ( .DIN1(\IDinst/n6737 ), .DIN2(n1172), 
        .Q(\IDinst/n6739 ) );
  nnd2s1 \IDinst/U6753  ( .DIN1(\IDinst/n6734 ), .DIN2(n1138), 
        .Q(\IDinst/n6738 ) );
  nnd2s1 \IDinst/U6752  ( .DIN1(\IDinst/n6736 ), .DIN2(\IDinst/n6735 ), 
        .Q(\IDinst/n6737 ) );
  nnd2s1 \IDinst/U6751  ( .DIN1(\IDinst/RegFile[3][8] ), .DIN2(n1117), 
        .Q(\IDinst/n6736 ) );
  nnd2s1 \IDinst/U6750  ( .DIN1(\IDinst/RegFile[2][8] ), .DIN2(n1030), 
        .Q(\IDinst/n6735 ) );
  nnd2s1 \IDinst/U6749  ( .DIN1(\IDinst/n6733 ), .DIN2(\IDinst/n6732 ), 
        .Q(\IDinst/n6734 ) );
  nnd2s1 \IDinst/U6748  ( .DIN1(\IDinst/RegFile[1][8] ), .DIN2(n1117), 
        .Q(\IDinst/n6733 ) );
  nnd2s1 \IDinst/U6747  ( .DIN1(\IDinst/RegFile[0][8] ), .DIN2(n1045), 
        .Q(\IDinst/n6732 ) );
  nnd2s1 \IDinst/U6746  ( .DIN1(\IDinst/n6731 ), .DIN2(n539), 
        .Q(\IDinst/n5962 ) );
  nnd2s1 \IDinst/U6745  ( .DIN1(\IDinst/n6686 ), .DIN2(n635), 
        .Q(\IDinst/n5963 ) );
  nnd2s1 \IDinst/U6744  ( .DIN1(\IDinst/n6730 ), .DIN2(\IDinst/n6729 ), 
        .Q(\IDinst/n6731 ) );
  nnd2s1 \IDinst/U6743  ( .DIN1(\IDinst/n6728 ), .DIN2(n643), 
        .Q(\IDinst/n6730 ) );
  nnd2s1 \IDinst/U6742  ( .DIN1(\IDinst/n6707 ), .DIN2(n670), 
        .Q(\IDinst/n6729 ) );
  nnd2s1 \IDinst/U6741  ( .DIN1(\IDinst/n6727 ), .DIN2(\IDinst/n6726 ), 
        .Q(\IDinst/n6728 ) );
  nnd2s1 \IDinst/U6740  ( .DIN1(\IDinst/n6725 ), .DIN2(n1194), 
        .Q(\IDinst/n6727 ) );
  nnd2s1 \IDinst/U6739  ( .DIN1(\IDinst/n6716 ), .DIN2(n1182), 
        .Q(\IDinst/n6726 ) );
  nnd2s1 \IDinst/U6738  ( .DIN1(\IDinst/n6724 ), .DIN2(\IDinst/n6723 ), 
        .Q(\IDinst/n6725 ) );
  nnd2s1 \IDinst/U6737  ( .DIN1(\IDinst/n6722 ), .DIN2(n1172), 
        .Q(\IDinst/n6724 ) );
  nnd2s1 \IDinst/U6736  ( .DIN1(\IDinst/n6719 ), .DIN2(n1138), 
        .Q(\IDinst/n6723 ) );
  nnd2s1 \IDinst/U6735  ( .DIN1(\IDinst/n6721 ), .DIN2(\IDinst/n6720 ), 
        .Q(\IDinst/n6722 ) );
  nnd2s1 \IDinst/U6734  ( .DIN1(\IDinst/RegFile[31][7] ), .DIN2(n1117), 
        .Q(\IDinst/n6721 ) );
  nnd2s1 \IDinst/U6733  ( .DIN1(\IDinst/RegFile[30][7] ), .DIN2(n1045), 
        .Q(\IDinst/n6720 ) );
  nnd2s1 \IDinst/U6732  ( .DIN1(\IDinst/n6718 ), .DIN2(\IDinst/n6717 ), 
        .Q(\IDinst/n6719 ) );
  nnd2s1 \IDinst/U6731  ( .DIN1(\IDinst/RegFile[29][7] ), .DIN2(n1117), 
        .Q(\IDinst/n6718 ) );
  nnd2s1 \IDinst/U6730  ( .DIN1(\IDinst/RegFile[28][7] ), .DIN2(n1045), 
        .Q(\IDinst/n6717 ) );
  nnd2s1 \IDinst/U6729  ( .DIN1(\IDinst/n6715 ), .DIN2(\IDinst/n6714 ), 
        .Q(\IDinst/n6716 ) );
  nnd2s1 \IDinst/U6728  ( .DIN1(\IDinst/n6713 ), .DIN2(n1172), 
        .Q(\IDinst/n6715 ) );
  nnd2s1 \IDinst/U6727  ( .DIN1(\IDinst/n6710 ), .DIN2(n1138), 
        .Q(\IDinst/n6714 ) );
  nnd2s1 \IDinst/U6726  ( .DIN1(\IDinst/n6712 ), .DIN2(\IDinst/n6711 ), 
        .Q(\IDinst/n6713 ) );
  nnd2s1 \IDinst/U6725  ( .DIN1(\IDinst/RegFile[27][7] ), .DIN2(n1116), 
        .Q(\IDinst/n6712 ) );
  nnd2s1 \IDinst/U6724  ( .DIN1(\IDinst/RegFile[26][7] ), .DIN2(n1045), 
        .Q(\IDinst/n6711 ) );
  nnd2s1 \IDinst/U6723  ( .DIN1(\IDinst/n6709 ), .DIN2(\IDinst/n6708 ), 
        .Q(\IDinst/n6710 ) );
  nnd2s1 \IDinst/U6722  ( .DIN1(\IDinst/RegFile[25][7] ), .DIN2(n1116), 
        .Q(\IDinst/n6709 ) );
  nnd2s1 \IDinst/U6721  ( .DIN1(\IDinst/RegFile[24][7] ), .DIN2(n1045), 
        .Q(\IDinst/n6708 ) );
  nnd2s1 \IDinst/U6720  ( .DIN1(\IDinst/n6706 ), .DIN2(\IDinst/n6705 ), 
        .Q(\IDinst/n6707 ) );
  nnd2s1 \IDinst/U6719  ( .DIN1(\IDinst/n6704 ), .DIN2(n1194), 
        .Q(\IDinst/n6706 ) );
  nnd2s1 \IDinst/U6718  ( .DIN1(\IDinst/n6695 ), .DIN2(n1182), 
        .Q(\IDinst/n6705 ) );
  nnd2s1 \IDinst/U6717  ( .DIN1(\IDinst/n6703 ), .DIN2(\IDinst/n6702 ), 
        .Q(\IDinst/n6704 ) );
  nnd2s1 \IDinst/U6716  ( .DIN1(\IDinst/n6701 ), .DIN2(n1172), 
        .Q(\IDinst/n6703 ) );
  nnd2s1 \IDinst/U6715  ( .DIN1(\IDinst/n6698 ), .DIN2(n1138), 
        .Q(\IDinst/n6702 ) );
  nnd2s1 \IDinst/U6714  ( .DIN1(\IDinst/n6700 ), .DIN2(\IDinst/n6699 ), 
        .Q(\IDinst/n6701 ) );
  nnd2s1 \IDinst/U6713  ( .DIN1(\IDinst/RegFile[23][7] ), .DIN2(n1116), 
        .Q(\IDinst/n6700 ) );
  nnd2s1 \IDinst/U6712  ( .DIN1(\IDinst/RegFile[22][7] ), .DIN2(n1044), 
        .Q(\IDinst/n6699 ) );
  nnd2s1 \IDinst/U6711  ( .DIN1(\IDinst/n6697 ), .DIN2(\IDinst/n6696 ), 
        .Q(\IDinst/n6698 ) );
  nnd2s1 \IDinst/U6710  ( .DIN1(\IDinst/RegFile[21][7] ), .DIN2(n1116), 
        .Q(\IDinst/n6697 ) );
  nnd2s1 \IDinst/U6709  ( .DIN1(\IDinst/RegFile[20][7] ), .DIN2(n1044), 
        .Q(\IDinst/n6696 ) );
  nnd2s1 \IDinst/U6708  ( .DIN1(\IDinst/n6694 ), .DIN2(\IDinst/n6693 ), 
        .Q(\IDinst/n6695 ) );
  nnd2s1 \IDinst/U6707  ( .DIN1(\IDinst/n6692 ), .DIN2(\IDinst/N40 ), 
        .Q(\IDinst/n6694 ) );
  nnd2s1 \IDinst/U6706  ( .DIN1(\IDinst/n6689 ), .DIN2(n1139), 
        .Q(\IDinst/n6693 ) );
  nnd2s1 \IDinst/U6705  ( .DIN1(\IDinst/n6691 ), .DIN2(\IDinst/n6690 ), 
        .Q(\IDinst/n6692 ) );
  nnd2s1 \IDinst/U6704  ( .DIN1(\IDinst/RegFile[19][7] ), .DIN2(n1116), 
        .Q(\IDinst/n6691 ) );
  nnd2s1 \IDinst/U6703  ( .DIN1(\IDinst/RegFile[18][7] ), .DIN2(n1044), 
        .Q(\IDinst/n6690 ) );
  nnd2s1 \IDinst/U6702  ( .DIN1(\IDinst/n6688 ), .DIN2(\IDinst/n6687 ), 
        .Q(\IDinst/n6689 ) );
  nnd2s1 \IDinst/U6701  ( .DIN1(\IDinst/RegFile[17][7] ), .DIN2(n1116), 
        .Q(\IDinst/n6688 ) );
  nnd2s1 \IDinst/U6700  ( .DIN1(\IDinst/RegFile[16][7] ), .DIN2(n1044), 
        .Q(\IDinst/n6687 ) );
  nnd2s1 \IDinst/U6699  ( .DIN1(\IDinst/n6685 ), .DIN2(\IDinst/n6684 ), 
        .Q(\IDinst/n6686 ) );
  nnd2s1 \IDinst/U6698  ( .DIN1(\IDinst/n6683 ), .DIN2(n642), 
        .Q(\IDinst/n6685 ) );
  nnd2s1 \IDinst/U6697  ( .DIN1(\IDinst/n6662 ), .DIN2(n673), 
        .Q(\IDinst/n6684 ) );
  nnd2s1 \IDinst/U6696  ( .DIN1(\IDinst/n6682 ), .DIN2(\IDinst/n6681 ), 
        .Q(\IDinst/n6683 ) );
  nnd2s1 \IDinst/U6695  ( .DIN1(\IDinst/n6680 ), .DIN2(n1194), 
        .Q(\IDinst/n6682 ) );
  nnd2s1 \IDinst/U6694  ( .DIN1(\IDinst/n6671 ), .DIN2(n1182), 
        .Q(\IDinst/n6681 ) );
  nnd2s1 \IDinst/U6693  ( .DIN1(\IDinst/n6679 ), .DIN2(\IDinst/n6678 ), 
        .Q(\IDinst/n6680 ) );
  nnd2s1 \IDinst/U6692  ( .DIN1(\IDinst/n6677 ), .DIN2(\IDinst/N40 ), 
        .Q(\IDinst/n6679 ) );
  nnd2s1 \IDinst/U6691  ( .DIN1(\IDinst/n6674 ), .DIN2(n1139), 
        .Q(\IDinst/n6678 ) );
  nnd2s1 \IDinst/U6690  ( .DIN1(\IDinst/n6676 ), .DIN2(\IDinst/n6675 ), 
        .Q(\IDinst/n6677 ) );
  nnd2s1 \IDinst/U6689  ( .DIN1(\IDinst/RegFile[15][7] ), .DIN2(n1116), 
        .Q(\IDinst/n6676 ) );
  nnd2s1 \IDinst/U6688  ( .DIN1(\IDinst/RegFile[14][7] ), .DIN2(n1044), 
        .Q(\IDinst/n6675 ) );
  nnd2s1 \IDinst/U6687  ( .DIN1(\IDinst/n6673 ), .DIN2(\IDinst/n6672 ), 
        .Q(\IDinst/n6674 ) );
  nnd2s1 \IDinst/U6686  ( .DIN1(\IDinst/RegFile[13][7] ), .DIN2(n1116), 
        .Q(\IDinst/n6673 ) );
  nnd2s1 \IDinst/U6685  ( .DIN1(\IDinst/RegFile[12][7] ), .DIN2(n1044), 
        .Q(\IDinst/n6672 ) );
  nnd2s1 \IDinst/U6684  ( .DIN1(\IDinst/n6670 ), .DIN2(\IDinst/n6669 ), 
        .Q(\IDinst/n6671 ) );
  nnd2s1 \IDinst/U6683  ( .DIN1(\IDinst/n6668 ), .DIN2(\IDinst/N40 ), 
        .Q(\IDinst/n6670 ) );
  nnd2s1 \IDinst/U6682  ( .DIN1(\IDinst/n6665 ), .DIN2(n1139), 
        .Q(\IDinst/n6669 ) );
  nnd2s1 \IDinst/U6681  ( .DIN1(\IDinst/n6667 ), .DIN2(\IDinst/n6666 ), 
        .Q(\IDinst/n6668 ) );
  nnd2s1 \IDinst/U6680  ( .DIN1(\IDinst/RegFile[11][7] ), .DIN2(n1103), 
        .Q(\IDinst/n6667 ) );
  nnd2s1 \IDinst/U6679  ( .DIN1(\IDinst/RegFile[10][7] ), .DIN2(n1044), 
        .Q(\IDinst/n6666 ) );
  nnd2s1 \IDinst/U6678  ( .DIN1(\IDinst/n6664 ), .DIN2(\IDinst/n6663 ), 
        .Q(\IDinst/n6665 ) );
  nnd2s1 \IDinst/U6677  ( .DIN1(\IDinst/RegFile[9][7] ), .DIN2(n1096), 
        .Q(\IDinst/n6664 ) );
  nnd2s1 \IDinst/U6676  ( .DIN1(\IDinst/RegFile[8][7] ), .DIN2(n1044), 
        .Q(\IDinst/n6663 ) );
  nnd2s1 \IDinst/U6675  ( .DIN1(\IDinst/n6661 ), .DIN2(\IDinst/n6660 ), 
        .Q(\IDinst/n6662 ) );
  nnd2s1 \IDinst/U6674  ( .DIN1(\IDinst/n6659 ), .DIN2(n1194), 
        .Q(\IDinst/n6661 ) );
  nnd2s1 \IDinst/U6673  ( .DIN1(\IDinst/n6650 ), .DIN2(n1182), 
        .Q(\IDinst/n6660 ) );
  nnd2s1 \IDinst/U6672  ( .DIN1(\IDinst/n6658 ), .DIN2(\IDinst/n6657 ), 
        .Q(\IDinst/n6659 ) );
  nnd2s1 \IDinst/U6671  ( .DIN1(\IDinst/n6656 ), .DIN2(\IDinst/N40 ), 
        .Q(\IDinst/n6658 ) );
  nnd2s1 \IDinst/U6670  ( .DIN1(\IDinst/n6653 ), .DIN2(n1139), 
        .Q(\IDinst/n6657 ) );
  nnd2s1 \IDinst/U6669  ( .DIN1(\IDinst/n6655 ), .DIN2(\IDinst/n6654 ), 
        .Q(\IDinst/n6656 ) );
  nnd2s1 \IDinst/U6668  ( .DIN1(\IDinst/RegFile[7][7] ), .DIN2(n1096), 
        .Q(\IDinst/n6655 ) );
  nnd2s1 \IDinst/U6667  ( .DIN1(\IDinst/RegFile[6][7] ), .DIN2(n1044), 
        .Q(\IDinst/n6654 ) );
  nnd2s1 \IDinst/U6666  ( .DIN1(\IDinst/n6652 ), .DIN2(\IDinst/n6651 ), 
        .Q(\IDinst/n6653 ) );
  nnd2s1 \IDinst/U6665  ( .DIN1(\IDinst/RegFile[5][7] ), .DIN2(n1096), 
        .Q(\IDinst/n6652 ) );
  nnd2s1 \IDinst/U6664  ( .DIN1(\IDinst/RegFile[4][7] ), .DIN2(n1044), 
        .Q(\IDinst/n6651 ) );
  nnd2s1 \IDinst/U6663  ( .DIN1(\IDinst/n6649 ), .DIN2(\IDinst/n6648 ), 
        .Q(\IDinst/n6650 ) );
  nnd2s1 \IDinst/U6662  ( .DIN1(\IDinst/n6647 ), .DIN2(\IDinst/N40 ), 
        .Q(\IDinst/n6649 ) );
  nnd2s1 \IDinst/U6661  ( .DIN1(\IDinst/n6644 ), .DIN2(n1139), 
        .Q(\IDinst/n6648 ) );
  nnd2s1 \IDinst/U6660  ( .DIN1(\IDinst/n6646 ), .DIN2(\IDinst/n6645 ), 
        .Q(\IDinst/n6647 ) );
  nnd2s1 \IDinst/U6659  ( .DIN1(\IDinst/RegFile[3][7] ), .DIN2(n1096), 
        .Q(\IDinst/n6646 ) );
  nnd2s1 \IDinst/U6658  ( .DIN1(\IDinst/RegFile[2][7] ), .DIN2(n1044), 
        .Q(\IDinst/n6645 ) );
  nnd2s1 \IDinst/U6657  ( .DIN1(\IDinst/n6643 ), .DIN2(\IDinst/n6642 ), 
        .Q(\IDinst/n6644 ) );
  nnd2s1 \IDinst/U6656  ( .DIN1(\IDinst/RegFile[1][7] ), .DIN2(n1097), 
        .Q(\IDinst/n6643 ) );
  nnd2s1 \IDinst/U6655  ( .DIN1(\IDinst/RegFile[0][7] ), .DIN2(n1044), 
        .Q(\IDinst/n6642 ) );
  nnd2s1 \IDinst/U6654  ( .DIN1(\IDinst/n6641 ), .DIN2(n539), 
        .Q(\IDinst/n5960 ) );
  nnd2s1 \IDinst/U6653  ( .DIN1(\IDinst/n6596 ), .DIN2(n636), 
        .Q(\IDinst/n5961 ) );
  nnd2s1 \IDinst/U6652  ( .DIN1(\IDinst/n6640 ), .DIN2(\IDinst/n6639 ), 
        .Q(\IDinst/n6641 ) );
  nnd2s1 \IDinst/U6651  ( .DIN1(\IDinst/n6638 ), .DIN2(n641), 
        .Q(\IDinst/n6640 ) );
  nnd2s1 \IDinst/U6650  ( .DIN1(\IDinst/n6617 ), .DIN2(n671), 
        .Q(\IDinst/n6639 ) );
  nnd2s1 \IDinst/U6649  ( .DIN1(\IDinst/n6637 ), .DIN2(\IDinst/n6636 ), 
        .Q(\IDinst/n6638 ) );
  nnd2s1 \IDinst/U6648  ( .DIN1(\IDinst/n6635 ), .DIN2(n1195), 
        .Q(\IDinst/n6637 ) );
  nnd2s1 \IDinst/U6647  ( .DIN1(\IDinst/n6626 ), .DIN2(n1182), 
        .Q(\IDinst/n6636 ) );
  nnd2s1 \IDinst/U6646  ( .DIN1(\IDinst/n6634 ), .DIN2(\IDinst/n6633 ), 
        .Q(\IDinst/n6635 ) );
  nnd2s1 \IDinst/U6645  ( .DIN1(\IDinst/n6632 ), .DIN2(\IDinst/N40 ), 
        .Q(\IDinst/n6634 ) );
  nnd2s1 \IDinst/U6644  ( .DIN1(\IDinst/n6629 ), .DIN2(n1139), 
        .Q(\IDinst/n6633 ) );
  nnd2s1 \IDinst/U6643  ( .DIN1(\IDinst/n6631 ), .DIN2(\IDinst/n6630 ), 
        .Q(\IDinst/n6632 ) );
  nnd2s1 \IDinst/U6642  ( .DIN1(\IDinst/RegFile[31][6] ), .DIN2(n1097), 
        .Q(\IDinst/n6631 ) );
  nnd2s1 \IDinst/U6641  ( .DIN1(\IDinst/RegFile[30][6] ), .DIN2(n1044), 
        .Q(\IDinst/n6630 ) );
  nnd2s1 \IDinst/U6640  ( .DIN1(\IDinst/n6628 ), .DIN2(\IDinst/n6627 ), 
        .Q(\IDinst/n6629 ) );
  nnd2s1 \IDinst/U6639  ( .DIN1(\IDinst/RegFile[29][6] ), .DIN2(n1097), 
        .Q(\IDinst/n6628 ) );
  nnd2s1 \IDinst/U6638  ( .DIN1(\IDinst/RegFile[28][6] ), .DIN2(n1043), 
        .Q(\IDinst/n6627 ) );
  nnd2s1 \IDinst/U6637  ( .DIN1(\IDinst/n6625 ), .DIN2(\IDinst/n6624 ), 
        .Q(\IDinst/n6626 ) );
  nnd2s1 \IDinst/U6636  ( .DIN1(\IDinst/n6623 ), .DIN2(n1177), 
        .Q(\IDinst/n6625 ) );
  nnd2s1 \IDinst/U6635  ( .DIN1(\IDinst/n6620 ), .DIN2(n1139), 
        .Q(\IDinst/n6624 ) );
  nnd2s1 \IDinst/U6634  ( .DIN1(\IDinst/n6622 ), .DIN2(\IDinst/n6621 ), 
        .Q(\IDinst/n6623 ) );
  nnd2s1 \IDinst/U6633  ( .DIN1(\IDinst/RegFile[27][6] ), .DIN2(n1097), 
        .Q(\IDinst/n6622 ) );
  nnd2s1 \IDinst/U6632  ( .DIN1(\IDinst/RegFile[26][6] ), .DIN2(n1043), 
        .Q(\IDinst/n6621 ) );
  nnd2s1 \IDinst/U6631  ( .DIN1(\IDinst/n6619 ), .DIN2(\IDinst/n6618 ), 
        .Q(\IDinst/n6620 ) );
  nnd2s1 \IDinst/U6630  ( .DIN1(\IDinst/RegFile[25][6] ), .DIN2(n1097), 
        .Q(\IDinst/n6619 ) );
  nnd2s1 \IDinst/U6629  ( .DIN1(\IDinst/RegFile[24][6] ), .DIN2(n1043), 
        .Q(\IDinst/n6618 ) );
  nnd2s1 \IDinst/U6628  ( .DIN1(\IDinst/n6616 ), .DIN2(\IDinst/n6615 ), 
        .Q(\IDinst/n6617 ) );
  nnd2s1 \IDinst/U6627  ( .DIN1(\IDinst/n6614 ), .DIN2(n1195), 
        .Q(\IDinst/n6616 ) );
  nnd2s1 \IDinst/U6626  ( .DIN1(\IDinst/n6605 ), .DIN2(n1182), 
        .Q(\IDinst/n6615 ) );
  nnd2s1 \IDinst/U6625  ( .DIN1(\IDinst/n6613 ), .DIN2(\IDinst/n6612 ), 
        .Q(\IDinst/n6614 ) );
  nnd2s1 \IDinst/U6624  ( .DIN1(\IDinst/n6611 ), .DIN2(n1165), 
        .Q(\IDinst/n6613 ) );
  nnd2s1 \IDinst/U6623  ( .DIN1(\IDinst/n6608 ), .DIN2(n1139), 
        .Q(\IDinst/n6612 ) );
  nnd2s1 \IDinst/U6622  ( .DIN1(\IDinst/n6610 ), .DIN2(\IDinst/n6609 ), 
        .Q(\IDinst/n6611 ) );
  nnd2s1 \IDinst/U6621  ( .DIN1(\IDinst/RegFile[23][6] ), .DIN2(n1097), 
        .Q(\IDinst/n6610 ) );
  nnd2s1 \IDinst/U6620  ( .DIN1(\IDinst/RegFile[22][6] ), .DIN2(n1043), 
        .Q(\IDinst/n6609 ) );
  nnd2s1 \IDinst/U6619  ( .DIN1(\IDinst/n6607 ), .DIN2(\IDinst/n6606 ), 
        .Q(\IDinst/n6608 ) );
  nnd2s1 \IDinst/U6618  ( .DIN1(\IDinst/RegFile[21][6] ), .DIN2(n1097), 
        .Q(\IDinst/n6607 ) );
  nnd2s1 \IDinst/U6617  ( .DIN1(\IDinst/RegFile[20][6] ), .DIN2(n1043), 
        .Q(\IDinst/n6606 ) );
  nnd2s1 \IDinst/U6616  ( .DIN1(\IDinst/n6604 ), .DIN2(\IDinst/n6603 ), 
        .Q(\IDinst/n6605 ) );
  nnd2s1 \IDinst/U6615  ( .DIN1(\IDinst/n6602 ), .DIN2(n1171), 
        .Q(\IDinst/n6604 ) );
  nnd2s1 \IDinst/U6614  ( .DIN1(\IDinst/n6599 ), .DIN2(n1139), 
        .Q(\IDinst/n6603 ) );
  nnd2s1 \IDinst/U6613  ( .DIN1(\IDinst/n6601 ), .DIN2(\IDinst/n6600 ), 
        .Q(\IDinst/n6602 ) );
  nnd2s1 \IDinst/U6612  ( .DIN1(\IDinst/RegFile[19][6] ), .DIN2(n1097), 
        .Q(\IDinst/n6601 ) );
  nnd2s1 \IDinst/U6611  ( .DIN1(\IDinst/RegFile[18][6] ), .DIN2(n1043), 
        .Q(\IDinst/n6600 ) );
  nnd2s1 \IDinst/U6610  ( .DIN1(\IDinst/n6598 ), .DIN2(\IDinst/n6597 ), 
        .Q(\IDinst/n6599 ) );
  nnd2s1 \IDinst/U6609  ( .DIN1(\IDinst/RegFile[17][6] ), .DIN2(n1097), 
        .Q(\IDinst/n6598 ) );
  nnd2s1 \IDinst/U6608  ( .DIN1(\IDinst/RegFile[16][6] ), .DIN2(n1043), 
        .Q(\IDinst/n6597 ) );
  nnd2s1 \IDinst/U6607  ( .DIN1(\IDinst/n6595 ), .DIN2(\IDinst/n6594 ), 
        .Q(\IDinst/n6596 ) );
  nnd2s1 \IDinst/U6606  ( .DIN1(\IDinst/n6593 ), .DIN2(n644), 
        .Q(\IDinst/n6595 ) );
  nnd2s1 \IDinst/U6605  ( .DIN1(\IDinst/n6572 ), .DIN2(n672), 
        .Q(\IDinst/n6594 ) );
  nnd2s1 \IDinst/U6604  ( .DIN1(\IDinst/n6592 ), .DIN2(\IDinst/n6591 ), 
        .Q(\IDinst/n6593 ) );
  nnd2s1 \IDinst/U6603  ( .DIN1(\IDinst/n6590 ), .DIN2(n1195), 
        .Q(\IDinst/n6592 ) );
  nnd2s1 \IDinst/U6602  ( .DIN1(\IDinst/n6581 ), .DIN2(n1182), 
        .Q(\IDinst/n6591 ) );
  nnd2s1 \IDinst/U6601  ( .DIN1(\IDinst/n6589 ), .DIN2(\IDinst/n6588 ), 
        .Q(\IDinst/n6590 ) );
  nnd2s1 \IDinst/U6600  ( .DIN1(\IDinst/n6587 ), .DIN2(n1171), 
        .Q(\IDinst/n6589 ) );
  nnd2s1 \IDinst/U6599  ( .DIN1(\IDinst/n6584 ), .DIN2(n1139), 
        .Q(\IDinst/n6588 ) );
  nnd2s1 \IDinst/U6598  ( .DIN1(\IDinst/n6586 ), .DIN2(\IDinst/n6585 ), 
        .Q(\IDinst/n6587 ) );
  nnd2s1 \IDinst/U6597  ( .DIN1(\IDinst/RegFile[15][6] ), .DIN2(n1098), 
        .Q(\IDinst/n6586 ) );
  nnd2s1 \IDinst/U6596  ( .DIN1(\IDinst/RegFile[14][6] ), .DIN2(n1043), 
        .Q(\IDinst/n6585 ) );
  nnd2s1 \IDinst/U6595  ( .DIN1(\IDinst/n6583 ), .DIN2(\IDinst/n6582 ), 
        .Q(\IDinst/n6584 ) );
  nnd2s1 \IDinst/U6594  ( .DIN1(\IDinst/RegFile[13][6] ), .DIN2(n1098), 
        .Q(\IDinst/n6583 ) );
  nnd2s1 \IDinst/U6593  ( .DIN1(\IDinst/RegFile[12][6] ), .DIN2(n1043), 
        .Q(\IDinst/n6582 ) );
  nnd2s1 \IDinst/U6592  ( .DIN1(\IDinst/n6580 ), .DIN2(\IDinst/n6579 ), 
        .Q(\IDinst/n6581 ) );
  nnd2s1 \IDinst/U6591  ( .DIN1(\IDinst/n6578 ), .DIN2(n1171), 
        .Q(\IDinst/n6580 ) );
  nnd2s1 \IDinst/U6590  ( .DIN1(\IDinst/n6575 ), .DIN2(n1139), 
        .Q(\IDinst/n6579 ) );
  nnd2s1 \IDinst/U6589  ( .DIN1(\IDinst/n6577 ), .DIN2(\IDinst/n6576 ), 
        .Q(\IDinst/n6578 ) );
  nnd2s1 \IDinst/U6588  ( .DIN1(\IDinst/RegFile[11][6] ), .DIN2(n1098), 
        .Q(\IDinst/n6577 ) );
  nnd2s1 \IDinst/U6587  ( .DIN1(\IDinst/RegFile[10][6] ), .DIN2(n1043), 
        .Q(\IDinst/n6576 ) );
  nnd2s1 \IDinst/U6586  ( .DIN1(\IDinst/n6574 ), .DIN2(\IDinst/n6573 ), 
        .Q(\IDinst/n6575 ) );
  nnd2s1 \IDinst/U6585  ( .DIN1(\IDinst/RegFile[9][6] ), .DIN2(n1098), 
        .Q(\IDinst/n6574 ) );
  nnd2s1 \IDinst/U6584  ( .DIN1(\IDinst/RegFile[8][6] ), .DIN2(n1043), 
        .Q(\IDinst/n6573 ) );
  nnd2s1 \IDinst/U6583  ( .DIN1(\IDinst/n6571 ), .DIN2(\IDinst/n6570 ), 
        .Q(\IDinst/n6572 ) );
  nnd2s1 \IDinst/U6582  ( .DIN1(\IDinst/n6569 ), .DIN2(n1195), 
        .Q(\IDinst/n6571 ) );
  nnd2s1 \IDinst/U6581  ( .DIN1(\IDinst/n6560 ), .DIN2(n1182), 
        .Q(\IDinst/n6570 ) );
  nnd2s1 \IDinst/U6580  ( .DIN1(\IDinst/n6568 ), .DIN2(\IDinst/n6567 ), 
        .Q(\IDinst/n6569 ) );
  nnd2s1 \IDinst/U6579  ( .DIN1(\IDinst/n6566 ), .DIN2(n1171), 
        .Q(\IDinst/n6568 ) );
  nnd2s1 \IDinst/U6578  ( .DIN1(\IDinst/n6563 ), .DIN2(n1139), 
        .Q(\IDinst/n6567 ) );
  nnd2s1 \IDinst/U6577  ( .DIN1(\IDinst/n6565 ), .DIN2(\IDinst/n6564 ), 
        .Q(\IDinst/n6566 ) );
  nnd2s1 \IDinst/U6576  ( .DIN1(\IDinst/RegFile[7][6] ), .DIN2(n1098), 
        .Q(\IDinst/n6565 ) );
  nnd2s1 \IDinst/U6575  ( .DIN1(\IDinst/RegFile[6][6] ), .DIN2(n1043), 
        .Q(\IDinst/n6564 ) );
  nnd2s1 \IDinst/U6574  ( .DIN1(\IDinst/n6562 ), .DIN2(\IDinst/n6561 ), 
        .Q(\IDinst/n6563 ) );
  nnd2s1 \IDinst/U6573  ( .DIN1(\IDinst/RegFile[5][6] ), .DIN2(n1098), 
        .Q(\IDinst/n6562 ) );
  nnd2s1 \IDinst/U6572  ( .DIN1(\IDinst/RegFile[4][6] ), .DIN2(n1043), 
        .Q(\IDinst/n6561 ) );
  nnd2s1 \IDinst/U6571  ( .DIN1(\IDinst/n6559 ), .DIN2(\IDinst/n6558 ), 
        .Q(\IDinst/n6560 ) );
  nnd2s1 \IDinst/U6570  ( .DIN1(\IDinst/n6557 ), .DIN2(n1171), 
        .Q(\IDinst/n6559 ) );
  nnd2s1 \IDinst/U6569  ( .DIN1(\IDinst/n6554 ), .DIN2(n1139), 
        .Q(\IDinst/n6558 ) );
  nnd2s1 \IDinst/U6568  ( .DIN1(\IDinst/n6556 ), .DIN2(\IDinst/n6555 ), 
        .Q(\IDinst/n6557 ) );
  nnd2s1 \IDinst/U6567  ( .DIN1(\IDinst/RegFile[3][6] ), .DIN2(n1098), 
        .Q(\IDinst/n6556 ) );
  nnd2s1 \IDinst/U6566  ( .DIN1(\IDinst/RegFile[2][6] ), .DIN2(n1042), 
        .Q(\IDinst/n6555 ) );
  nnd2s1 \IDinst/U6565  ( .DIN1(\IDinst/n6553 ), .DIN2(\IDinst/n6552 ), 
        .Q(\IDinst/n6554 ) );
  nnd2s1 \IDinst/U6564  ( .DIN1(\IDinst/RegFile[1][6] ), .DIN2(n1098), 
        .Q(\IDinst/n6553 ) );
  nnd2s1 \IDinst/U6563  ( .DIN1(\IDinst/RegFile[0][6] ), .DIN2(n1042), 
        .Q(\IDinst/n6552 ) );
  nnd2s1 \IDinst/U6562  ( .DIN1(\IDinst/n6551 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n5958 ) );
  nnd2s1 \IDinst/U6561  ( .DIN1(\IDinst/n6506 ), .DIN2(n635), 
        .Q(\IDinst/n5959 ) );
  nnd2s1 \IDinst/U6560  ( .DIN1(\IDinst/n6550 ), .DIN2(\IDinst/n6549 ), 
        .Q(\IDinst/n6551 ) );
  nnd2s1 \IDinst/U6559  ( .DIN1(\IDinst/n6548 ), .DIN2(n643), 
        .Q(\IDinst/n6550 ) );
  nnd2s1 \IDinst/U6558  ( .DIN1(\IDinst/n6527 ), .DIN2(n670), 
        .Q(\IDinst/n6549 ) );
  nnd2s1 \IDinst/U6557  ( .DIN1(\IDinst/n6547 ), .DIN2(\IDinst/n6546 ), 
        .Q(\IDinst/n6548 ) );
  nnd2s1 \IDinst/U6556  ( .DIN1(\IDinst/n6545 ), .DIN2(n1195), 
        .Q(\IDinst/n6547 ) );
  nnd2s1 \IDinst/U6555  ( .DIN1(\IDinst/n6536 ), .DIN2(n1182), 
        .Q(\IDinst/n6546 ) );
  nnd2s1 \IDinst/U6554  ( .DIN1(\IDinst/n6544 ), .DIN2(\IDinst/n6543 ), 
        .Q(\IDinst/n6545 ) );
  nnd2s1 \IDinst/U6553  ( .DIN1(\IDinst/n6542 ), .DIN2(n1171), 
        .Q(\IDinst/n6544 ) );
  nnd2s1 \IDinst/U6552  ( .DIN1(\IDinst/n6539 ), .DIN2(n1140), 
        .Q(\IDinst/n6543 ) );
  nnd2s1 \IDinst/U6551  ( .DIN1(\IDinst/n6541 ), .DIN2(\IDinst/n6540 ), 
        .Q(\IDinst/n6542 ) );
  nnd2s1 \IDinst/U6550  ( .DIN1(\IDinst/RegFile[31][5] ), .DIN2(n1098), 
        .Q(\IDinst/n6541 ) );
  nnd2s1 \IDinst/U6549  ( .DIN1(\IDinst/RegFile[30][5] ), .DIN2(n1042), 
        .Q(\IDinst/n6540 ) );
  nnd2s1 \IDinst/U6548  ( .DIN1(\IDinst/n6538 ), .DIN2(\IDinst/n6537 ), 
        .Q(\IDinst/n6539 ) );
  nnd2s1 \IDinst/U6547  ( .DIN1(\IDinst/RegFile[29][5] ), .DIN2(n1099), 
        .Q(\IDinst/n6538 ) );
  nnd2s1 \IDinst/U6546  ( .DIN1(\IDinst/RegFile[28][5] ), .DIN2(n1042), 
        .Q(\IDinst/n6537 ) );
  nnd2s1 \IDinst/U6545  ( .DIN1(\IDinst/n6535 ), .DIN2(\IDinst/n6534 ), 
        .Q(\IDinst/n6536 ) );
  nnd2s1 \IDinst/U6544  ( .DIN1(\IDinst/n6533 ), .DIN2(n1171), 
        .Q(\IDinst/n6535 ) );
  nnd2s1 \IDinst/U6543  ( .DIN1(\IDinst/n6530 ), .DIN2(n1140), 
        .Q(\IDinst/n6534 ) );
  nnd2s1 \IDinst/U6542  ( .DIN1(\IDinst/n6532 ), .DIN2(\IDinst/n6531 ), 
        .Q(\IDinst/n6533 ) );
  nnd2s1 \IDinst/U6541  ( .DIN1(\IDinst/RegFile[27][5] ), .DIN2(n1099), 
        .Q(\IDinst/n6532 ) );
  nnd2s1 \IDinst/U6540  ( .DIN1(\IDinst/RegFile[26][5] ), .DIN2(n1042), 
        .Q(\IDinst/n6531 ) );
  nnd2s1 \IDinst/U6539  ( .DIN1(\IDinst/n6529 ), .DIN2(\IDinst/n6528 ), 
        .Q(\IDinst/n6530 ) );
  nnd2s1 \IDinst/U6538  ( .DIN1(\IDinst/RegFile[25][5] ), .DIN2(n1099), 
        .Q(\IDinst/n6529 ) );
  nnd2s1 \IDinst/U6537  ( .DIN1(\IDinst/RegFile[24][5] ), .DIN2(n1042), 
        .Q(\IDinst/n6528 ) );
  nnd2s1 \IDinst/U6536  ( .DIN1(\IDinst/n6526 ), .DIN2(\IDinst/n6525 ), 
        .Q(\IDinst/n6527 ) );
  nnd2s1 \IDinst/U6535  ( .DIN1(\IDinst/n6524 ), .DIN2(n1195), 
        .Q(\IDinst/n6526 ) );
  nnd2s1 \IDinst/U6534  ( .DIN1(\IDinst/n6515 ), .DIN2(n1182), 
        .Q(\IDinst/n6525 ) );
  nnd2s1 \IDinst/U6533  ( .DIN1(\IDinst/n6523 ), .DIN2(\IDinst/n6522 ), 
        .Q(\IDinst/n6524 ) );
  nnd2s1 \IDinst/U6532  ( .DIN1(\IDinst/n6521 ), .DIN2(n1171), 
        .Q(\IDinst/n6523 ) );
  nnd2s1 \IDinst/U6531  ( .DIN1(\IDinst/n6518 ), .DIN2(n1140), 
        .Q(\IDinst/n6522 ) );
  nnd2s1 \IDinst/U6530  ( .DIN1(\IDinst/n6520 ), .DIN2(\IDinst/n6519 ), 
        .Q(\IDinst/n6521 ) );
  nnd2s1 \IDinst/U6529  ( .DIN1(\IDinst/RegFile[23][5] ), .DIN2(n1099), 
        .Q(\IDinst/n6520 ) );
  nnd2s1 \IDinst/U6528  ( .DIN1(\IDinst/RegFile[22][5] ), .DIN2(n1042), 
        .Q(\IDinst/n6519 ) );
  nnd2s1 \IDinst/U6527  ( .DIN1(\IDinst/n6517 ), .DIN2(\IDinst/n6516 ), 
        .Q(\IDinst/n6518 ) );
  nnd2s1 \IDinst/U6526  ( .DIN1(\IDinst/RegFile[21][5] ), .DIN2(n1099), 
        .Q(\IDinst/n6517 ) );
  nnd2s1 \IDinst/U6525  ( .DIN1(\IDinst/RegFile[20][5] ), .DIN2(n1042), 
        .Q(\IDinst/n6516 ) );
  nnd2s1 \IDinst/U6524  ( .DIN1(\IDinst/n6514 ), .DIN2(\IDinst/n6513 ), 
        .Q(\IDinst/n6515 ) );
  nnd2s1 \IDinst/U6523  ( .DIN1(\IDinst/n6512 ), .DIN2(n1171), 
        .Q(\IDinst/n6514 ) );
  nnd2s1 \IDinst/U6522  ( .DIN1(\IDinst/n6509 ), .DIN2(n1140), 
        .Q(\IDinst/n6513 ) );
  nnd2s1 \IDinst/U6521  ( .DIN1(\IDinst/n6511 ), .DIN2(\IDinst/n6510 ), 
        .Q(\IDinst/n6512 ) );
  nnd2s1 \IDinst/U6520  ( .DIN1(\IDinst/RegFile[19][5] ), .DIN2(n1099), 
        .Q(\IDinst/n6511 ) );
  nnd2s1 \IDinst/U6519  ( .DIN1(\IDinst/RegFile[18][5] ), .DIN2(n1042), 
        .Q(\IDinst/n6510 ) );
  nnd2s1 \IDinst/U6518  ( .DIN1(\IDinst/n6508 ), .DIN2(\IDinst/n6507 ), 
        .Q(\IDinst/n6509 ) );
  nnd2s1 \IDinst/U6517  ( .DIN1(\IDinst/RegFile[17][5] ), .DIN2(n1099), 
        .Q(\IDinst/n6508 ) );
  nnd2s1 \IDinst/U6516  ( .DIN1(\IDinst/RegFile[16][5] ), .DIN2(n1042), 
        .Q(\IDinst/n6507 ) );
  nnd2s1 \IDinst/U6515  ( .DIN1(\IDinst/n6505 ), .DIN2(\IDinst/n6504 ), 
        .Q(\IDinst/n6506 ) );
  nnd2s1 \IDinst/U6514  ( .DIN1(\IDinst/n6503 ), .DIN2(n642), 
        .Q(\IDinst/n6505 ) );
  nnd2s1 \IDinst/U6513  ( .DIN1(\IDinst/n6482 ), .DIN2(n673), 
        .Q(\IDinst/n6504 ) );
  nnd2s1 \IDinst/U6512  ( .DIN1(\IDinst/n6502 ), .DIN2(\IDinst/n6501 ), 
        .Q(\IDinst/n6503 ) );
  nnd2s1 \IDinst/U6511  ( .DIN1(\IDinst/n6500 ), .DIN2(n1195), 
        .Q(\IDinst/n6502 ) );
  nnd2s1 \IDinst/U6510  ( .DIN1(\IDinst/n6491 ), .DIN2(n1182), 
        .Q(\IDinst/n6501 ) );
  nnd2s1 \IDinst/U6509  ( .DIN1(\IDinst/n6499 ), .DIN2(\IDinst/n6498 ), 
        .Q(\IDinst/n6500 ) );
  nnd2s1 \IDinst/U6508  ( .DIN1(\IDinst/n6497 ), .DIN2(n1170), 
        .Q(\IDinst/n6499 ) );
  nnd2s1 \IDinst/U6507  ( .DIN1(\IDinst/n6494 ), .DIN2(n1140), 
        .Q(\IDinst/n6498 ) );
  nnd2s1 \IDinst/U6506  ( .DIN1(\IDinst/n6496 ), .DIN2(\IDinst/n6495 ), 
        .Q(\IDinst/n6497 ) );
  nnd2s1 \IDinst/U6505  ( .DIN1(\IDinst/RegFile[15][5] ), .DIN2(n1099), 
        .Q(\IDinst/n6496 ) );
  nnd2s1 \IDinst/U6504  ( .DIN1(\IDinst/RegFile[14][5] ), .DIN2(n1042), 
        .Q(\IDinst/n6495 ) );
  nnd2s1 \IDinst/U6503  ( .DIN1(\IDinst/n6493 ), .DIN2(\IDinst/n6492 ), 
        .Q(\IDinst/n6494 ) );
  nnd2s1 \IDinst/U6502  ( .DIN1(\IDinst/RegFile[13][5] ), .DIN2(n1099), 
        .Q(\IDinst/n6493 ) );
  nnd2s1 \IDinst/U6501  ( .DIN1(\IDinst/RegFile[12][5] ), .DIN2(n1042), 
        .Q(\IDinst/n6492 ) );
  nnd2s1 \IDinst/U6500  ( .DIN1(\IDinst/n6490 ), .DIN2(\IDinst/n6489 ), 
        .Q(\IDinst/n6491 ) );
  nnd2s1 \IDinst/U6499  ( .DIN1(\IDinst/n6488 ), .DIN2(n1170), 
        .Q(\IDinst/n6490 ) );
  nnd2s1 \IDinst/U6498  ( .DIN1(\IDinst/n6485 ), .DIN2(n1140), 
        .Q(\IDinst/n6489 ) );
  nnd2s1 \IDinst/U6497  ( .DIN1(\IDinst/n6487 ), .DIN2(\IDinst/n6486 ), 
        .Q(\IDinst/n6488 ) );
  nnd2s1 \IDinst/U6496  ( .DIN1(\IDinst/RegFile[11][5] ), .DIN2(n1100), 
        .Q(\IDinst/n6487 ) );
  nnd2s1 \IDinst/U6495  ( .DIN1(\IDinst/RegFile[10][5] ), .DIN2(n1042), 
        .Q(\IDinst/n6486 ) );
  nnd2s1 \IDinst/U6494  ( .DIN1(\IDinst/n6484 ), .DIN2(\IDinst/n6483 ), 
        .Q(\IDinst/n6485 ) );
  nnd2s1 \IDinst/U6493  ( .DIN1(\IDinst/RegFile[9][5] ), .DIN2(n1100), 
        .Q(\IDinst/n6484 ) );
  nnd2s1 \IDinst/U6492  ( .DIN1(\IDinst/RegFile[8][5] ), .DIN2(n1041), 
        .Q(\IDinst/n6483 ) );
  nnd2s1 \IDinst/U6491  ( .DIN1(\IDinst/n6481 ), .DIN2(\IDinst/n6480 ), 
        .Q(\IDinst/n6482 ) );
  nnd2s1 \IDinst/U6490  ( .DIN1(\IDinst/n6479 ), .DIN2(n1195), 
        .Q(\IDinst/n6481 ) );
  nnd2s1 \IDinst/U6489  ( .DIN1(\IDinst/n6470 ), .DIN2(n1182), 
        .Q(\IDinst/n6480 ) );
  nnd2s1 \IDinst/U6488  ( .DIN1(\IDinst/n6478 ), .DIN2(\IDinst/n6477 ), 
        .Q(\IDinst/n6479 ) );
  nnd2s1 \IDinst/U6487  ( .DIN1(\IDinst/n6476 ), .DIN2(n1170), 
        .Q(\IDinst/n6478 ) );
  nnd2s1 \IDinst/U6486  ( .DIN1(\IDinst/n6473 ), .DIN2(n1140), 
        .Q(\IDinst/n6477 ) );
  nnd2s1 \IDinst/U6485  ( .DIN1(\IDinst/n6475 ), .DIN2(\IDinst/n6474 ), 
        .Q(\IDinst/n6476 ) );
  nnd2s1 \IDinst/U6484  ( .DIN1(\IDinst/RegFile[7][5] ), .DIN2(n1100), 
        .Q(\IDinst/n6475 ) );
  nnd2s1 \IDinst/U6483  ( .DIN1(\IDinst/RegFile[6][5] ), .DIN2(n1041), 
        .Q(\IDinst/n6474 ) );
  nnd2s1 \IDinst/U6482  ( .DIN1(\IDinst/n6472 ), .DIN2(\IDinst/n6471 ), 
        .Q(\IDinst/n6473 ) );
  nnd2s1 \IDinst/U6481  ( .DIN1(\IDinst/RegFile[5][5] ), .DIN2(n1100), 
        .Q(\IDinst/n6472 ) );
  nnd2s1 \IDinst/U6480  ( .DIN1(\IDinst/RegFile[4][5] ), .DIN2(n1041), 
        .Q(\IDinst/n6471 ) );
  nnd2s1 \IDinst/U6479  ( .DIN1(\IDinst/n6469 ), .DIN2(\IDinst/n6468 ), 
        .Q(\IDinst/n6470 ) );
  nnd2s1 \IDinst/U6478  ( .DIN1(\IDinst/n6467 ), .DIN2(n1170), 
        .Q(\IDinst/n6469 ) );
  nnd2s1 \IDinst/U6477  ( .DIN1(\IDinst/n6464 ), .DIN2(n1140), 
        .Q(\IDinst/n6468 ) );
  nnd2s1 \IDinst/U6476  ( .DIN1(\IDinst/n6466 ), .DIN2(\IDinst/n6465 ), 
        .Q(\IDinst/n6467 ) );
  nnd2s1 \IDinst/U6475  ( .DIN1(\IDinst/RegFile[3][5] ), .DIN2(n1100), 
        .Q(\IDinst/n6466 ) );
  nnd2s1 \IDinst/U6474  ( .DIN1(\IDinst/RegFile[2][5] ), .DIN2(n1041), 
        .Q(\IDinst/n6465 ) );
  nnd2s1 \IDinst/U6473  ( .DIN1(\IDinst/n6463 ), .DIN2(\IDinst/n6462 ), 
        .Q(\IDinst/n6464 ) );
  nnd2s1 \IDinst/U6472  ( .DIN1(\IDinst/RegFile[1][5] ), .DIN2(n1100), 
        .Q(\IDinst/n6463 ) );
  nnd2s1 \IDinst/U6471  ( .DIN1(\IDinst/RegFile[0][5] ), .DIN2(n1041), 
        .Q(\IDinst/n6462 ) );
  nnd2s1 \IDinst/U6470  ( .DIN1(\IDinst/n6461 ), .DIN2(n539), 
        .Q(\IDinst/n5956 ) );
  nnd2s1 \IDinst/U6469  ( .DIN1(\IDinst/n6416 ), .DIN2(n636), 
        .Q(\IDinst/n5957 ) );
  nnd2s1 \IDinst/U6468  ( .DIN1(\IDinst/n6460 ), .DIN2(\IDinst/n6459 ), 
        .Q(\IDinst/n6461 ) );
  nnd2s1 \IDinst/U6467  ( .DIN1(\IDinst/n6458 ), .DIN2(n644), 
        .Q(\IDinst/n6460 ) );
  nnd2s1 \IDinst/U6466  ( .DIN1(\IDinst/n6437 ), .DIN2(n671), 
        .Q(\IDinst/n6459 ) );
  nnd2s1 \IDinst/U6465  ( .DIN1(\IDinst/n6457 ), .DIN2(\IDinst/n6456 ), 
        .Q(\IDinst/n6458 ) );
  nnd2s1 \IDinst/U6464  ( .DIN1(\IDinst/n6455 ), .DIN2(n1195), 
        .Q(\IDinst/n6457 ) );
  nnd2s1 \IDinst/U6463  ( .DIN1(\IDinst/n6446 ), .DIN2(n1182), 
        .Q(\IDinst/n6456 ) );
  nnd2s1 \IDinst/U6462  ( .DIN1(\IDinst/n6454 ), .DIN2(\IDinst/n6453 ), 
        .Q(\IDinst/n6455 ) );
  nnd2s1 \IDinst/U6461  ( .DIN1(\IDinst/n6452 ), .DIN2(n1170), 
        .Q(\IDinst/n6454 ) );
  nnd2s1 \IDinst/U6460  ( .DIN1(\IDinst/n6449 ), .DIN2(n1140), 
        .Q(\IDinst/n6453 ) );
  nnd2s1 \IDinst/U6459  ( .DIN1(\IDinst/n6451 ), .DIN2(\IDinst/n6450 ), 
        .Q(\IDinst/n6452 ) );
  nnd2s1 \IDinst/U6458  ( .DIN1(\IDinst/RegFile[31][4] ), .DIN2(n1100), 
        .Q(\IDinst/n6451 ) );
  nnd2s1 \IDinst/U6457  ( .DIN1(\IDinst/RegFile[30][4] ), .DIN2(n1041), 
        .Q(\IDinst/n6450 ) );
  nnd2s1 \IDinst/U6456  ( .DIN1(\IDinst/n6448 ), .DIN2(\IDinst/n6447 ), 
        .Q(\IDinst/n6449 ) );
  nnd2s1 \IDinst/U6455  ( .DIN1(\IDinst/RegFile[29][4] ), .DIN2(n1100), 
        .Q(\IDinst/n6448 ) );
  nnd2s1 \IDinst/U6454  ( .DIN1(\IDinst/RegFile[28][4] ), .DIN2(n1041), 
        .Q(\IDinst/n6447 ) );
  nnd2s1 \IDinst/U6453  ( .DIN1(\IDinst/n6445 ), .DIN2(\IDinst/n6444 ), 
        .Q(\IDinst/n6446 ) );
  nnd2s1 \IDinst/U6452  ( .DIN1(\IDinst/n6443 ), .DIN2(n1170), 
        .Q(\IDinst/n6445 ) );
  nnd2s1 \IDinst/U6451  ( .DIN1(\IDinst/n6440 ), .DIN2(n1140), 
        .Q(\IDinst/n6444 ) );
  nnd2s1 \IDinst/U6450  ( .DIN1(\IDinst/n6442 ), .DIN2(\IDinst/n6441 ), 
        .Q(\IDinst/n6443 ) );
  nnd2s1 \IDinst/U6449  ( .DIN1(\IDinst/RegFile[27][4] ), .DIN2(n1100), 
        .Q(\IDinst/n6442 ) );
  nnd2s1 \IDinst/U6448  ( .DIN1(\IDinst/RegFile[26][4] ), .DIN2(n1041), 
        .Q(\IDinst/n6441 ) );
  nnd2s1 \IDinst/U6447  ( .DIN1(\IDinst/n6439 ), .DIN2(\IDinst/n6438 ), 
        .Q(\IDinst/n6440 ) );
  nnd2s1 \IDinst/U6446  ( .DIN1(\IDinst/RegFile[25][4] ), .DIN2(n1101), 
        .Q(\IDinst/n6439 ) );
  nnd2s1 \IDinst/U6445  ( .DIN1(\IDinst/RegFile[24][4] ), .DIN2(n1041), 
        .Q(\IDinst/n6438 ) );
  nnd2s1 \IDinst/U6444  ( .DIN1(\IDinst/n6436 ), .DIN2(\IDinst/n6435 ), 
        .Q(\IDinst/n6437 ) );
  nnd2s1 \IDinst/U6443  ( .DIN1(\IDinst/n6434 ), .DIN2(n1196), 
        .Q(\IDinst/n6436 ) );
  nnd2s1 \IDinst/U6442  ( .DIN1(\IDinst/n6425 ), .DIN2(n1181), 
        .Q(\IDinst/n6435 ) );
  nnd2s1 \IDinst/U6441  ( .DIN1(\IDinst/n6433 ), .DIN2(\IDinst/n6432 ), 
        .Q(\IDinst/n6434 ) );
  nnd2s1 \IDinst/U6440  ( .DIN1(\IDinst/n6431 ), .DIN2(n1170), 
        .Q(\IDinst/n6433 ) );
  nnd2s1 \IDinst/U6439  ( .DIN1(\IDinst/n6428 ), .DIN2(n1140), 
        .Q(\IDinst/n6432 ) );
  nnd2s1 \IDinst/U6438  ( .DIN1(\IDinst/n6430 ), .DIN2(\IDinst/n6429 ), 
        .Q(\IDinst/n6431 ) );
  nnd2s1 \IDinst/U6437  ( .DIN1(\IDinst/RegFile[23][4] ), .DIN2(n1101), 
        .Q(\IDinst/n6430 ) );
  nnd2s1 \IDinst/U6436  ( .DIN1(\IDinst/RegFile[22][4] ), .DIN2(n1041), 
        .Q(\IDinst/n6429 ) );
  nnd2s1 \IDinst/U6435  ( .DIN1(\IDinst/n6427 ), .DIN2(\IDinst/n6426 ), 
        .Q(\IDinst/n6428 ) );
  nnd2s1 \IDinst/U6434  ( .DIN1(\IDinst/RegFile[21][4] ), .DIN2(n1101), 
        .Q(\IDinst/n6427 ) );
  nnd2s1 \IDinst/U6433  ( .DIN1(\IDinst/RegFile[20][4] ), .DIN2(n1041), 
        .Q(\IDinst/n6426 ) );
  nnd2s1 \IDinst/U6432  ( .DIN1(\IDinst/n6424 ), .DIN2(\IDinst/n6423 ), 
        .Q(\IDinst/n6425 ) );
  nnd2s1 \IDinst/U6431  ( .DIN1(\IDinst/n6422 ), .DIN2(n1170), 
        .Q(\IDinst/n6424 ) );
  nnd2s1 \IDinst/U6430  ( .DIN1(\IDinst/n6419 ), .DIN2(n1140), 
        .Q(\IDinst/n6423 ) );
  nnd2s1 \IDinst/U6429  ( .DIN1(\IDinst/n6421 ), .DIN2(\IDinst/n6420 ), 
        .Q(\IDinst/n6422 ) );
  nnd2s1 \IDinst/U6428  ( .DIN1(\IDinst/RegFile[19][4] ), .DIN2(n1101), 
        .Q(\IDinst/n6421 ) );
  nnd2s1 \IDinst/U6427  ( .DIN1(\IDinst/RegFile[18][4] ), .DIN2(n1041), 
        .Q(\IDinst/n6420 ) );
  nnd2s1 \IDinst/U6426  ( .DIN1(\IDinst/n6418 ), .DIN2(\IDinst/n6417 ), 
        .Q(\IDinst/n6419 ) );
  nnd2s1 \IDinst/U6425  ( .DIN1(\IDinst/RegFile[17][4] ), .DIN2(n1101), 
        .Q(\IDinst/n6418 ) );
  nnd2s1 \IDinst/U6424  ( .DIN1(\IDinst/RegFile[16][4] ), .DIN2(n1041), 
        .Q(\IDinst/n6417 ) );
  nnd2s1 \IDinst/U6423  ( .DIN1(\IDinst/n6415 ), .DIN2(\IDinst/n6414 ), 
        .Q(\IDinst/n6416 ) );
  nnd2s1 \IDinst/U6422  ( .DIN1(\IDinst/n6413 ), .DIN2(n643), 
        .Q(\IDinst/n6415 ) );
  nnd2s1 \IDinst/U6421  ( .DIN1(\IDinst/n6392 ), .DIN2(n672), 
        .Q(\IDinst/n6414 ) );
  nnd2s1 \IDinst/U6420  ( .DIN1(\IDinst/n6412 ), .DIN2(\IDinst/n6411 ), 
        .Q(\IDinst/n6413 ) );
  nnd2s1 \IDinst/U6419  ( .DIN1(\IDinst/n6410 ), .DIN2(n1196), 
        .Q(\IDinst/n6412 ) );
  nnd2s1 \IDinst/U6418  ( .DIN1(\IDinst/n6401 ), .DIN2(n1181), 
        .Q(\IDinst/n6411 ) );
  nnd2s1 \IDinst/U6417  ( .DIN1(\IDinst/n6409 ), .DIN2(\IDinst/n6408 ), 
        .Q(\IDinst/n6410 ) );
  nnd2s1 \IDinst/U6416  ( .DIN1(\IDinst/n6407 ), .DIN2(n1170), 
        .Q(\IDinst/n6409 ) );
  nnd2s1 \IDinst/U6415  ( .DIN1(\IDinst/n6404 ), .DIN2(n1140), 
        .Q(\IDinst/n6408 ) );
  nnd2s1 \IDinst/U6414  ( .DIN1(\IDinst/n6406 ), .DIN2(\IDinst/n6405 ), 
        .Q(\IDinst/n6407 ) );
  nnd2s1 \IDinst/U6413  ( .DIN1(\IDinst/RegFile[15][4] ), .DIN2(n1101), 
        .Q(\IDinst/n6406 ) );
  nnd2s1 \IDinst/U6412  ( .DIN1(\IDinst/RegFile[14][4] ), .DIN2(n1040), 
        .Q(\IDinst/n6405 ) );
  nnd2s1 \IDinst/U6411  ( .DIN1(\IDinst/n6403 ), .DIN2(\IDinst/n6402 ), 
        .Q(\IDinst/n6404 ) );
  nnd2s1 \IDinst/U6410  ( .DIN1(\IDinst/RegFile[13][4] ), .DIN2(n1101), 
        .Q(\IDinst/n6403 ) );
  nnd2s1 \IDinst/U6409  ( .DIN1(\IDinst/RegFile[12][4] ), .DIN2(n1040), 
        .Q(\IDinst/n6402 ) );
  nnd2s1 \IDinst/U6408  ( .DIN1(\IDinst/n6400 ), .DIN2(\IDinst/n6399 ), 
        .Q(\IDinst/n6401 ) );
  nnd2s1 \IDinst/U6407  ( .DIN1(\IDinst/n6398 ), .DIN2(n1169), 
        .Q(\IDinst/n6400 ) );
  nnd2s1 \IDinst/U6406  ( .DIN1(\IDinst/n6395 ), .DIN2(n1141), 
        .Q(\IDinst/n6399 ) );
  nnd2s1 \IDinst/U6405  ( .DIN1(\IDinst/n6397 ), .DIN2(\IDinst/n6396 ), 
        .Q(\IDinst/n6398 ) );
  nnd2s1 \IDinst/U6404  ( .DIN1(\IDinst/RegFile[11][4] ), .DIN2(n1101), 
        .Q(\IDinst/n6397 ) );
  nnd2s1 \IDinst/U6403  ( .DIN1(\IDinst/RegFile[10][4] ), .DIN2(n1040), 
        .Q(\IDinst/n6396 ) );
  nnd2s1 \IDinst/U6402  ( .DIN1(\IDinst/n6394 ), .DIN2(\IDinst/n6393 ), 
        .Q(\IDinst/n6395 ) );
  nnd2s1 \IDinst/U6401  ( .DIN1(\IDinst/RegFile[9][4] ), .DIN2(n1101), 
        .Q(\IDinst/n6394 ) );
  nnd2s1 \IDinst/U6400  ( .DIN1(\IDinst/RegFile[8][4] ), .DIN2(n1040), 
        .Q(\IDinst/n6393 ) );
  nnd2s1 \IDinst/U6399  ( .DIN1(\IDinst/n6391 ), .DIN2(\IDinst/n6390 ), 
        .Q(\IDinst/n6392 ) );
  nnd2s1 \IDinst/U6398  ( .DIN1(\IDinst/n6389 ), .DIN2(n1196), 
        .Q(\IDinst/n6391 ) );
  nnd2s1 \IDinst/U6397  ( .DIN1(\IDinst/n6380 ), .DIN2(n1183), 
        .Q(\IDinst/n6390 ) );
  nnd2s1 \IDinst/U6396  ( .DIN1(\IDinst/n6388 ), .DIN2(\IDinst/n6387 ), 
        .Q(\IDinst/n6389 ) );
  nnd2s1 \IDinst/U6395  ( .DIN1(\IDinst/n6386 ), .DIN2(n1169), 
        .Q(\IDinst/n6388 ) );
  nnd2s1 \IDinst/U6394  ( .DIN1(\IDinst/n6383 ), .DIN2(n1141), 
        .Q(\IDinst/n6387 ) );
  nnd2s1 \IDinst/U6393  ( .DIN1(\IDinst/n6385 ), .DIN2(\IDinst/n6384 ), 
        .Q(\IDinst/n6386 ) );
  nnd2s1 \IDinst/U6392  ( .DIN1(\IDinst/RegFile[7][4] ), .DIN2(n1102), 
        .Q(\IDinst/n6385 ) );
  nnd2s1 \IDinst/U6391  ( .DIN1(\IDinst/RegFile[6][4] ), .DIN2(n1040), 
        .Q(\IDinst/n6384 ) );
  nnd2s1 \IDinst/U6390  ( .DIN1(\IDinst/n6382 ), .DIN2(\IDinst/n6381 ), 
        .Q(\IDinst/n6383 ) );
  nnd2s1 \IDinst/U6389  ( .DIN1(\IDinst/RegFile[5][4] ), .DIN2(n1102), 
        .Q(\IDinst/n6382 ) );
  nnd2s1 \IDinst/U6388  ( .DIN1(\IDinst/RegFile[4][4] ), .DIN2(n1040), 
        .Q(\IDinst/n6381 ) );
  nnd2s1 \IDinst/U6387  ( .DIN1(\IDinst/n6379 ), .DIN2(\IDinst/n6378 ), 
        .Q(\IDinst/n6380 ) );
  nnd2s1 \IDinst/U6386  ( .DIN1(\IDinst/n6377 ), .DIN2(n1169), 
        .Q(\IDinst/n6379 ) );
  nnd2s1 \IDinst/U6385  ( .DIN1(\IDinst/n6374 ), .DIN2(n1141), 
        .Q(\IDinst/n6378 ) );
  nnd2s1 \IDinst/U6384  ( .DIN1(\IDinst/n6376 ), .DIN2(\IDinst/n6375 ), 
        .Q(\IDinst/n6377 ) );
  nnd2s1 \IDinst/U6383  ( .DIN1(\IDinst/RegFile[3][4] ), .DIN2(n1102), 
        .Q(\IDinst/n6376 ) );
  nnd2s1 \IDinst/U6382  ( .DIN1(\IDinst/RegFile[2][4] ), .DIN2(n1040), 
        .Q(\IDinst/n6375 ) );
  nnd2s1 \IDinst/U6381  ( .DIN1(\IDinst/n6373 ), .DIN2(\IDinst/n6372 ), 
        .Q(\IDinst/n6374 ) );
  nnd2s1 \IDinst/U6380  ( .DIN1(\IDinst/RegFile[1][4] ), .DIN2(n1102), 
        .Q(\IDinst/n6373 ) );
  nnd2s1 \IDinst/U6379  ( .DIN1(\IDinst/RegFile[0][4] ), .DIN2(n1040), 
        .Q(\IDinst/n6372 ) );
  nnd2s1 \IDinst/U6378  ( .DIN1(\IDinst/n6371 ), .DIN2(n539), 
        .Q(\IDinst/n5954 ) );
  nnd2s1 \IDinst/U6377  ( .DIN1(\IDinst/n6326 ), .DIN2(n635), 
        .Q(\IDinst/n5955 ) );
  nnd2s1 \IDinst/U6376  ( .DIN1(\IDinst/n6370 ), .DIN2(\IDinst/n6369 ), 
        .Q(\IDinst/n6371 ) );
  nnd2s1 \IDinst/U6375  ( .DIN1(\IDinst/n6368 ), .DIN2(n642), 
        .Q(\IDinst/n6370 ) );
  nnd2s1 \IDinst/U6374  ( .DIN1(\IDinst/n6347 ), .DIN2(n670), 
        .Q(\IDinst/n6369 ) );
  nnd2s1 \IDinst/U6373  ( .DIN1(\IDinst/n6367 ), .DIN2(\IDinst/n6366 ), 
        .Q(\IDinst/n6368 ) );
  nnd2s1 \IDinst/U6372  ( .DIN1(\IDinst/n6365 ), .DIN2(n1196), 
        .Q(\IDinst/n6367 ) );
  nnd2s1 \IDinst/U6371  ( .DIN1(\IDinst/n6356 ), .DIN2(n1182), 
        .Q(\IDinst/n6366 ) );
  nnd2s1 \IDinst/U6370  ( .DIN1(\IDinst/n6364 ), .DIN2(\IDinst/n6363 ), 
        .Q(\IDinst/n6365 ) );
  nnd2s1 \IDinst/U6369  ( .DIN1(\IDinst/n6362 ), .DIN2(n1169), 
        .Q(\IDinst/n6364 ) );
  nnd2s1 \IDinst/U6368  ( .DIN1(\IDinst/n6359 ), .DIN2(n1141), 
        .Q(\IDinst/n6363 ) );
  nnd2s1 \IDinst/U6367  ( .DIN1(\IDinst/n6361 ), .DIN2(\IDinst/n6360 ), 
        .Q(\IDinst/n6362 ) );
  nnd2s1 \IDinst/U6366  ( .DIN1(\IDinst/RegFile[31][3] ), .DIN2(n1102), 
        .Q(\IDinst/n6361 ) );
  nnd2s1 \IDinst/U6365  ( .DIN1(\IDinst/RegFile[30][3] ), .DIN2(n1040), 
        .Q(\IDinst/n6360 ) );
  nnd2s1 \IDinst/U6364  ( .DIN1(\IDinst/n6358 ), .DIN2(\IDinst/n6357 ), 
        .Q(\IDinst/n6359 ) );
  nnd2s1 \IDinst/U6363  ( .DIN1(\IDinst/RegFile[29][3] ), .DIN2(n1102), 
        .Q(\IDinst/n6358 ) );
  nnd2s1 \IDinst/U6362  ( .DIN1(\IDinst/RegFile[28][3] ), .DIN2(n1040), 
        .Q(\IDinst/n6357 ) );
  nnd2s1 \IDinst/U6361  ( .DIN1(\IDinst/n6355 ), .DIN2(\IDinst/n6354 ), 
        .Q(\IDinst/n6356 ) );
  nnd2s1 \IDinst/U6360  ( .DIN1(\IDinst/n6353 ), .DIN2(n1169), 
        .Q(\IDinst/n6355 ) );
  nnd2s1 \IDinst/U6359  ( .DIN1(\IDinst/n6350 ), .DIN2(n1141), 
        .Q(\IDinst/n6354 ) );
  nnd2s1 \IDinst/U6358  ( .DIN1(\IDinst/n6352 ), .DIN2(\IDinst/n6351 ), 
        .Q(\IDinst/n6353 ) );
  nnd2s1 \IDinst/U6357  ( .DIN1(\IDinst/RegFile[27][3] ), .DIN2(n1102), 
        .Q(\IDinst/n6352 ) );
  nnd2s1 \IDinst/U6356  ( .DIN1(\IDinst/RegFile[26][3] ), .DIN2(n1040), 
        .Q(\IDinst/n6351 ) );
  nnd2s1 \IDinst/U6355  ( .DIN1(\IDinst/n6349 ), .DIN2(\IDinst/n6348 ), 
        .Q(\IDinst/n6350 ) );
  nnd2s1 \IDinst/U6354  ( .DIN1(\IDinst/RegFile[25][3] ), .DIN2(n1102), 
        .Q(\IDinst/n6349 ) );
  nnd2s1 \IDinst/U6353  ( .DIN1(\IDinst/RegFile[24][3] ), .DIN2(n1040), 
        .Q(\IDinst/n6348 ) );
  nnd2s1 \IDinst/U6352  ( .DIN1(\IDinst/n6346 ), .DIN2(\IDinst/n6345 ), 
        .Q(\IDinst/n6347 ) );
  nnd2s1 \IDinst/U6351  ( .DIN1(\IDinst/n6344 ), .DIN2(n1196), 
        .Q(\IDinst/n6346 ) );
  nnd2s1 \IDinst/U6350  ( .DIN1(\IDinst/n6335 ), .DIN2(n1189), 
        .Q(\IDinst/n6345 ) );
  nnd2s1 \IDinst/U6349  ( .DIN1(\IDinst/n6343 ), .DIN2(\IDinst/n6342 ), 
        .Q(\IDinst/n6344 ) );
  nnd2s1 \IDinst/U6348  ( .DIN1(\IDinst/n6341 ), .DIN2(n1169), 
        .Q(\IDinst/n6343 ) );
  nnd2s1 \IDinst/U6347  ( .DIN1(\IDinst/n6338 ), .DIN2(n1141), 
        .Q(\IDinst/n6342 ) );
  nnd2s1 \IDinst/U6346  ( .DIN1(\IDinst/n6340 ), .DIN2(\IDinst/n6339 ), 
        .Q(\IDinst/n6341 ) );
  nnd2s1 \IDinst/U6345  ( .DIN1(\IDinst/RegFile[23][3] ), .DIN2(n1102), 
        .Q(\IDinst/n6340 ) );
  nnd2s1 \IDinst/U6344  ( .DIN1(\IDinst/RegFile[22][3] ), .DIN2(n1039), 
        .Q(\IDinst/n6339 ) );
  nnd2s1 \IDinst/U6343  ( .DIN1(\IDinst/n6337 ), .DIN2(\IDinst/n6336 ), 
        .Q(\IDinst/n6338 ) );
  nnd2s1 \IDinst/U6342  ( .DIN1(\IDinst/RegFile[21][3] ), .DIN2(n1103), 
        .Q(\IDinst/n6337 ) );
  nnd2s1 \IDinst/U6341  ( .DIN1(\IDinst/RegFile[20][3] ), .DIN2(n1039), 
        .Q(\IDinst/n6336 ) );
  nnd2s1 \IDinst/U6340  ( .DIN1(\IDinst/n6334 ), .DIN2(\IDinst/n6333 ), 
        .Q(\IDinst/n6335 ) );
  nnd2s1 \IDinst/U6339  ( .DIN1(\IDinst/n6332 ), .DIN2(n1169), 
        .Q(\IDinst/n6334 ) );
  nnd2s1 \IDinst/U6338  ( .DIN1(\IDinst/n6329 ), .DIN2(n1141), 
        .Q(\IDinst/n6333 ) );
  nnd2s1 \IDinst/U6337  ( .DIN1(\IDinst/n6331 ), .DIN2(\IDinst/n6330 ), 
        .Q(\IDinst/n6332 ) );
  nnd2s1 \IDinst/U6336  ( .DIN1(\IDinst/RegFile[19][3] ), .DIN2(n1103), 
        .Q(\IDinst/n6331 ) );
  nnd2s1 \IDinst/U6335  ( .DIN1(\IDinst/RegFile[18][3] ), .DIN2(n1039), 
        .Q(\IDinst/n6330 ) );
  nnd2s1 \IDinst/U6334  ( .DIN1(\IDinst/n6328 ), .DIN2(\IDinst/n6327 ), 
        .Q(\IDinst/n6329 ) );
  nnd2s1 \IDinst/U6333  ( .DIN1(\IDinst/RegFile[17][3] ), .DIN2(n1103), 
        .Q(\IDinst/n6328 ) );
  nnd2s1 \IDinst/U6332  ( .DIN1(\IDinst/RegFile[16][3] ), .DIN2(n1039), 
        .Q(\IDinst/n6327 ) );
  nnd2s1 \IDinst/U6331  ( .DIN1(\IDinst/n6325 ), .DIN2(\IDinst/n6324 ), 
        .Q(\IDinst/n6326 ) );
  nnd2s1 \IDinst/U6330  ( .DIN1(\IDinst/n6323 ), .DIN2(n644), 
        .Q(\IDinst/n6325 ) );
  nnd2s1 \IDinst/U6329  ( .DIN1(\IDinst/n6302 ), .DIN2(n673), 
        .Q(\IDinst/n6324 ) );
  nnd2s1 \IDinst/U6328  ( .DIN1(\IDinst/n6322 ), .DIN2(\IDinst/n6321 ), 
        .Q(\IDinst/n6323 ) );
  nnd2s1 \IDinst/U6327  ( .DIN1(\IDinst/n6320 ), .DIN2(n1196), 
        .Q(\IDinst/n6322 ) );
  nnd2s1 \IDinst/U6326  ( .DIN1(\IDinst/n6311 ), .DIN2(n1188), 
        .Q(\IDinst/n6321 ) );
  nnd2s1 \IDinst/U6325  ( .DIN1(\IDinst/n6319 ), .DIN2(\IDinst/n6318 ), 
        .Q(\IDinst/n6320 ) );
  nnd2s1 \IDinst/U6324  ( .DIN1(\IDinst/n6317 ), .DIN2(n1169), 
        .Q(\IDinst/n6319 ) );
  nnd2s1 \IDinst/U6323  ( .DIN1(\IDinst/n6314 ), .DIN2(n1141), 
        .Q(\IDinst/n6318 ) );
  nnd2s1 \IDinst/U6322  ( .DIN1(\IDinst/n6316 ), .DIN2(\IDinst/n6315 ), 
        .Q(\IDinst/n6317 ) );
  nnd2s1 \IDinst/U6321  ( .DIN1(\IDinst/RegFile[15][3] ), .DIN2(n1103), 
        .Q(\IDinst/n6316 ) );
  nnd2s1 \IDinst/U6320  ( .DIN1(\IDinst/RegFile[14][3] ), .DIN2(n1039), 
        .Q(\IDinst/n6315 ) );
  nnd2s1 \IDinst/U6319  ( .DIN1(\IDinst/n6313 ), .DIN2(\IDinst/n6312 ), 
        .Q(\IDinst/n6314 ) );
  nnd2s1 \IDinst/U6318  ( .DIN1(\IDinst/RegFile[13][3] ), .DIN2(n1103), 
        .Q(\IDinst/n6313 ) );
  nnd2s1 \IDinst/U6317  ( .DIN1(\IDinst/RegFile[12][3] ), .DIN2(n1039), 
        .Q(\IDinst/n6312 ) );
  nnd2s1 \IDinst/U6316  ( .DIN1(\IDinst/n6310 ), .DIN2(\IDinst/n6309 ), 
        .Q(\IDinst/n6311 ) );
  nnd2s1 \IDinst/U6315  ( .DIN1(\IDinst/n6308 ), .DIN2(n1169), 
        .Q(\IDinst/n6310 ) );
  nnd2s1 \IDinst/U6314  ( .DIN1(\IDinst/n6305 ), .DIN2(n1141), 
        .Q(\IDinst/n6309 ) );
  nnd2s1 \IDinst/U6313  ( .DIN1(\IDinst/n6307 ), .DIN2(\IDinst/n6306 ), 
        .Q(\IDinst/n6308 ) );
  nnd2s1 \IDinst/U6312  ( .DIN1(\IDinst/RegFile[11][3] ), .DIN2(n1103), 
        .Q(\IDinst/n6307 ) );
  nnd2s1 \IDinst/U6311  ( .DIN1(\IDinst/RegFile[10][3] ), .DIN2(n1039), 
        .Q(\IDinst/n6306 ) );
  nnd2s1 \IDinst/U6310  ( .DIN1(\IDinst/n6304 ), .DIN2(\IDinst/n6303 ), 
        .Q(\IDinst/n6305 ) );
  nnd2s1 \IDinst/U6309  ( .DIN1(\IDinst/RegFile[9][3] ), .DIN2(n1103), 
        .Q(\IDinst/n6304 ) );
  nnd2s1 \IDinst/U6308  ( .DIN1(\IDinst/RegFile[8][3] ), .DIN2(n1039), 
        .Q(\IDinst/n6303 ) );
  nnd2s1 \IDinst/U6307  ( .DIN1(\IDinst/n6301 ), .DIN2(\IDinst/n6300 ), 
        .Q(\IDinst/n6302 ) );
  nnd2s1 \IDinst/U6306  ( .DIN1(\IDinst/n6299 ), .DIN2(n1196), 
        .Q(\IDinst/n6301 ) );
  nnd2s1 \IDinst/U6305  ( .DIN1(\IDinst/n6290 ), .DIN2(n1187), 
        .Q(\IDinst/n6300 ) );
  nnd2s1 \IDinst/U6304  ( .DIN1(\IDinst/n6298 ), .DIN2(\IDinst/n6297 ), 
        .Q(\IDinst/n6299 ) );
  nnd2s1 \IDinst/U6303  ( .DIN1(\IDinst/n6296 ), .DIN2(n1168), 
        .Q(\IDinst/n6298 ) );
  nnd2s1 \IDinst/U6302  ( .DIN1(\IDinst/n6293 ), .DIN2(n1141), 
        .Q(\IDinst/n6297 ) );
  nnd2s1 \IDinst/U6301  ( .DIN1(\IDinst/n6295 ), .DIN2(\IDinst/n6294 ), 
        .Q(\IDinst/n6296 ) );
  nnd2s1 \IDinst/U6300  ( .DIN1(\IDinst/RegFile[7][3] ), .DIN2(n1103), 
        .Q(\IDinst/n6295 ) );
  nnd2s1 \IDinst/U6299  ( .DIN1(\IDinst/RegFile[6][3] ), .DIN2(n1039), 
        .Q(\IDinst/n6294 ) );
  nnd2s1 \IDinst/U6298  ( .DIN1(\IDinst/n6292 ), .DIN2(\IDinst/n6291 ), 
        .Q(\IDinst/n6293 ) );
  nnd2s1 \IDinst/U6297  ( .DIN1(\IDinst/RegFile[5][3] ), .DIN2(n1104), 
        .Q(\IDinst/n6292 ) );
  nnd2s1 \IDinst/U6296  ( .DIN1(\IDinst/RegFile[4][3] ), .DIN2(n1039), 
        .Q(\IDinst/n6291 ) );
  nnd2s1 \IDinst/U6295  ( .DIN1(\IDinst/n6289 ), .DIN2(\IDinst/n6288 ), 
        .Q(\IDinst/n6290 ) );
  nnd2s1 \IDinst/U6294  ( .DIN1(\IDinst/n6287 ), .DIN2(n1168), 
        .Q(\IDinst/n6289 ) );
  nnd2s1 \IDinst/U6293  ( .DIN1(\IDinst/n6284 ), .DIN2(n1141), 
        .Q(\IDinst/n6288 ) );
  nnd2s1 \IDinst/U6292  ( .DIN1(\IDinst/n6286 ), .DIN2(\IDinst/n6285 ), 
        .Q(\IDinst/n6287 ) );
  nnd2s1 \IDinst/U6291  ( .DIN1(\IDinst/RegFile[3][3] ), .DIN2(n1104), 
        .Q(\IDinst/n6286 ) );
  nnd2s1 \IDinst/U6290  ( .DIN1(\IDinst/RegFile[2][3] ), .DIN2(n1039), 
        .Q(\IDinst/n6285 ) );
  nnd2s1 \IDinst/U6289  ( .DIN1(\IDinst/n6283 ), .DIN2(\IDinst/n6282 ), 
        .Q(\IDinst/n6284 ) );
  nnd2s1 \IDinst/U6288  ( .DIN1(\IDinst/RegFile[1][3] ), .DIN2(n1104), 
        .Q(\IDinst/n6283 ) );
  nnd2s1 \IDinst/U6287  ( .DIN1(\IDinst/RegFile[0][3] ), .DIN2(n1039), 
        .Q(\IDinst/n6282 ) );
  nnd2s1 \IDinst/U6286  ( .DIN1(\IDinst/n6281 ), .DIN2(\IDinst/N43 ), 
        .Q(\IDinst/n5952 ) );
  nnd2s1 \IDinst/U6285  ( .DIN1(\IDinst/n6236 ), .DIN2(n636), 
        .Q(\IDinst/n5953 ) );
  nnd2s1 \IDinst/U6284  ( .DIN1(\IDinst/n6280 ), .DIN2(\IDinst/n6279 ), 
        .Q(\IDinst/n6281 ) );
  nnd2s1 \IDinst/U6283  ( .DIN1(\IDinst/n6278 ), .DIN2(n643), 
        .Q(\IDinst/n6280 ) );
  nnd2s1 \IDinst/U6282  ( .DIN1(\IDinst/n6257 ), .DIN2(n671), 
        .Q(\IDinst/n6279 ) );
  nnd2s1 \IDinst/U6281  ( .DIN1(\IDinst/n6277 ), .DIN2(\IDinst/n6276 ), 
        .Q(\IDinst/n6278 ) );
  nnd2s1 \IDinst/U6280  ( .DIN1(\IDinst/n6275 ), .DIN2(n1196), 
        .Q(\IDinst/n6277 ) );
  nnd2s1 \IDinst/U6279  ( .DIN1(\IDinst/n6266 ), .DIN2(n1186), 
        .Q(\IDinst/n6276 ) );
  nnd2s1 \IDinst/U6278  ( .DIN1(\IDinst/n6274 ), .DIN2(\IDinst/n6273 ), 
        .Q(\IDinst/n6275 ) );
  nnd2s1 \IDinst/U6277  ( .DIN1(\IDinst/n6272 ), .DIN2(n1168), 
        .Q(\IDinst/n6274 ) );
  nnd2s1 \IDinst/U6276  ( .DIN1(\IDinst/n6269 ), .DIN2(n1141), 
        .Q(\IDinst/n6273 ) );
  nnd2s1 \IDinst/U6275  ( .DIN1(\IDinst/n6271 ), .DIN2(\IDinst/n6270 ), 
        .Q(\IDinst/n6272 ) );
  nnd2s1 \IDinst/U6274  ( .DIN1(\IDinst/RegFile[31][2] ), .DIN2(n1104), 
        .Q(\IDinst/n6271 ) );
  nnd2s1 \IDinst/U6273  ( .DIN1(\IDinst/RegFile[30][2] ), .DIN2(n1039), 
        .Q(\IDinst/n6270 ) );
  nnd2s1 \IDinst/U6272  ( .DIN1(\IDinst/n6268 ), .DIN2(\IDinst/n6267 ), 
        .Q(\IDinst/n6269 ) );
  nnd2s1 \IDinst/U6271  ( .DIN1(\IDinst/RegFile[29][2] ), .DIN2(n1104), 
        .Q(\IDinst/n6268 ) );
  nnd2s1 \IDinst/U6270  ( .DIN1(\IDinst/RegFile[28][2] ), .DIN2(n1038), 
        .Q(\IDinst/n6267 ) );
  nnd2s1 \IDinst/U6269  ( .DIN1(\IDinst/n6265 ), .DIN2(\IDinst/n6264 ), 
        .Q(\IDinst/n6266 ) );
  nnd2s1 \IDinst/U6268  ( .DIN1(\IDinst/n6263 ), .DIN2(n1168), 
        .Q(\IDinst/n6265 ) );
  nnd2s1 \IDinst/U6267  ( .DIN1(\IDinst/n6260 ), .DIN2(n1141), 
        .Q(\IDinst/n6264 ) );
  nnd2s1 \IDinst/U6266  ( .DIN1(\IDinst/n6262 ), .DIN2(\IDinst/n6261 ), 
        .Q(\IDinst/n6263 ) );
  nnd2s1 \IDinst/U6265  ( .DIN1(\IDinst/RegFile[27][2] ), .DIN2(n1104), 
        .Q(\IDinst/n6262 ) );
  nnd2s1 \IDinst/U6264  ( .DIN1(\IDinst/RegFile[26][2] ), .DIN2(n1038), 
        .Q(\IDinst/n6261 ) );
  nnd2s1 \IDinst/U6263  ( .DIN1(\IDinst/n6259 ), .DIN2(\IDinst/n6258 ), 
        .Q(\IDinst/n6260 ) );
  nnd2s1 \IDinst/U6262  ( .DIN1(\IDinst/RegFile[25][2] ), .DIN2(n1104), 
        .Q(\IDinst/n6259 ) );
  nnd2s1 \IDinst/U6261  ( .DIN1(\IDinst/RegFile[24][2] ), .DIN2(n1038), 
        .Q(\IDinst/n6258 ) );
  nnd2s1 \IDinst/U6260  ( .DIN1(\IDinst/n6256 ), .DIN2(\IDinst/n6255 ), 
        .Q(\IDinst/n6257 ) );
  nnd2s1 \IDinst/U6259  ( .DIN1(\IDinst/n6254 ), .DIN2(n1196), 
        .Q(\IDinst/n6256 ) );
  nnd2s1 \IDinst/U6258  ( .DIN1(\IDinst/n6245 ), .DIN2(n1185), 
        .Q(\IDinst/n6255 ) );
  nnd2s1 \IDinst/U6257  ( .DIN1(\IDinst/n6253 ), .DIN2(\IDinst/n6252 ), 
        .Q(\IDinst/n6254 ) );
  nnd2s1 \IDinst/U6256  ( .DIN1(\IDinst/n6251 ), .DIN2(n1168), 
        .Q(\IDinst/n6253 ) );
  nnd2s1 \IDinst/U6255  ( .DIN1(\IDinst/n6248 ), .DIN2(n1142), 
        .Q(\IDinst/n6252 ) );
  nnd2s1 \IDinst/U6254  ( .DIN1(\IDinst/n6250 ), .DIN2(\IDinst/n6249 ), 
        .Q(\IDinst/n6251 ) );
  nnd2s1 \IDinst/U6253  ( .DIN1(\IDinst/RegFile[23][2] ), .DIN2(n1104), 
        .Q(\IDinst/n6250 ) );
  nnd2s1 \IDinst/U6252  ( .DIN1(\IDinst/RegFile[22][2] ), .DIN2(n1038), 
        .Q(\IDinst/n6249 ) );
  nnd2s1 \IDinst/U6251  ( .DIN1(\IDinst/n6247 ), .DIN2(\IDinst/n6246 ), 
        .Q(\IDinst/n6248 ) );
  nnd2s1 \IDinst/U6250  ( .DIN1(\IDinst/RegFile[21][2] ), .DIN2(n1104), 
        .Q(\IDinst/n6247 ) );
  nnd2s1 \IDinst/U6249  ( .DIN1(\IDinst/RegFile[20][2] ), .DIN2(n1038), 
        .Q(\IDinst/n6246 ) );
  nnd2s1 \IDinst/U6248  ( .DIN1(\IDinst/n6244 ), .DIN2(\IDinst/n6243 ), 
        .Q(\IDinst/n6245 ) );
  nnd2s1 \IDinst/U6247  ( .DIN1(\IDinst/n6242 ), .DIN2(n1168), 
        .Q(\IDinst/n6244 ) );
  nnd2s1 \IDinst/U6246  ( .DIN1(\IDinst/n6239 ), .DIN2(n1142), 
        .Q(\IDinst/n6243 ) );
  nnd2s1 \IDinst/U6245  ( .DIN1(\IDinst/n6241 ), .DIN2(\IDinst/n6240 ), 
        .Q(\IDinst/n6242 ) );
  nnd2s1 \IDinst/U6244  ( .DIN1(\IDinst/RegFile[19][2] ), .DIN2(n1105), 
        .Q(\IDinst/n6241 ) );
  nnd2s1 \IDinst/U6243  ( .DIN1(\IDinst/RegFile[18][2] ), .DIN2(n1038), 
        .Q(\IDinst/n6240 ) );
  nnd2s1 \IDinst/U6242  ( .DIN1(\IDinst/n6238 ), .DIN2(\IDinst/n6237 ), 
        .Q(\IDinst/n6239 ) );
  nnd2s1 \IDinst/U6241  ( .DIN1(\IDinst/RegFile[17][2] ), .DIN2(n1105), 
        .Q(\IDinst/n6238 ) );
  nnd2s1 \IDinst/U6240  ( .DIN1(\IDinst/RegFile[16][2] ), .DIN2(n1038), 
        .Q(\IDinst/n6237 ) );
  nnd2s1 \IDinst/U6239  ( .DIN1(\IDinst/n6235 ), .DIN2(\IDinst/n6234 ), 
        .Q(\IDinst/n6236 ) );
  nnd2s1 \IDinst/U6238  ( .DIN1(\IDinst/n6233 ), .DIN2(n642), 
        .Q(\IDinst/n6235 ) );
  nnd2s1 \IDinst/U6237  ( .DIN1(\IDinst/n6212 ), .DIN2(n672), 
        .Q(\IDinst/n6234 ) );
  nnd2s1 \IDinst/U6236  ( .DIN1(\IDinst/n6232 ), .DIN2(\IDinst/n6231 ), 
        .Q(\IDinst/n6233 ) );
  nnd2s1 \IDinst/U6235  ( .DIN1(\IDinst/n6230 ), .DIN2(n1197), 
        .Q(\IDinst/n6232 ) );
  nnd2s1 \IDinst/U6234  ( .DIN1(\IDinst/n6221 ), .DIN2(n1184), 
        .Q(\IDinst/n6231 ) );
  nnd2s1 \IDinst/U6233  ( .DIN1(\IDinst/n6229 ), .DIN2(\IDinst/n6228 ), 
        .Q(\IDinst/n6230 ) );
  nnd2s1 \IDinst/U6232  ( .DIN1(\IDinst/n6227 ), .DIN2(n1168), 
        .Q(\IDinst/n6229 ) );
  nnd2s1 \IDinst/U6231  ( .DIN1(\IDinst/n6224 ), .DIN2(n1142), 
        .Q(\IDinst/n6228 ) );
  nnd2s1 \IDinst/U6230  ( .DIN1(\IDinst/n6226 ), .DIN2(\IDinst/n6225 ), 
        .Q(\IDinst/n6227 ) );
  nnd2s1 \IDinst/U6229  ( .DIN1(\IDinst/RegFile[15][2] ), .DIN2(n1105), 
        .Q(\IDinst/n6226 ) );
  nnd2s1 \IDinst/U6228  ( .DIN1(\IDinst/RegFile[14][2] ), .DIN2(n1038), 
        .Q(\IDinst/n6225 ) );
  nnd2s1 \IDinst/U6227  ( .DIN1(\IDinst/n6223 ), .DIN2(\IDinst/n6222 ), 
        .Q(\IDinst/n6224 ) );
  nnd2s1 \IDinst/U6226  ( .DIN1(\IDinst/RegFile[13][2] ), .DIN2(n1105), 
        .Q(\IDinst/n6223 ) );
  nnd2s1 \IDinst/U6225  ( .DIN1(\IDinst/RegFile[12][2] ), .DIN2(n1038), 
        .Q(\IDinst/n6222 ) );
  nnd2s1 \IDinst/U6224  ( .DIN1(\IDinst/n6220 ), .DIN2(\IDinst/n6219 ), 
        .Q(\IDinst/n6221 ) );
  nnd2s1 \IDinst/U6223  ( .DIN1(\IDinst/n6218 ), .DIN2(n1168), 
        .Q(\IDinst/n6220 ) );
  nnd2s1 \IDinst/U6222  ( .DIN1(\IDinst/n6215 ), .DIN2(n1142), 
        .Q(\IDinst/n6219 ) );
  nnd2s1 \IDinst/U6221  ( .DIN1(\IDinst/n6217 ), .DIN2(\IDinst/n6216 ), 
        .Q(\IDinst/n6218 ) );
  nnd2s1 \IDinst/U6220  ( .DIN1(\IDinst/RegFile[11][2] ), .DIN2(n1105), 
        .Q(\IDinst/n6217 ) );
  nnd2s1 \IDinst/U6219  ( .DIN1(\IDinst/RegFile[10][2] ), .DIN2(n1038), 
        .Q(\IDinst/n6216 ) );
  nnd2s1 \IDinst/U6218  ( .DIN1(\IDinst/n6214 ), .DIN2(\IDinst/n6213 ), 
        .Q(\IDinst/n6215 ) );
  nnd2s1 \IDinst/U6217  ( .DIN1(\IDinst/RegFile[9][2] ), .DIN2(n1105), 
        .Q(\IDinst/n6214 ) );
  nnd2s1 \IDinst/U6216  ( .DIN1(\IDinst/RegFile[8][2] ), .DIN2(n1038), 
        .Q(\IDinst/n6213 ) );
  nnd2s1 \IDinst/U6215  ( .DIN1(\IDinst/n6211 ), .DIN2(\IDinst/n6210 ), 
        .Q(\IDinst/n6212 ) );
  nnd2s1 \IDinst/U6214  ( .DIN1(\IDinst/n6209 ), .DIN2(n1197), 
        .Q(\IDinst/n6211 ) );
  nnd2s1 \IDinst/U6213  ( .DIN1(\IDinst/n6200 ), .DIN2(n1181), 
        .Q(\IDinst/n6210 ) );
  nnd2s1 \IDinst/U6212  ( .DIN1(\IDinst/n6208 ), .DIN2(\IDinst/n6207 ), 
        .Q(\IDinst/n6209 ) );
  nnd2s1 \IDinst/U6211  ( .DIN1(\IDinst/n6206 ), .DIN2(n1168), 
        .Q(\IDinst/n6208 ) );
  nnd2s1 \IDinst/U6210  ( .DIN1(\IDinst/n6203 ), .DIN2(n1142), 
        .Q(\IDinst/n6207 ) );
  nnd2s1 \IDinst/U6209  ( .DIN1(\IDinst/n6205 ), .DIN2(\IDinst/n6204 ), 
        .Q(\IDinst/n6206 ) );
  nnd2s1 \IDinst/U6208  ( .DIN1(\IDinst/RegFile[7][2] ), .DIN2(n1105), 
        .Q(\IDinst/n6205 ) );
  nnd2s1 \IDinst/U6207  ( .DIN1(\IDinst/RegFile[6][2] ), .DIN2(n1038), 
        .Q(\IDinst/n6204 ) );
  nnd2s1 \IDinst/U6206  ( .DIN1(\IDinst/n6202 ), .DIN2(\IDinst/n6201 ), 
        .Q(\IDinst/n6203 ) );
  nnd2s1 \IDinst/U6205  ( .DIN1(\IDinst/RegFile[5][2] ), .DIN2(n1105), 
        .Q(\IDinst/n6202 ) );
  nnd2s1 \IDinst/U6204  ( .DIN1(\IDinst/RegFile[4][2] ), .DIN2(n1038), 
        .Q(\IDinst/n6201 ) );
  nnd2s1 \IDinst/U6203  ( .DIN1(\IDinst/n6199 ), .DIN2(\IDinst/n6198 ), 
        .Q(\IDinst/n6200 ) );
  nnd2s1 \IDinst/U6202  ( .DIN1(\IDinst/n6197 ), .DIN2(n1167), 
        .Q(\IDinst/n6199 ) );
  nnd2s1 \IDinst/U6201  ( .DIN1(\IDinst/n6194 ), .DIN2(n1142), 
        .Q(\IDinst/n6198 ) );
  nnd2s1 \IDinst/U6200  ( .DIN1(\IDinst/n6196 ), .DIN2(\IDinst/n6195 ), 
        .Q(\IDinst/n6197 ) );
  nnd2s1 \IDinst/U6199  ( .DIN1(\IDinst/RegFile[3][2] ), .DIN2(n1105), 
        .Q(\IDinst/n6196 ) );
  nnd2s1 \IDinst/U6198  ( .DIN1(\IDinst/RegFile[2][2] ), .DIN2(n1037), 
        .Q(\IDinst/n6195 ) );
  nnd2s1 \IDinst/U6197  ( .DIN1(\IDinst/n6193 ), .DIN2(\IDinst/n6192 ), 
        .Q(\IDinst/n6194 ) );
  nnd2s1 \IDinst/U6196  ( .DIN1(\IDinst/RegFile[1][2] ), .DIN2(n1106), 
        .Q(\IDinst/n6193 ) );
  nnd2s1 \IDinst/U6195  ( .DIN1(\IDinst/RegFile[0][2] ), .DIN2(n1037), 
        .Q(\IDinst/n6192 ) );
  nnd2s1 \IDinst/U6194  ( .DIN1(\IDinst/n6191 ), .DIN2(n539), 
        .Q(\IDinst/n5950 ) );
  nnd2s1 \IDinst/U6193  ( .DIN1(\IDinst/n6146 ), .DIN2(n635), 
        .Q(\IDinst/n5951 ) );
  nnd2s1 \IDinst/U6192  ( .DIN1(\IDinst/n6190 ), .DIN2(\IDinst/n6189 ), 
        .Q(\IDinst/n6191 ) );
  nnd2s1 \IDinst/U6191  ( .DIN1(\IDinst/n6188 ), .DIN2(n644), 
        .Q(\IDinst/n6190 ) );
  nnd2s1 \IDinst/U6190  ( .DIN1(\IDinst/n6167 ), .DIN2(n670), 
        .Q(\IDinst/n6189 ) );
  nnd2s1 \IDinst/U6189  ( .DIN1(\IDinst/n6187 ), .DIN2(\IDinst/n6186 ), 
        .Q(\IDinst/n6188 ) );
  nnd2s1 \IDinst/U6188  ( .DIN1(\IDinst/n6185 ), .DIN2(n1197), 
        .Q(\IDinst/n6187 ) );
  nnd2s1 \IDinst/U6187  ( .DIN1(\IDinst/n6176 ), .DIN2(n1183), 
        .Q(\IDinst/n6186 ) );
  nnd2s1 \IDinst/U6186  ( .DIN1(\IDinst/n6184 ), .DIN2(\IDinst/n6183 ), 
        .Q(\IDinst/n6185 ) );
  nnd2s1 \IDinst/U6185  ( .DIN1(\IDinst/n6182 ), .DIN2(n1167), 
        .Q(\IDinst/n6184 ) );
  nnd2s1 \IDinst/U6184  ( .DIN1(\IDinst/n6179 ), .DIN2(n1142), 
        .Q(\IDinst/n6183 ) );
  nnd2s1 \IDinst/U6183  ( .DIN1(\IDinst/n6181 ), .DIN2(\IDinst/n6180 ), 
        .Q(\IDinst/n6182 ) );
  nnd2s1 \IDinst/U6182  ( .DIN1(\IDinst/RegFile[31][1] ), .DIN2(n1106), 
        .Q(\IDinst/n6181 ) );
  nnd2s1 \IDinst/U6181  ( .DIN1(\IDinst/RegFile[30][1] ), .DIN2(n1037), 
        .Q(\IDinst/n6180 ) );
  nnd2s1 \IDinst/U6180  ( .DIN1(\IDinst/n6178 ), .DIN2(\IDinst/n6177 ), 
        .Q(\IDinst/n6179 ) );
  nnd2s1 \IDinst/U6179  ( .DIN1(\IDinst/RegFile[29][1] ), .DIN2(n1106), 
        .Q(\IDinst/n6178 ) );
  nnd2s1 \IDinst/U6178  ( .DIN1(\IDinst/RegFile[28][1] ), .DIN2(n1037), 
        .Q(\IDinst/n6177 ) );
  nnd2s1 \IDinst/U6177  ( .DIN1(\IDinst/n6175 ), .DIN2(\IDinst/n6174 ), 
        .Q(\IDinst/n6176 ) );
  nnd2s1 \IDinst/U6176  ( .DIN1(\IDinst/n6173 ), .DIN2(n1167), 
        .Q(\IDinst/n6175 ) );
  nnd2s1 \IDinst/U6175  ( .DIN1(\IDinst/n6170 ), .DIN2(n1142), 
        .Q(\IDinst/n6174 ) );
  nnd2s1 \IDinst/U6174  ( .DIN1(\IDinst/n6172 ), .DIN2(\IDinst/n6171 ), 
        .Q(\IDinst/n6173 ) );
  nnd2s1 \IDinst/U6173  ( .DIN1(\IDinst/RegFile[27][1] ), .DIN2(n1106), 
        .Q(\IDinst/n6172 ) );
  nnd2s1 \IDinst/U6172  ( .DIN1(\IDinst/RegFile[26][1] ), .DIN2(n1037), 
        .Q(\IDinst/n6171 ) );
  nnd2s1 \IDinst/U6171  ( .DIN1(\IDinst/n6169 ), .DIN2(\IDinst/n6168 ), 
        .Q(\IDinst/n6170 ) );
  nnd2s1 \IDinst/U6170  ( .DIN1(\IDinst/RegFile[25][1] ), .DIN2(n1106), 
        .Q(\IDinst/n6169 ) );
  nnd2s1 \IDinst/U6169  ( .DIN1(\IDinst/RegFile[24][1] ), .DIN2(n1037), 
        .Q(\IDinst/n6168 ) );
  nnd2s1 \IDinst/U6168  ( .DIN1(\IDinst/n6166 ), .DIN2(\IDinst/n6165 ), 
        .Q(\IDinst/n6167 ) );
  nnd2s1 \IDinst/U6167  ( .DIN1(\IDinst/n6164 ), .DIN2(n1197), 
        .Q(\IDinst/n6166 ) );
  nnd2s1 \IDinst/U6166  ( .DIN1(\IDinst/n6155 ), .DIN2(n1182), 
        .Q(\IDinst/n6165 ) );
  nnd2s1 \IDinst/U6165  ( .DIN1(\IDinst/n6163 ), .DIN2(\IDinst/n6162 ), 
        .Q(\IDinst/n6164 ) );
  nnd2s1 \IDinst/U6164  ( .DIN1(\IDinst/n6161 ), .DIN2(n1167), 
        .Q(\IDinst/n6163 ) );
  nnd2s1 \IDinst/U6163  ( .DIN1(\IDinst/n6158 ), .DIN2(n1142), 
        .Q(\IDinst/n6162 ) );
  nnd2s1 \IDinst/U6162  ( .DIN1(\IDinst/n6160 ), .DIN2(\IDinst/n6159 ), 
        .Q(\IDinst/n6161 ) );
  nnd2s1 \IDinst/U6161  ( .DIN1(\IDinst/RegFile[23][1] ), .DIN2(n1106), 
        .Q(\IDinst/n6160 ) );
  nnd2s1 \IDinst/U6160  ( .DIN1(\IDinst/RegFile[22][1] ), .DIN2(n1037), 
        .Q(\IDinst/n6159 ) );
  nnd2s1 \IDinst/U6159  ( .DIN1(\IDinst/n6157 ), .DIN2(\IDinst/n6156 ), 
        .Q(\IDinst/n6158 ) );
  nnd2s1 \IDinst/U6158  ( .DIN1(\IDinst/RegFile[21][1] ), .DIN2(n1106), 
        .Q(\IDinst/n6157 ) );
  nnd2s1 \IDinst/U6157  ( .DIN1(\IDinst/RegFile[20][1] ), .DIN2(n1037), 
        .Q(\IDinst/n6156 ) );
  nnd2s1 \IDinst/U6156  ( .DIN1(\IDinst/n6154 ), .DIN2(\IDinst/n6153 ), 
        .Q(\IDinst/n6155 ) );
  nnd2s1 \IDinst/U6155  ( .DIN1(\IDinst/n6152 ), .DIN2(n1167), 
        .Q(\IDinst/n6154 ) );
  nnd2s1 \IDinst/U6154  ( .DIN1(\IDinst/n6149 ), .DIN2(n1142), 
        .Q(\IDinst/n6153 ) );
  nnd2s1 \IDinst/U6153  ( .DIN1(\IDinst/n6151 ), .DIN2(\IDinst/n6150 ), 
        .Q(\IDinst/n6152 ) );
  nnd2s1 \IDinst/U6152  ( .DIN1(\IDinst/RegFile[19][1] ), .DIN2(n1106), 
        .Q(\IDinst/n6151 ) );
  nnd2s1 \IDinst/U6151  ( .DIN1(\IDinst/RegFile[18][1] ), .DIN2(n1037), 
        .Q(\IDinst/n6150 ) );
  nnd2s1 \IDinst/U6150  ( .DIN1(\IDinst/n6148 ), .DIN2(\IDinst/n6147 ), 
        .Q(\IDinst/n6149 ) );
  nnd2s1 \IDinst/U6149  ( .DIN1(\IDinst/RegFile[17][1] ), .DIN2(n1106), 
        .Q(\IDinst/n6148 ) );
  nnd2s1 \IDinst/U6148  ( .DIN1(\IDinst/RegFile[16][1] ), .DIN2(n1037), 
        .Q(\IDinst/n6147 ) );
  nnd2s1 \IDinst/U6147  ( .DIN1(\IDinst/n6145 ), .DIN2(\IDinst/n6144 ), 
        .Q(\IDinst/n6146 ) );
  nnd2s1 \IDinst/U6146  ( .DIN1(\IDinst/n6143 ), .DIN2(n643), 
        .Q(\IDinst/n6145 ) );
  nnd2s1 \IDinst/U6145  ( .DIN1(\IDinst/n6122 ), .DIN2(n673), 
        .Q(\IDinst/n6144 ) );
  nnd2s1 \IDinst/U6144  ( .DIN1(\IDinst/n6142 ), .DIN2(\IDinst/n6141 ), 
        .Q(\IDinst/n6143 ) );
  nnd2s1 \IDinst/U6143  ( .DIN1(\IDinst/n6140 ), .DIN2(n1197), 
        .Q(\IDinst/n6142 ) );
  nnd2s1 \IDinst/U6142  ( .DIN1(\IDinst/n6131 ), .DIN2(n1181), 
        .Q(\IDinst/n6141 ) );
  nnd2s1 \IDinst/U6141  ( .DIN1(\IDinst/n6139 ), .DIN2(\IDinst/n6138 ), 
        .Q(\IDinst/n6140 ) );
  nnd2s1 \IDinst/U6140  ( .DIN1(\IDinst/n6137 ), .DIN2(n1167), 
        .Q(\IDinst/n6139 ) );
  nnd2s1 \IDinst/U6139  ( .DIN1(\IDinst/n6134 ), .DIN2(n1142), 
        .Q(\IDinst/n6138 ) );
  nnd2s1 \IDinst/U6138  ( .DIN1(\IDinst/n6136 ), .DIN2(\IDinst/n6135 ), 
        .Q(\IDinst/n6137 ) );
  nnd2s1 \IDinst/U6137  ( .DIN1(\IDinst/RegFile[15][1] ), .DIN2(n1107), 
        .Q(\IDinst/n6136 ) );
  nnd2s1 \IDinst/U6136  ( .DIN1(\IDinst/RegFile[14][1] ), .DIN2(n1037), 
        .Q(\IDinst/n6135 ) );
  nnd2s1 \IDinst/U6135  ( .DIN1(\IDinst/n6133 ), .DIN2(\IDinst/n6132 ), 
        .Q(\IDinst/n6134 ) );
  nnd2s1 \IDinst/U6134  ( .DIN1(\IDinst/RegFile[13][1] ), .DIN2(n1107), 
        .Q(\IDinst/n6133 ) );
  nnd2s1 \IDinst/U6133  ( .DIN1(\IDinst/RegFile[12][1] ), .DIN2(n1037), 
        .Q(\IDinst/n6132 ) );
  nnd2s1 \IDinst/U6132  ( .DIN1(\IDinst/n6130 ), .DIN2(\IDinst/n6129 ), 
        .Q(\IDinst/n6131 ) );
  nnd2s1 \IDinst/U6131  ( .DIN1(\IDinst/n6128 ), .DIN2(n1167), 
        .Q(\IDinst/n6130 ) );
  nnd2s1 \IDinst/U6130  ( .DIN1(\IDinst/n6125 ), .DIN2(n1142), 
        .Q(\IDinst/n6129 ) );
  nnd2s1 \IDinst/U6129  ( .DIN1(\IDinst/n6127 ), .DIN2(\IDinst/n6126 ), 
        .Q(\IDinst/n6128 ) );
  nnd2s1 \IDinst/U6128  ( .DIN1(\IDinst/RegFile[11][1] ), .DIN2(n1107), 
        .Q(\IDinst/n6127 ) );
  nnd2s1 \IDinst/U6127  ( .DIN1(\IDinst/RegFile[10][1] ), .DIN2(n1037), 
        .Q(\IDinst/n6126 ) );
  nnd2s1 \IDinst/U6126  ( .DIN1(\IDinst/n6124 ), .DIN2(\IDinst/n6123 ), 
        .Q(\IDinst/n6125 ) );
  nnd2s1 \IDinst/U6125  ( .DIN1(\IDinst/RegFile[9][1] ), .DIN2(n1107), 
        .Q(\IDinst/n6124 ) );
  nnd2s1 \IDinst/U6124  ( .DIN1(\IDinst/RegFile[8][1] ), .DIN2(n1036), 
        .Q(\IDinst/n6123 ) );
  nnd2s1 \IDinst/U6123  ( .DIN1(\IDinst/n6121 ), .DIN2(\IDinst/n6120 ), 
        .Q(\IDinst/n6122 ) );
  nnd2s1 \IDinst/U6122  ( .DIN1(\IDinst/n6119 ), .DIN2(n1197), 
        .Q(\IDinst/n6121 ) );
  nnd2s1 \IDinst/U6121  ( .DIN1(\IDinst/n6110 ), .DIN2(n1181), 
        .Q(\IDinst/n6120 ) );
  nnd2s1 \IDinst/U6120  ( .DIN1(\IDinst/n6118 ), .DIN2(\IDinst/n6117 ), 
        .Q(\IDinst/n6119 ) );
  nnd2s1 \IDinst/U6119  ( .DIN1(\IDinst/n6116 ), .DIN2(n1167), 
        .Q(\IDinst/n6118 ) );
  nnd2s1 \IDinst/U6118  ( .DIN1(\IDinst/n6113 ), .DIN2(n1142), 
        .Q(\IDinst/n6117 ) );
  nnd2s1 \IDinst/U6117  ( .DIN1(\IDinst/n6115 ), .DIN2(\IDinst/n6114 ), 
        .Q(\IDinst/n6116 ) );
  nnd2s1 \IDinst/U6116  ( .DIN1(\IDinst/RegFile[7][1] ), .DIN2(n1107), 
        .Q(\IDinst/n6115 ) );
  nnd2s1 \IDinst/U6115  ( .DIN1(\IDinst/RegFile[6][1] ), .DIN2(n1036), 
        .Q(\IDinst/n6114 ) );
  nnd2s1 \IDinst/U6114  ( .DIN1(\IDinst/n6112 ), .DIN2(\IDinst/n6111 ), 
        .Q(\IDinst/n6113 ) );
  nnd2s1 \IDinst/U6113  ( .DIN1(\IDinst/RegFile[5][1] ), .DIN2(n1107), 
        .Q(\IDinst/n6112 ) );
  nnd2s1 \IDinst/U6112  ( .DIN1(\IDinst/RegFile[4][1] ), .DIN2(n1036), 
        .Q(\IDinst/n6111 ) );
  nnd2s1 \IDinst/U6111  ( .DIN1(\IDinst/n6109 ), .DIN2(\IDinst/n6108 ), 
        .Q(\IDinst/n6110 ) );
  nnd2s1 \IDinst/U6110  ( .DIN1(\IDinst/n6107 ), .DIN2(n1167), 
        .Q(\IDinst/n6109 ) );
  nnd2s1 \IDinst/U6109  ( .DIN1(\IDinst/n6104 ), .DIN2(n1143), 
        .Q(\IDinst/n6108 ) );
  nnd2s1 \IDinst/U6108  ( .DIN1(\IDinst/n6106 ), .DIN2(\IDinst/n6105 ), 
        .Q(\IDinst/n6107 ) );
  nnd2s1 \IDinst/U6107  ( .DIN1(\IDinst/RegFile[3][1] ), .DIN2(n1107), 
        .Q(\IDinst/n6106 ) );
  nnd2s1 \IDinst/U6106  ( .DIN1(\IDinst/RegFile[2][1] ), .DIN2(n1036), 
        .Q(\IDinst/n6105 ) );
  nnd2s1 \IDinst/U6105  ( .DIN1(\IDinst/n6103 ), .DIN2(\IDinst/n6102 ), 
        .Q(\IDinst/n6104 ) );
  nnd2s1 \IDinst/U6104  ( .DIN1(\IDinst/RegFile[1][1] ), .DIN2(n1107), 
        .Q(\IDinst/n6103 ) );
  nnd2s1 \IDinst/U6103  ( .DIN1(\IDinst/RegFile[0][1] ), .DIN2(n1036), 
        .Q(\IDinst/n6102 ) );
  nnd2s1 \IDinst/U6102  ( .DIN1(n539), .DIN2(\IDinst/n6101 ), 
        .Q(\IDinst/n5948 ) );
  nnd2s1 \IDinst/U6101  ( .DIN1(\IDinst/n6056 ), .DIN2(n636), 
        .Q(\IDinst/n5949 ) );
  nnd2s1 \IDinst/U6100  ( .DIN1(\IDinst/n6100 ), .DIN2(\IDinst/n6099 ), 
        .Q(\IDinst/n6101 ) );
  nnd2s1 \IDinst/U6099  ( .DIN1(\IDinst/n6098 ), .DIN2(n642), 
        .Q(\IDinst/n6100 ) );
  nnd2s1 \IDinst/U6098  ( .DIN1(\IDinst/n6077 ), .DIN2(n671), 
        .Q(\IDinst/n6099 ) );
  nnd2s1 \IDinst/U6097  ( .DIN1(\IDinst/n6097 ), .DIN2(\IDinst/n6096 ), 
        .Q(\IDinst/n6098 ) );
  nnd2s1 \IDinst/U6096  ( .DIN1(\IDinst/n6095 ), .DIN2(n1197), 
        .Q(\IDinst/n6097 ) );
  nnd2s1 \IDinst/U6095  ( .DIN1(\IDinst/n6086 ), .DIN2(n1181), 
        .Q(\IDinst/n6096 ) );
  nnd2s1 \IDinst/U6094  ( .DIN1(\IDinst/n6094 ), .DIN2(\IDinst/n6093 ), 
        .Q(\IDinst/n6095 ) );
  nnd2s1 \IDinst/U6093  ( .DIN1(\IDinst/n6092 ), .DIN2(n1166), 
        .Q(\IDinst/n6094 ) );
  nnd2s1 \IDinst/U6092  ( .DIN1(\IDinst/n6089 ), .DIN2(n1143), 
        .Q(\IDinst/n6093 ) );
  nnd2s1 \IDinst/U6091  ( .DIN1(\IDinst/n6091 ), .DIN2(\IDinst/n6090 ), 
        .Q(\IDinst/n6092 ) );
  nnd2s1 \IDinst/U6090  ( .DIN1(\IDinst/RegFile[31][0] ), .DIN2(n1107), 
        .Q(\IDinst/n6091 ) );
  nnd2s1 \IDinst/U6089  ( .DIN1(\IDinst/RegFile[30][0] ), .DIN2(n1036), 
        .Q(\IDinst/n6090 ) );
  nnd2s1 \IDinst/U6088  ( .DIN1(\IDinst/n6088 ), .DIN2(\IDinst/n6087 ), 
        .Q(\IDinst/n6089 ) );
  nnd2s1 \IDinst/U6087  ( .DIN1(\IDinst/RegFile[29][0] ), .DIN2(n1108), 
        .Q(\IDinst/n6088 ) );
  nnd2s1 \IDinst/U6086  ( .DIN1(\IDinst/RegFile[28][0] ), .DIN2(n1036), 
        .Q(\IDinst/n6087 ) );
  nnd2s1 \IDinst/U6085  ( .DIN1(\IDinst/n6085 ), .DIN2(\IDinst/n6084 ), 
        .Q(\IDinst/n6086 ) );
  nnd2s1 \IDinst/U6084  ( .DIN1(\IDinst/n6083 ), .DIN2(n1166), 
        .Q(\IDinst/n6085 ) );
  nnd2s1 \IDinst/U6083  ( .DIN1(\IDinst/n6080 ), .DIN2(n1143), 
        .Q(\IDinst/n6084 ) );
  nnd2s1 \IDinst/U6082  ( .DIN1(\IDinst/n6082 ), .DIN2(\IDinst/n6081 ), 
        .Q(\IDinst/n6083 ) );
  nnd2s1 \IDinst/U6081  ( .DIN1(\IDinst/RegFile[27][0] ), .DIN2(n1108), 
        .Q(\IDinst/n6082 ) );
  nnd2s1 \IDinst/U6080  ( .DIN1(\IDinst/RegFile[26][0] ), .DIN2(n1036), 
        .Q(\IDinst/n6081 ) );
  nnd2s1 \IDinst/U6079  ( .DIN1(\IDinst/n6079 ), .DIN2(\IDinst/n6078 ), 
        .Q(\IDinst/n6080 ) );
  nnd2s1 \IDinst/U6078  ( .DIN1(\IDinst/RegFile[25][0] ), .DIN2(n1108), 
        .Q(\IDinst/n6079 ) );
  nnd2s1 \IDinst/U6077  ( .DIN1(\IDinst/RegFile[24][0] ), .DIN2(n1036), 
        .Q(\IDinst/n6078 ) );
  nnd2s1 \IDinst/U6076  ( .DIN1(\IDinst/n6076 ), .DIN2(\IDinst/n6075 ), 
        .Q(\IDinst/n6077 ) );
  nnd2s1 \IDinst/U6075  ( .DIN1(\IDinst/n6074 ), .DIN2(n1197), 
        .Q(\IDinst/n6076 ) );
  nnd2s1 \IDinst/U6074  ( .DIN1(\IDinst/n6065 ), .DIN2(n1181), 
        .Q(\IDinst/n6075 ) );
  nnd2s1 \IDinst/U6073  ( .DIN1(\IDinst/n6073 ), .DIN2(\IDinst/n6072 ), 
        .Q(\IDinst/n6074 ) );
  nnd2s1 \IDinst/U6072  ( .DIN1(\IDinst/n6071 ), .DIN2(n1166), 
        .Q(\IDinst/n6073 ) );
  nnd2s1 \IDinst/U6071  ( .DIN1(\IDinst/n6068 ), .DIN2(n1143), 
        .Q(\IDinst/n6072 ) );
  nnd2s1 \IDinst/U6070  ( .DIN1(\IDinst/n6070 ), .DIN2(\IDinst/n6069 ), 
        .Q(\IDinst/n6071 ) );
  nnd2s1 \IDinst/U6069  ( .DIN1(\IDinst/RegFile[23][0] ), .DIN2(n1108), 
        .Q(\IDinst/n6070 ) );
  nnd2s1 \IDinst/U6068  ( .DIN1(\IDinst/RegFile[22][0] ), .DIN2(n1036), 
        .Q(\IDinst/n6069 ) );
  nnd2s1 \IDinst/U6067  ( .DIN1(\IDinst/n6067 ), .DIN2(\IDinst/n6066 ), 
        .Q(\IDinst/n6068 ) );
  nnd2s1 \IDinst/U6066  ( .DIN1(\IDinst/RegFile[21][0] ), .DIN2(n1108), 
        .Q(\IDinst/n6067 ) );
  nnd2s1 \IDinst/U6065  ( .DIN1(\IDinst/RegFile[20][0] ), .DIN2(n1036), 
        .Q(\IDinst/n6066 ) );
  nnd2s1 \IDinst/U6064  ( .DIN1(\IDinst/n6064 ), .DIN2(\IDinst/n6063 ), 
        .Q(\IDinst/n6065 ) );
  nnd2s1 \IDinst/U6063  ( .DIN1(\IDinst/n6062 ), .DIN2(n1166), 
        .Q(\IDinst/n6064 ) );
  nnd2s1 \IDinst/U6062  ( .DIN1(\IDinst/n6059 ), .DIN2(n1143), 
        .Q(\IDinst/n6063 ) );
  nnd2s1 \IDinst/U6061  ( .DIN1(\IDinst/n6061 ), .DIN2(\IDinst/n6060 ), 
        .Q(\IDinst/n6062 ) );
  nnd2s1 \IDinst/U6060  ( .DIN1(\IDinst/RegFile[19][0] ), .DIN2(n1108), 
        .Q(\IDinst/n6061 ) );
  nnd2s1 \IDinst/U6059  ( .DIN1(\IDinst/RegFile[18][0] ), .DIN2(n1036), 
        .Q(\IDinst/n6060 ) );
  nnd2s1 \IDinst/U6058  ( .DIN1(\IDinst/n6058 ), .DIN2(\IDinst/n6057 ), 
        .Q(\IDinst/n6059 ) );
  nnd2s1 \IDinst/U6057  ( .DIN1(\IDinst/RegFile[17][0] ), .DIN2(n1108), 
        .Q(\IDinst/n6058 ) );
  nnd2s1 \IDinst/U6056  ( .DIN1(\IDinst/RegFile[16][0] ), .DIN2(n1036), 
        .Q(\IDinst/n6057 ) );
  nnd2s1 \IDinst/U6055  ( .DIN1(\IDinst/n6055 ), .DIN2(\IDinst/n6054 ), 
        .Q(\IDinst/n6056 ) );
  nnd2s1 \IDinst/U6054  ( .DIN1(n644), .DIN2(\IDinst/n6053 ), 
        .Q(\IDinst/n6055 ) );
  nnd2s1 \IDinst/U6053  ( .DIN1(\IDinst/n6032 ), .DIN2(n672), 
        .Q(\IDinst/n6054 ) );
  nnd2s1 \IDinst/U6052  ( .DIN1(\IDinst/n6052 ), .DIN2(\IDinst/n6051 ), 
        .Q(\IDinst/n6053 ) );
  nnd2s1 \IDinst/U6051  ( .DIN1(\IDinst/n6050 ), .DIN2(n1197), 
        .Q(\IDinst/n6052 ) );
  nnd2s1 \IDinst/U6050  ( .DIN1(\IDinst/n6041 ), .DIN2(n1181), 
        .Q(\IDinst/n6051 ) );
  nnd2s1 \IDinst/U6049  ( .DIN1(\IDinst/n6049 ), .DIN2(\IDinst/n6048 ), 
        .Q(\IDinst/n6050 ) );
  nnd2s1 \IDinst/U6048  ( .DIN1(\IDinst/n6047 ), .DIN2(n1166), 
        .Q(\IDinst/n6049 ) );
  nnd2s1 \IDinst/U6047  ( .DIN1(\IDinst/n6044 ), .DIN2(n1143), 
        .Q(\IDinst/n6048 ) );
  nnd2s1 \IDinst/U6046  ( .DIN1(\IDinst/n6046 ), .DIN2(\IDinst/n6045 ), 
        .Q(\IDinst/n6047 ) );
  nnd2s1 \IDinst/U6045  ( .DIN1(\IDinst/RegFile[15][0] ), .DIN2(n1108), 
        .Q(\IDinst/n6046 ) );
  nnd2s1 \IDinst/U6044  ( .DIN1(\IDinst/RegFile[14][0] ), .DIN2(n1035), 
        .Q(\IDinst/n6045 ) );
  nnd2s1 \IDinst/U6043  ( .DIN1(\IDinst/n6043 ), .DIN2(\IDinst/n6042 ), 
        .Q(\IDinst/n6044 ) );
  nnd2s1 \IDinst/U6042  ( .DIN1(\IDinst/RegFile[13][0] ), .DIN2(n1108), 
        .Q(\IDinst/n6043 ) );
  nnd2s1 \IDinst/U6041  ( .DIN1(\IDinst/RegFile[12][0] ), .DIN2(n1035), 
        .Q(\IDinst/n6042 ) );
  nnd2s1 \IDinst/U6040  ( .DIN1(\IDinst/n6040 ), .DIN2(\IDinst/n6039 ), 
        .Q(\IDinst/n6041 ) );
  nnd2s1 \IDinst/U6039  ( .DIN1(\IDinst/n6038 ), .DIN2(n1166), 
        .Q(\IDinst/n6040 ) );
  nnd2s1 \IDinst/U6038  ( .DIN1(\IDinst/n6035 ), .DIN2(n1143), 
        .Q(\IDinst/n6039 ) );
  nnd2s1 \IDinst/U6037  ( .DIN1(\IDinst/n6037 ), .DIN2(\IDinst/n6036 ), 
        .Q(\IDinst/n6038 ) );
  nnd2s1 \IDinst/U6036  ( .DIN1(\IDinst/RegFile[11][0] ), .DIN2(n1109), 
        .Q(\IDinst/n6037 ) );
  nnd2s1 \IDinst/U6035  ( .DIN1(\IDinst/RegFile[10][0] ), .DIN2(n1035), 
        .Q(\IDinst/n6036 ) );
  nnd2s1 \IDinst/U6034  ( .DIN1(\IDinst/n6034 ), .DIN2(\IDinst/n6033 ), 
        .Q(\IDinst/n6035 ) );
  nnd2s1 \IDinst/U6033  ( .DIN1(\IDinst/RegFile[9][0] ), .DIN2(n1109), 
        .Q(\IDinst/n6034 ) );
  nnd2s1 \IDinst/U6032  ( .DIN1(\IDinst/RegFile[8][0] ), .DIN2(n1035), 
        .Q(\IDinst/n6033 ) );
  nnd2s1 \IDinst/U6031  ( .DIN1(\IDinst/n6031 ), .DIN2(\IDinst/n6030 ), 
        .Q(\IDinst/n6032 ) );
  nnd2s1 \IDinst/U6030  ( .DIN1(n1196), .DIN2(\IDinst/n6029 ), 
        .Q(\IDinst/n6031 ) );
  nnd2s1 \IDinst/U6029  ( .DIN1(\IDinst/n6020 ), .DIN2(n1185), 
        .Q(\IDinst/n6030 ) );
  nnd2s1 \IDinst/U6028  ( .DIN1(\IDinst/n6028 ), .DIN2(\IDinst/n6027 ), 
        .Q(\IDinst/n6029 ) );
  nnd2s1 \IDinst/U6027  ( .DIN1(\IDinst/n6026 ), .DIN2(n1166), 
        .Q(\IDinst/n6028 ) );
  nnd2s1 \IDinst/U6026  ( .DIN1(\IDinst/n6023 ), .DIN2(n1133), 
        .Q(\IDinst/n6027 ) );
  nnd2s1 \IDinst/U6025  ( .DIN1(\IDinst/n6025 ), .DIN2(\IDinst/n6024 ), 
        .Q(\IDinst/n6026 ) );
  nnd2s1 \IDinst/U6024  ( .DIN1(\IDinst/RegFile[7][0] ), .DIN2(n1109), 
        .Q(\IDinst/n6025 ) );
  nnd2s1 \IDinst/U6023  ( .DIN1(\IDinst/RegFile[6][0] ), .DIN2(n1035), 
        .Q(\IDinst/n6024 ) );
  nnd2s1 \IDinst/U6022  ( .DIN1(\IDinst/n6022 ), .DIN2(\IDinst/n6021 ), 
        .Q(\IDinst/n6023 ) );
  nnd2s1 \IDinst/U6021  ( .DIN1(\IDinst/RegFile[5][0] ), .DIN2(n1109), 
        .Q(\IDinst/n6022 ) );
  nnd2s1 \IDinst/U6020  ( .DIN1(\IDinst/RegFile[4][0] ), .DIN2(n1040), 
        .Q(\IDinst/n6021 ) );
  nnd2s1 \IDinst/U6019  ( .DIN1(\IDinst/n6019 ), .DIN2(\IDinst/n6018 ), 
        .Q(\IDinst/n6020 ) );
  nnd2s1 \IDinst/U6018  ( .DIN1(n1153), .DIN2(\IDinst/n6017 ), 
        .Q(\IDinst/n6019 ) );
  nnd2s1 \IDinst/U6017  ( .DIN1(\IDinst/n6014 ), .DIN2(n1143), 
        .Q(\IDinst/n6018 ) );
  nnd2s1 \IDinst/U6016  ( .DIN1(\IDinst/n6016 ), .DIN2(\IDinst/n6015 ), 
        .Q(\IDinst/n6017 ) );
  nnd2s1 \IDinst/U6015  ( .DIN1(\IDinst/RegFile[3][0] ), .DIN2(n1109), 
        .Q(\IDinst/n6016 ) );
  nnd2s1 \IDinst/U6014  ( .DIN1(\IDinst/RegFile[2][0] ), .DIN2(n1025), 
        .Q(\IDinst/n6015 ) );
  nnd2s1 \IDinst/U6013  ( .DIN1(\IDinst/n6013 ), .DIN2(\IDinst/n6012 ), 
        .Q(\IDinst/n6014 ) );
  nnd2s1 \IDinst/U6012  ( .DIN1(\IDinst/RegFile[1][0] ), .DIN2(n1096), 
        .Q(\IDinst/n6013 ) );
  nnd2s1 \IDinst/U6011  ( .DIN1(\IDinst/RegFile[0][0] ), .DIN2(n1045), 
        .Q(\IDinst/n6012 ) );
  nnd2s1 \IDinst/U6010  ( .DIN1(\IDinst/n6010 ), .DIN2(\IDinst/n6011 ), 
        .Q(\IDinst/N54 ) );
  nnd2s1 \IDinst/U6009  ( .DIN1(\IDinst/n6008 ), .DIN2(\IDinst/n6009 ), 
        .Q(\IDinst/N55 ) );
  nnd2s1 \IDinst/U6008  ( .DIN1(\IDinst/n6006 ), .DIN2(\IDinst/n6007 ), 
        .Q(\IDinst/N56 ) );
  nnd2s1 \IDinst/U6007  ( .DIN1(\IDinst/n6004 ), .DIN2(\IDinst/n6005 ), 
        .Q(\IDinst/N57 ) );
  nnd2s1 \IDinst/U6006  ( .DIN1(\IDinst/n6002 ), .DIN2(\IDinst/n6003 ), 
        .Q(\IDinst/N58 ) );
  nnd2s1 \IDinst/U6005  ( .DIN1(\IDinst/n6000 ), .DIN2(\IDinst/n6001 ), 
        .Q(\IDinst/N59 ) );
  nnd2s1 \IDinst/U6004  ( .DIN1(\IDinst/n5998 ), .DIN2(\IDinst/n5999 ), 
        .Q(\IDinst/N60 ) );
  nnd2s1 \IDinst/U6003  ( .DIN1(\IDinst/n5996 ), .DIN2(\IDinst/n5997 ), 
        .Q(\IDinst/N61 ) );
  nnd2s1 \IDinst/U6002  ( .DIN1(\IDinst/n5994 ), .DIN2(\IDinst/n5995 ), 
        .Q(\IDinst/N62 ) );
  nnd2s1 \IDinst/U6001  ( .DIN1(\IDinst/n5992 ), .DIN2(\IDinst/n5993 ), 
        .Q(\IDinst/N63 ) );
  nnd2s1 \IDinst/U6000  ( .DIN1(\IDinst/n5990 ), .DIN2(\IDinst/n5991 ), 
        .Q(\IDinst/N64 ) );
  nnd2s1 \IDinst/U5999  ( .DIN1(\IDinst/n5988 ), .DIN2(\IDinst/n5989 ), 
        .Q(\IDinst/N65 ) );
  nnd2s1 \IDinst/U5998  ( .DIN1(\IDinst/n5986 ), .DIN2(\IDinst/n5987 ), 
        .Q(\IDinst/N66 ) );
  nnd2s1 \IDinst/U5997  ( .DIN1(\IDinst/n5984 ), .DIN2(\IDinst/n5985 ), 
        .Q(\IDinst/N67 ) );
  nnd2s1 \IDinst/U5996  ( .DIN1(\IDinst/n5982 ), .DIN2(\IDinst/n5983 ), 
        .Q(\IDinst/N68 ) );
  nnd2s1 \IDinst/U5995  ( .DIN1(\IDinst/n5980 ), .DIN2(\IDinst/n5981 ), 
        .Q(\IDinst/N69 ) );
  nnd2s1 \IDinst/U5994  ( .DIN1(\IDinst/n5978 ), .DIN2(\IDinst/n5979 ), 
        .Q(\IDinst/N70 ) );
  nnd2s1 \IDinst/U5993  ( .DIN1(\IDinst/n5976 ), .DIN2(\IDinst/n5977 ), 
        .Q(\IDinst/N71 ) );
  nnd2s1 \IDinst/U5992  ( .DIN1(\IDinst/n5974 ), .DIN2(\IDinst/n5975 ), 
        .Q(\IDinst/N72 ) );
  nnd2s1 \IDinst/U5991  ( .DIN1(\IDinst/n5972 ), .DIN2(\IDinst/n5973 ), 
        .Q(\IDinst/N73 ) );
  nnd2s1 \IDinst/U5990  ( .DIN1(\IDinst/n5970 ), .DIN2(\IDinst/n5971 ), 
        .Q(\IDinst/N74 ) );
  nnd2s1 \IDinst/U5989  ( .DIN1(\IDinst/n5968 ), .DIN2(\IDinst/n5969 ), 
        .Q(\IDinst/N75 ) );
  nnd2s1 \IDinst/U5988  ( .DIN1(\IDinst/n5966 ), .DIN2(\IDinst/n5967 ), 
        .Q(\IDinst/N76 ) );
  nnd2s1 \IDinst/U5987  ( .DIN1(\IDinst/n5964 ), .DIN2(\IDinst/n5965 ), 
        .Q(\IDinst/N77 ) );
  nnd2s1 \IDinst/U5986  ( .DIN1(\IDinst/n5962 ), .DIN2(\IDinst/n5963 ), 
        .Q(\IDinst/N78 ) );
  nnd2s1 \IDinst/U5985  ( .DIN1(\IDinst/n5960 ), .DIN2(\IDinst/n5961 ), 
        .Q(\IDinst/N79 ) );
  nnd2s1 \IDinst/U5984  ( .DIN1(\IDinst/n5958 ), .DIN2(\IDinst/n5959 ), 
        .Q(\IDinst/N80 ) );
  nnd2s1 \IDinst/U5983  ( .DIN1(\IDinst/n5956 ), .DIN2(\IDinst/n5957 ), 
        .Q(\IDinst/N81 ) );
  nnd2s1 \IDinst/U5982  ( .DIN1(\IDinst/n5954 ), .DIN2(\IDinst/n5955 ), 
        .Q(\IDinst/N82 ) );
  nnd2s1 \IDinst/U5981  ( .DIN1(\IDinst/n5952 ), .DIN2(\IDinst/n5953 ), 
        .Q(\IDinst/N83 ) );
  nnd2s1 \IDinst/U5980  ( .DIN1(\IDinst/n5950 ), .DIN2(\IDinst/n5951 ), 
        .Q(\IDinst/N84 ) );
  nnd2s1 \IDinst/U5979  ( .DIN1(\IDinst/n5948 ), .DIN2(\IDinst/n5949 ), 
        .Q(\IDinst/N85 ) );
  dffascs1 \IDinst/reg_out_A_reg[0]  ( .DIN(\IDinst/N992 ), .CLK(clk), 
        .CLRB(n926), .SETB(1'b1), .Q(n33), .QN(n331) );
  dffascs1 \IDinst/Cause_Reg_reg[0]  ( .DIN(\IDinst/n4729 ), .CLK(clk), 
        .CLRB(n950), .SETB(1'b1), .Q(n271) );
  dffascs1 \IDinst/Imm_reg[0]  ( .DIN(\IDinst/n4730 ), .CLK(clk), .CLRB(n950), 
        .SETB(1'b1), .QN(n9489) );
  dffascs1 \IDinst/reg_out_A_reg[1]  ( .DIN(\IDinst/N993 ), .CLK(clk), 
        .CLRB(n830), .SETB(1'b1), .Q(n35), .QN(n330) );
  dffascs1 \IDinst/Cause_Reg_reg[1]  ( .DIN(\IDinst/n4731 ), .CLK(clk), 
        .CLRB(n950), .SETB(1'b1), .Q(n270) );
  dffascs1 \IDinst/Imm_reg[1]  ( .DIN(\IDinst/n4732 ), .CLK(clk), .CLRB(n950), 
        .SETB(1'b1), .Q(n711), .QN(n9488) );
  dffascs1 \IDinst/reg_out_A_reg[2]  ( .DIN(\IDinst/N994 ), .CLK(clk), 
        .CLRB(n830), .SETB(1'b1), .QN(n80) );
  dffascs1 \IDinst/Cause_Reg_reg[2]  ( .DIN(\IDinst/n4733 ), .CLK(clk), 
        .CLRB(n950), .SETB(1'b1), .Q(n269) );
  dffascs1 \IDinst/Imm_reg[2]  ( .DIN(\IDinst/n4734 ), .CLK(clk), .CLRB(n950), 
        .SETB(1'b1), .Q(n207), .QN(n29) );
  dffascs1 \IDinst/reg_out_A_reg[3]  ( .DIN(\IDinst/N995 ), .CLK(clk), 
        .CLRB(n833), .SETB(1'b1), .QN(n77) );
  dffascs1 \IDinst/Cause_Reg_reg[3]  ( .DIN(\IDinst/n4735 ), .CLK(clk), 
        .CLRB(n949), .SETB(1'b1), .Q(n268) );
  dffascs1 \IDinst/Imm_reg[3]  ( .DIN(\IDinst/n4736 ), .CLK(clk), .CLRB(n949), 
        .SETB(1'b1), .Q(n735), .QN(n9487) );
  dffascs1 \IDinst/reg_out_A_reg[4]  ( .DIN(\IDinst/N996 ), .CLK(clk), 
        .CLRB(n832), .SETB(1'b1), .Q(n10), .QN(n334) );
  dffascs1 \IDinst/Cause_Reg_reg[4]  ( .DIN(\IDinst/n4737 ), .CLK(clk), 
        .CLRB(n949), .SETB(1'b1), .Q(n267) );
  dffascs1 \IDinst/Imm_reg[4]  ( .DIN(\IDinst/n4738 ), .CLK(clk), .CLRB(n949), 
        .SETB(1'b1), .Q(n206), .QN(n56) );
  dffascs1 \IDinst/reg_out_A_reg[5]  ( .DIN(\IDinst/N997 ), .CLK(clk), 
        .CLRB(n832), .SETB(1'b1), .QN(n81) );
  dffascs1 \IDinst/Cause_Reg_reg[5]  ( .DIN(\IDinst/n4739 ), .CLK(clk), 
        .CLRB(n949), .SETB(1'b1), .Q(n266) );
  dffascs1 \IDinst/Imm_reg[5]  ( .DIN(\IDinst/n4740 ), .CLK(clk), .CLRB(n949), 
        .SETB(1'b1), .QN(n9486) );
  dffascs1 \IDinst/reg_out_A_reg[6]  ( .DIN(\IDinst/N998 ), .CLK(clk), 
        .CLRB(n845), .SETB(1'b1), .Q(n34), .QN(n333) );
  dffascs1 \IDinst/Cause_Reg_reg[6]  ( .DIN(\IDinst/n4741 ), .CLK(clk), 
        .CLRB(n949), .SETB(1'b1), .Q(n265) );
  dffascs1 \IDinst/Imm_reg[6]  ( .DIN(\IDinst/n4742 ), .CLK(clk), .CLRB(n949), 
        .SETB(1'b1), .Q(n105), .QN(n9485) );
  dffascs1 \IDinst/reg_out_A_reg[7]  ( .DIN(\IDinst/N999 ), .CLK(clk), 
        .CLRB(n849), .SETB(1'b1), .QN(n63) );
  dffascs1 \IDinst/Cause_Reg_reg[7]  ( .DIN(\IDinst/n4743 ), .CLK(clk), 
        .CLRB(n949), .SETB(1'b1), .Q(n264) );
  dffascs1 \IDinst/Imm_reg[7]  ( .DIN(\IDinst/n4744 ), .CLK(clk), .CLRB(n949), 
        .SETB(1'b1), .Q(n76), .QN(n9484) );
  dffascs1 \IDinst/reg_out_A_reg[8]  ( .DIN(\IDinst/N1000 ), .CLK(clk), 
        .CLRB(n845), .SETB(1'b1), .Q(n36), .QN(n332) );
  dffascs1 \IDinst/Cause_Reg_reg[8]  ( .DIN(\IDinst/n4745 ), .CLK(clk), 
        .CLRB(n948), .SETB(1'b1), .Q(n305) );
  dffascs1 \IDinst/Imm_reg[8]  ( .DIN(\IDinst/n4746 ), .CLK(clk), .CLRB(n948), 
        .SETB(1'b1), .Q(n107), .QN(n9483) );
  dffascs1 \IDinst/reg_out_A_reg[9]  ( .DIN(\IDinst/N1001 ), .CLK(clk), 
        .CLRB(n844), .SETB(1'b1), .QN(n66) );
  dffascs1 \IDinst/Cause_Reg_reg[9]  ( .DIN(\IDinst/n4747 ), .CLK(clk), 
        .CLRB(n948), .SETB(1'b1), .Q(n304) );
  dffascs1 \IDinst/Imm_reg[9]  ( .DIN(\IDinst/n4748 ), .CLK(clk), .CLRB(n948), 
        .SETB(1'b1), .Q(n75), .QN(n9482) );
  dffascs1 \IDinst/reg_out_A_reg[10]  ( .DIN(\IDinst/N1002 ), .CLK(clk), 
        .CLRB(n856), .SETB(1'b1), .QN(n65) );
  dffascs1 \IDinst/Cause_Reg_reg[10]  ( .DIN(\IDinst/n4749 ), .CLK(clk), 
        .CLRB(n948), .SETB(1'b1), .Q(n303) );
  dffascs1 \IDinst/Imm_reg[10]  ( .DIN(\IDinst/n4750 ), .CLK(clk), .CLRB(n948), 
        .SETB(1'b1), .Q(n104), .QN(n9481) );
  dffascs1 \IDinst/reg_out_A_reg[11]  ( .DIN(\IDinst/N1003 ), .CLK(clk), 
        .CLRB(n856), .SETB(1'b1), .QN(n84) );
  dffascs1 \IDinst/Cause_Reg_reg[11]  ( .DIN(\IDinst/n4751 ), .CLK(clk), 
        .CLRB(n948), .SETB(1'b1), .Q(n302) );
  dffascs1 \IDinst/Imm_reg[11]  ( .DIN(\IDinst/n4752 ), .CLK(clk), .CLRB(n948), 
        .SETB(1'b1), .Q(n8), .QN(n9480) );
  dffascs1 \IDinst/reg_out_A_reg[12]  ( .DIN(\IDinst/N1004 ), .CLK(clk), 
        .CLRB(n831), .SETB(1'b1), .QN(n64) );
  dffascs1 \IDinst/Cause_Reg_reg[12]  ( .DIN(\IDinst/n4753 ), .CLK(clk), 
        .CLRB(n948), .SETB(1'b1), .Q(n301) );
  dffascs1 \IDinst/Imm_reg[12]  ( .DIN(\IDinst/n4754 ), .CLK(clk), .CLRB(n948), 
        .SETB(1'b1), .Q(n106), .QN(n9479) );
  dffascs1 \IDinst/reg_out_A_reg[13]  ( .DIN(\IDinst/N1005 ), .CLK(clk), 
        .CLRB(n875), .SETB(1'b1), .QN(n86) );
  dffascs1 \IDinst/Cause_Reg_reg[13]  ( .DIN(\IDinst/n4755 ), .CLK(clk), 
        .CLRB(n947), .SETB(1'b1), .Q(n300) );
  dffascs1 \IDinst/Imm_reg[13]  ( .DIN(\IDinst/n4756 ), .CLK(clk), .CLRB(n947), 
        .SETB(1'b1), .Q(n9), .QN(n9478) );
  dffascs1 \IDinst/reg_out_A_reg[14]  ( .DIN(\IDinst/N1006 ), .CLK(clk), 
        .CLRB(n864), .SETB(1'b1), .QN(n31) );
  dffascs1 \IDinst/Cause_Reg_reg[14]  ( .DIN(\IDinst/n4757 ), .CLK(clk), 
        .CLRB(n947), .SETB(1'b1), .Q(n299) );
  dffascs1 \IDinst/Imm_reg[14]  ( .DIN(\IDinst/n4758 ), .CLK(clk), .CLRB(n947), 
        .SETB(1'b1), .Q(n108), .QN(n9477) );
  dffascs1 \IDinst/reg_out_A_reg[15]  ( .DIN(\IDinst/N1007 ), .CLK(clk), 
        .CLRB(n864), .SETB(1'b1), .QN(n85) );
  dffascs1 \IDinst/Cause_Reg_reg[15]  ( .DIN(\IDinst/n4759 ), .CLK(clk), 
        .CLRB(n947), .SETB(1'b1), .Q(n298) );
  dffascs1 \IDinst/Imm_reg[15]  ( .DIN(\IDinst/n4760 ), .CLK(clk), .CLRB(n947), 
        .SETB(1'b1), .Q(n7), .QN(n9476) );
  dffascs1 \IDinst/reg_out_A_reg[16]  ( .DIN(\IDinst/N1008 ), .CLK(clk), 
        .CLRB(n914), .SETB(1'b1), .QN(n71) );
  dffascs1 \IDinst/Cause_Reg_reg[16]  ( .DIN(\IDinst/n4761 ), .CLK(clk), 
        .CLRB(n947), .SETB(1'b1), .Q(n297) );
  dffascs1 \IDinst/Imm_reg[16]  ( .DIN(\IDinst/n4762 ), .CLK(clk), .CLRB(n947), 
        .SETB(1'b1), .Q(n109), .QN(n9475) );
  dffascs1 \IDinst/reg_out_A_reg[17]  ( .DIN(\IDinst/N1009 ), .CLK(clk), 
        .CLRB(n913), .SETB(1'b1), .QN(n82) );
  dffascs1 \IDinst/Cause_Reg_reg[17]  ( .DIN(\IDinst/n4763 ), .CLK(clk), 
        .CLRB(n947), .SETB(1'b1), .Q(n296) );
  dffascs1 \IDinst/Imm_reg[17]  ( .DIN(\IDinst/n4764 ), .CLK(clk), .CLRB(n947), 
        .SETB(1'b1), .Q(n13), .QN(n9474) );
  dffascs1 \IDinst/reg_out_A_reg[18]  ( .DIN(\IDinst/N1010 ), .CLK(clk), 
        .CLRB(n872), .SETB(1'b1), .QN(n70) );
  dffascs1 \IDinst/Cause_Reg_reg[18]  ( .DIN(\IDinst/n4765 ), .CLK(clk), 
        .CLRB(n946), .SETB(1'b1), .Q(n295) );
  dffascs1 \IDinst/Imm_reg[18]  ( .DIN(\IDinst/n4766 ), .CLK(clk), .CLRB(n946), 
        .SETB(1'b1), .Q(n122), .QN(n9473) );
  dffascs1 \IDinst/reg_out_A_reg[19]  ( .DIN(\IDinst/N1011 ), .CLK(clk), 
        .CLRB(n871), .SETB(1'b1), .QN(n37) );
  dffascs1 \IDinst/Cause_Reg_reg[19]  ( .DIN(\IDinst/n4767 ), .CLK(clk), 
        .CLRB(n946), .SETB(1'b1), .Q(n294) );
  dffascs1 \IDinst/Imm_reg[19]  ( .DIN(\IDinst/n4768 ), .CLK(clk), .CLRB(n946), 
        .SETB(1'b1), .Q(n94), .QN(n9472) );
  dffascs1 \IDinst/reg_out_A_reg[20]  ( .DIN(\IDinst/N1012 ), .CLK(clk), 
        .CLRB(n884), .SETB(1'b1), .QN(n69) );
  dffascs1 \IDinst/Cause_Reg_reg[20]  ( .DIN(\IDinst/n4769 ), .CLK(clk), 
        .CLRB(n946), .SETB(1'b1), .Q(n293) );
  dffascs1 \IDinst/Imm_reg[20]  ( .DIN(\IDinst/n4770 ), .CLK(clk), .CLRB(n946), 
        .SETB(1'b1), .Q(n123), .QN(n9471) );
  dffascs1 \IDinst/reg_out_A_reg[21]  ( .DIN(\IDinst/N1013 ), .CLK(clk), 
        .CLRB(n884), .SETB(1'b1), .QN(n78) );
  dffascs1 \IDinst/Cause_Reg_reg[21]  ( .DIN(\IDinst/n4771 ), .CLK(clk), 
        .CLRB(n946), .SETB(1'b1), .Q(n292) );
  dffascs1 \IDinst/Imm_reg[21]  ( .DIN(\IDinst/n4772 ), .CLK(clk), .CLRB(n946), 
        .SETB(1'b1), .Q(n16), .QN(n9470) );
  dffascs1 \IDinst/reg_out_A_reg[22]  ( .DIN(\IDinst/N1014 ), .CLK(clk), 
        .CLRB(n880), .SETB(1'b1), .QN(n67) );
  dffascs1 \IDinst/Cause_Reg_reg[22]  ( .DIN(\IDinst/n4773 ), .CLK(clk), 
        .CLRB(n946), .SETB(1'b1), .Q(n291) );
  dffascs1 \IDinst/Imm_reg[22]  ( .DIN(\IDinst/n4774 ), .CLK(clk), .CLRB(n946), 
        .SETB(1'b1), .Q(n121), .QN(n9469) );
  dffascs1 \IDinst/reg_out_A_reg[23]  ( .DIN(\IDinst/N1015 ), .CLK(clk), 
        .CLRB(n888), .SETB(1'b1), .QN(n68) );
  dffascs1 \IDinst/Cause_Reg_reg[23]  ( .DIN(\IDinst/n4775 ), .CLK(clk), 
        .CLRB(n945), .SETB(1'b1), .Q(n290) );
  dffascs1 \IDinst/Imm_reg[23]  ( .DIN(\IDinst/n4776 ), .CLK(clk), .CLRB(n945), 
        .SETB(1'b1), .Q(n93), .QN(n9468) );
  dffascs1 \IDinst/reg_out_A_reg[24]  ( .DIN(\IDinst/N1016 ), .CLK(clk), 
        .CLRB(n880), .SETB(1'b1), .QN(n30) );
  dffascs1 \IDinst/Cause_Reg_reg[24]  ( .DIN(\IDinst/n4777 ), .CLK(clk), 
        .CLRB(n945), .SETB(1'b1), .Q(n289) );
  dffascs1 \IDinst/Imm_reg[24]  ( .DIN(\IDinst/n4778 ), .CLK(clk), .CLRB(n945), 
        .SETB(1'b1), .Q(n120), .QN(n9467) );
  dffascs1 \IDinst/reg_out_A_reg[25]  ( .DIN(\IDinst/N1017 ), .CLK(clk), 
        .CLRB(n899), .SETB(1'b1), .QN(n83) );
  dffascs1 \IDinst/Cause_Reg_reg[25]  ( .DIN(\IDinst/n4779 ), .CLK(clk), 
        .CLRB(n945), .SETB(1'b1), .Q(n288) );
  dffascs1 \IDinst/Imm_reg[25]  ( .DIN(\IDinst/n4780 ), .CLK(clk), .CLRB(n945), 
        .SETB(1'b1), .Q(n15), .QN(n9466) );
  dffascs1 \IDinst/reg_out_A_reg[26]  ( .DIN(\IDinst/N1018 ), .CLK(clk), 
        .CLRB(n879), .SETB(1'b1), .Q(n6), .QN(n336) );
  dffascs1 \IDinst/Cause_Reg_reg[26]  ( .DIN(\IDinst/n4781 ), .CLK(clk), 
        .CLRB(n945), .SETB(1'b1), .Q(n287) );
  dffascs1 \IDinst/Imm_reg[26]  ( .DIN(\IDinst/n4782 ), .CLK(clk), .CLRB(n945), 
        .SETB(1'b1), .Q(n103), .QN(n9465) );
  dffascs1 \IDinst/reg_out_A_reg[27]  ( .DIN(\IDinst/N1019 ), .CLK(clk), 
        .CLRB(n906), .SETB(1'b1), .QN(n38) );
  dffascs1 \IDinst/Cause_Reg_reg[27]  ( .DIN(\IDinst/n4783 ), .CLK(clk), 
        .CLRB(n945), .SETB(1'b1), .Q(n286) );
  dffascs1 \IDinst/Imm_reg[27]  ( .DIN(\IDinst/n4784 ), .CLK(clk), .CLRB(n945), 
        .SETB(1'b1), .Q(n95), .QN(n9464) );
  dffascs1 \IDinst/reg_out_A_reg[28]  ( .DIN(\IDinst/N1020 ), .CLK(clk), 
        .CLRB(n918), .SETB(1'b1), .Q(n12), .QN(n335) );
  dffascs1 \IDinst/Cause_Reg_reg[28]  ( .DIN(\IDinst/n4785 ), .CLK(clk), 
        .CLRB(n944), .SETB(1'b1), .Q(n285) );
  dffascs1 \IDinst/Imm_reg[28]  ( .DIN(\IDinst/n4786 ), .CLK(clk), .CLRB(n944), 
        .SETB(1'b1), .Q(n102), .QN(n9463) );
  dffascs1 \IDinst/reg_out_A_reg[29]  ( .DIN(\IDinst/N1021 ), .CLK(clk), 
        .CLRB(n831), .SETB(1'b1), .QN(n79) );
  dffascs1 \IDinst/Cause_Reg_reg[29]  ( .DIN(\IDinst/n4787 ), .CLK(clk), 
        .CLRB(n944), .SETB(1'b1), .Q(n284) );
  dffascs1 \IDinst/Imm_reg[29]  ( .DIN(\IDinst/n4788 ), .CLK(clk), .CLRB(n944), 
        .SETB(1'b1), .Q(n14), .QN(n9462) );
  dffascs1 \IDinst/reg_out_A_reg[30]  ( .DIN(\IDinst/N1022 ), .CLK(clk), 
        .CLRB(n830), .SETB(1'b1), .Q(reg_out_A[30]), .QN(n717) );
  dffascs1 \IDinst/Cause_Reg_reg[30]  ( .DIN(\IDinst/n4789 ), .CLK(clk), 
        .CLRB(n944), .SETB(1'b1), .Q(n283) );
  dffascs1 \IDinst/Imm_reg[30]  ( .DIN(\IDinst/n4790 ), .CLK(clk), .CLRB(n944), 
        .SETB(1'b1), .Q(n96), .QN(n9461) );
  dffascs1 \IDinst/reg_out_A_reg[31]  ( .DIN(\IDinst/N1023 ), .CLK(clk), 
        .CLRB(n918), .SETB(1'b1), .Q(reg_out_A[31]), .QN(n62) );
  dffascs1 \IDinst/Cause_Reg_reg[31]  ( .DIN(\IDinst/n4791 ), .CLK(clk), 
        .CLRB(n944), .SETB(1'b1), .Q(n282) );
  dffascs1 \IDinst/Imm_reg[31]  ( .DIN(\IDinst/n4792 ), .CLK(clk), .CLRB(n944), 
        .SETB(1'b1), .Q(n124), .QN(n9460) );
  dffascs1 \IDinst/reg_out_B_reg[31]  ( .DIN(\IDinst/N1055 ), .CLK(clk), 
        .CLRB(n963), .SETB(1'b1), .Q(reg_out_B[31]), .QN(n133) );
  dffascs1 \IDinst/reg_out_B_reg[30]  ( .DIN(\IDinst/N1054 ), .CLK(clk), 
        .CLRB(n962), .SETB(1'b1), .Q(reg_out_B[30]), .QN(n18) );
  dffascs1 \IDinst/reg_out_B_reg[29]  ( .DIN(\IDinst/N1053 ), .CLK(clk), 
        .CLRB(n809), .SETB(1'b1), .Q(reg_out_B[29]), .QN(n43) );
  dffascs1 \IDinst/reg_out_B_reg[28]  ( .DIN(\IDinst/N1052 ), .CLK(clk), 
        .CLRB(n809), .SETB(1'b1), .Q(reg_out_B[28]), .QN(n44) );
  dffascs1 \IDinst/reg_out_B_reg[27]  ( .DIN(\IDinst/N1051 ), .CLK(clk), 
        .CLRB(n810), .SETB(1'b1), .Q(reg_out_B[27]), .QN(n134) );
  dffascs1 \IDinst/reg_out_B_reg[26]  ( .DIN(\IDinst/N1050 ), .CLK(clk), 
        .CLRB(n910), .SETB(1'b1), .Q(reg_out_B[26]), .QN(n20) );
  dffascs1 \IDinst/reg_out_B_reg[25]  ( .DIN(\IDinst/N1049 ), .CLK(clk), 
        .CLRB(n810), .SETB(1'b1), .Q(reg_out_B[25]), .QN(n25) );
  dffascs1 \IDinst/reg_out_B_reg[24]  ( .DIN(\IDinst/N1048 ), .CLK(clk), 
        .CLRB(n902), .SETB(1'b1), .Q(reg_out_B[24]), .QN(n145) );
  dffascs1 \IDinst/reg_out_B_reg[23]  ( .DIN(\IDinst/N1047 ), .CLK(clk), 
        .CLRB(n811), .SETB(1'b1), .Q(reg_out_B[23]), .QN(n53) );
  dffascs1 \IDinst/reg_out_B_reg[22]  ( .DIN(\IDinst/N1046 ), .CLK(clk), 
        .CLRB(n812), .SETB(1'b1), .Q(reg_out_B[22]), .QN(n3) );
  dffascs1 \IDinst/reg_out_B_reg[21]  ( .DIN(\IDinst/N1045 ), .CLK(clk), 
        .CLRB(n824), .SETB(1'b1), .Q(reg_out_B[21]), .QN(n23) );
  dffascs1 \IDinst/reg_out_B_reg[20]  ( .DIN(\IDinst/N1044 ), .CLK(clk), 
        .CLRB(n811), .SETB(1'b1), .Q(reg_out_B[20]), .QN(n52) );
  dffascs1 \IDinst/reg_out_B_reg[19]  ( .DIN(\IDinst/N1043 ), .CLK(clk), 
        .CLRB(n813), .SETB(1'b1), .Q(reg_out_B[19]), .QN(n144) );
  dffascs1 \IDinst/reg_out_B_reg[18]  ( .DIN(\IDinst/N1042 ), .CLK(clk), 
        .CLRB(n812), .SETB(1'b1), .Q(reg_out_B[18]), .QN(n45) );
  dffascs1 \IDinst/reg_out_B_reg[17]  ( .DIN(\IDinst/N1041 ), .CLK(clk), 
        .CLRB(n817), .SETB(1'b1), .Q(reg_out_B[17]), .QN(n135) );
  dffascs1 \IDinst/reg_out_B_reg[16]  ( .DIN(\IDinst/N1040 ), .CLK(clk), 
        .CLRB(n922), .SETB(1'b1), .Q(reg_out_B[16]), .QN(n21) );
  dffascs1 \IDinst/reg_out_B_reg[15]  ( .DIN(\IDinst/N1039 ), .CLK(clk), 
        .CLRB(n821), .SETB(1'b1), .Q(reg_out_B[15]), .QN(n26) );
  dffascs1 \IDinst/reg_out_B_reg[14]  ( .DIN(\IDinst/N1038 ), .CLK(clk), 
        .CLRB(n820), .SETB(1'b1), .Q(reg_out_B[14]), .QN(n146) );
  dffascs1 \IDinst/reg_out_B_reg[13]  ( .DIN(\IDinst/N1037 ), .CLK(clk), 
        .CLRB(n812), .SETB(1'b1), .Q(reg_out_B[13]), .QN(n54) );
  dffascs1 \IDinst/reg_out_B_reg[12]  ( .DIN(\IDinst/N1036 ), .CLK(clk), 
        .CLRB(n914), .SETB(1'b1), .Q(reg_out_B[12]), .QN(n46) );
  dffascs1 \IDinst/reg_out_B_reg[11]  ( .DIN(\IDinst/N1035 ), .CLK(clk), 
        .CLRB(n892), .SETB(1'b1), .Q(reg_out_B[11]), .QN(n136) );
  dffascs1 \IDinst/reg_out_B_reg[10]  ( .DIN(\IDinst/N1034 ), .CLK(clk), 
        .CLRB(n828), .SETB(1'b1), .Q(reg_out_B[10]), .QN(n22) );
  dffascs1 \IDinst/reg_out_B_reg[9]  ( .DIN(\IDinst/N1033 ), .CLK(clk), 
        .CLRB(n860), .SETB(1'b1), .Q(reg_out_B[9]), .QN(n4) );
  dffascs1 \IDinst/reg_out_B_reg[8]  ( .DIN(\IDinst/N1032 ), .CLK(clk), 
        .CLRB(n895), .SETB(1'b1), .Q(reg_out_B[8]), .QN(n24) );
  dffascs1 \IDinst/reg_out_B_reg[7]  ( .DIN(\IDinst/N1031 ), .CLK(clk), 
        .CLRB(n828), .SETB(1'b1), .Q(reg_out_B[7]), .QN(n51) );
  dffascs1 \IDinst/reg_out_B_reg[6]  ( .DIN(\IDinst/N1030 ), .CLK(clk), 
        .CLRB(n829), .SETB(1'b1), .Q(reg_out_B[6]), .QN(n143) );
  dffascs1 \IDinst/reg_out_B_reg[5]  ( .DIN(\IDinst/N1029 ), .CLK(clk), 
        .CLRB(n853), .SETB(1'b1), .Q(reg_out_B[5]) );
  dffascs1 \IDinst/reg_out_B_reg[4]  ( .DIN(\IDinst/N1028 ), .CLK(clk), 
        .CLRB(n868), .SETB(1'b1), .Q(n55), .QN(n204) );
  dffascs1 \IDinst/reg_out_B_reg[3]  ( .DIN(\IDinst/N1027 ), .CLK(clk), 
        .CLRB(n841), .SETB(1'b1), .Q(n61), .QN(n337) );
  dffascs1 \IDinst/reg_out_B_reg[2]  ( .DIN(\IDinst/N1026 ), .CLK(clk), 
        .CLRB(n837), .SETB(1'b1), .Q(n32), .QN(n205) );
  dffascs1 \IDinst/reg_out_B_reg[1]  ( .DIN(\IDinst/N1025 ), .CLK(clk), 
        .CLRB(n829), .SETB(1'b1), .Q(reg_out_B[1]), .QN(n714) );
  dffascs1 \IDinst/reg_out_B_reg[0]  ( .DIN(\IDinst/N1024 ), .CLK(clk), 
        .CLRB(n963), .SETB(1'b1), .QN(n1) );
  dffascs1 \IDinst/branch_address_reg[31]  ( .DIN(\IDinst/n4793 ), .CLK(clk), 
        .CLRB(n809), .SETB(1'b1), .QN(n9406) );
  dffascs1 \IDinst/branch_address_reg[30]  ( .DIN(\IDinst/n4794 ), .CLK(clk), 
        .CLRB(n830), .SETB(1'b1), .Q(n263) );
  dffascs1 \IDinst/branch_address_reg[29]  ( .DIN(\IDinst/n4795 ), .CLK(clk), 
        .CLRB(n831), .SETB(1'b1), .Q(n262) );
  dffascs1 \IDinst/branch_address_reg[28]  ( .DIN(\IDinst/n4796 ), .CLK(clk), 
        .CLRB(n918), .SETB(1'b1), .Q(n261) );
  dffascs1 \IDinst/branch_address_reg[27]  ( .DIN(\IDinst/n4797 ), .CLK(clk), 
        .CLRB(n906), .SETB(1'b1), .Q(n260) );
  dffascs1 \IDinst/branch_address_reg[26]  ( .DIN(\IDinst/n4798 ), .CLK(clk), 
        .CLRB(n812), .SETB(1'b1), .Q(n259) );
  dffascs1 \IDinst/branch_address_reg[25]  ( .DIN(\IDinst/n4799 ), .CLK(clk), 
        .CLRB(n899), .SETB(1'b1), .Q(n258) );
  dffascs1 \IDinst/branch_address_reg[24]  ( .DIN(\IDinst/n4800 ), .CLK(clk), 
        .CLRB(n831), .SETB(1'b1), .Q(n257) );
  dffascs1 \IDinst/branch_address_reg[23]  ( .DIN(\IDinst/n4801 ), .CLK(clk), 
        .CLRB(n888), .SETB(1'b1), .Q(n256) );
  dffascs1 \IDinst/branch_address_reg[22]  ( .DIN(\IDinst/n4802 ), .CLK(clk), 
        .CLRB(n880), .SETB(1'b1), .Q(n255) );
  dffascs1 \IDinst/branch_address_reg[21]  ( .DIN(\IDinst/n4803 ), .CLK(clk), 
        .CLRB(n811), .SETB(1'b1), .Q(n254) );
  dffascs1 \IDinst/branch_address_reg[20]  ( .DIN(\IDinst/n4804 ), .CLK(clk), 
        .CLRB(n884), .SETB(1'b1), .Q(n253) );
  dffascs1 \IDinst/branch_address_reg[19]  ( .DIN(\IDinst/n4805 ), .CLK(clk), 
        .CLRB(n813), .SETB(1'b1), .Q(n252) );
  dffascs1 \IDinst/branch_address_reg[18]  ( .DIN(\IDinst/n4806 ), .CLK(clk), 
        .CLRB(n872), .SETB(1'b1), .Q(n251) );
  dffascs1 \IDinst/branch_address_reg[17]  ( .DIN(\IDinst/n4807 ), .CLK(clk), 
        .CLRB(n810), .SETB(1'b1), .Q(n250) );
  dffascs1 \IDinst/branch_address_reg[16]  ( .DIN(\IDinst/n4808 ), .CLK(clk), 
        .CLRB(n914), .SETB(1'b1), .Q(n249) );
  dffascs1 \IDinst/branch_address_reg[15]  ( .DIN(\IDinst/n4809 ), .CLK(clk), 
        .CLRB(n820), .SETB(1'b1), .Q(n248) );
  dffascs1 \IDinst/branch_address_reg[14]  ( .DIN(\IDinst/n4810 ), .CLK(clk), 
        .CLRB(n864), .SETB(1'b1), .Q(n247) );
  dffascs1 \IDinst/branch_address_reg[13]  ( .DIN(\IDinst/n4811 ), .CLK(clk), 
        .CLRB(n876), .SETB(1'b1), .Q(n246) );
  dffascs1 \IDinst/branch_address_reg[12]  ( .DIN(\IDinst/n4812 ), .CLK(clk), 
        .CLRB(n832), .SETB(1'b1), .Q(n245) );
  dffascs1 \IDinst/branch_address_reg[11]  ( .DIN(\IDinst/n4813 ), .CLK(clk), 
        .CLRB(n828), .SETB(1'b1), .Q(n244) );
  dffascs1 \IDinst/branch_address_reg[10]  ( .DIN(\IDinst/n4814 ), .CLK(clk), 
        .CLRB(n857), .SETB(1'b1), .Q(n243) );
  dffascs1 \IDinst/branch_address_reg[9]  ( .DIN(\IDinst/n4815 ), .CLK(clk), 
        .CLRB(n829), .SETB(1'b1), .Q(n242) );
  dffascs1 \IDinst/branch_address_reg[8]  ( .DIN(\IDinst/n4816 ), .CLK(clk), 
        .CLRB(n832), .SETB(1'b1), .Q(n241) );
  dffascs1 \IDinst/branch_address_reg[7]  ( .DIN(\IDinst/n4817 ), .CLK(clk), 
        .CLRB(n849), .SETB(1'b1), .Q(n240) );
  dffascs1 \IDinst/branch_address_reg[6]  ( .DIN(\IDinst/n4818 ), .CLK(clk), 
        .CLRB(n845), .SETB(1'b1), .Q(n239) );
  dffascs1 \IDinst/branch_address_reg[5]  ( .DIN(\IDinst/n4819 ), .CLK(clk), 
        .CLRB(n832), .SETB(1'b1), .Q(n238) );
  dffascs1 \IDinst/branch_address_reg[4]  ( .DIN(\IDinst/n4820 ), .CLK(clk), 
        .CLRB(n833), .SETB(1'b1), .Q(n237) );
  dffascs1 \IDinst/branch_address_reg[3]  ( .DIN(\IDinst/n4821 ), .CLK(clk), 
        .CLRB(n833), .SETB(1'b1), .Q(n236) );
  dffascs1 \IDinst/branch_address_reg[2]  ( .DIN(\IDinst/n4822 ), .CLK(clk), 
        .CLRB(n833), .SETB(1'b1), .Q(n235) );
  dffascs1 \IDinst/branch_address_reg[1]  ( .DIN(\IDinst/n4823 ), .CLK(clk), 
        .CLRB(n834), .SETB(1'b1), .Q(n234) );
  dffascs1 \IDinst/branch_address_reg[0]  ( .DIN(\IDinst/n4824 ), .CLK(clk), 
        .CLRB(n925), .SETB(1'b1), .Q(n233) );
  dffascs1 \IDinst/branch_sig_reg  ( .DIN(\IDinst/n4860 ), .CLK(clk), 
        .CLRB(n958), .SETB(1'b1), .QN(n9459) );
  dffascs1 \IDinst/EPC_reg[31]  ( .DIN(\IDinst/n4825 ), .CLK(clk), .CLRB(n918), 
        .SETB(1'b1), .Q(n156) );
  dffascs1 \IDinst/EPC_reg[30]  ( .DIN(\IDinst/n4826 ), .CLK(clk), .CLRB(n830), 
        .SETB(1'b1), .Q(n158) );
  dffascs1 \IDinst/EPC_reg[29]  ( .DIN(\IDinst/n4827 ), .CLK(clk), .CLRB(n831), 
        .SETB(1'b1), .Q(n160) );
  dffascs1 \IDinst/EPC_reg[28]  ( .DIN(\IDinst/n4828 ), .CLK(clk), .CLRB(n918), 
        .SETB(1'b1), .Q(n162) );
  dffascs1 \IDinst/EPC_reg[27]  ( .DIN(\IDinst/n4829 ), .CLK(clk), .CLRB(n906), 
        .SETB(1'b1), .Q(n164) );
  dffascs1 \IDinst/EPC_reg[26]  ( .DIN(\IDinst/n4830 ), .CLK(clk), .CLRB(n879), 
        .SETB(1'b1), .Q(n166) );
  dffascs1 \IDinst/EPC_reg[25]  ( .DIN(\IDinst/n4831 ), .CLK(clk), .CLRB(n899), 
        .SETB(1'b1), .Q(n168) );
  dffascs1 \IDinst/EPC_reg[24]  ( .DIN(\IDinst/n4832 ), .CLK(clk), .CLRB(n880), 
        .SETB(1'b1), .Q(n170) );
  dffascs1 \IDinst/EPC_reg[23]  ( .DIN(\IDinst/n4833 ), .CLK(clk), .CLRB(n888), 
        .SETB(1'b1), .Q(n172) );
  dffascs1 \IDinst/EPC_reg[22]  ( .DIN(\IDinst/n4834 ), .CLK(clk), .CLRB(n880), 
        .SETB(1'b1), .Q(n174) );
  dffascs1 \IDinst/EPC_reg[21]  ( .DIN(\IDinst/n4835 ), .CLK(clk), .CLRB(n884), 
        .SETB(1'b1), .Q(n176) );
  dffascs1 \IDinst/EPC_reg[20]  ( .DIN(\IDinst/n4836 ), .CLK(clk), .CLRB(n884), 
        .SETB(1'b1), .Q(n178) );
  dffascs1 \IDinst/EPC_reg[19]  ( .DIN(\IDinst/n4837 ), .CLK(clk), .CLRB(n871), 
        .SETB(1'b1), .Q(n180) );
  dffascs1 \IDinst/EPC_reg[18]  ( .DIN(\IDinst/n4838 ), .CLK(clk), .CLRB(n872), 
        .SETB(1'b1), .Q(n182) );
  dffascs1 \IDinst/EPC_reg[17]  ( .DIN(\IDinst/n4839 ), .CLK(clk), .CLRB(n913), 
        .SETB(1'b1), .Q(n184) );
  dffascs1 \IDinst/EPC_reg[16]  ( .DIN(\IDinst/n4840 ), .CLK(clk), .CLRB(n914), 
        .SETB(1'b1), .Q(n186) );
  dffascs1 \IDinst/EPC_reg[15]  ( .DIN(\IDinst/n4841 ), .CLK(clk), .CLRB(n864), 
        .SETB(1'b1), .Q(n187) );
  dffascs1 \IDinst/EPC_reg[14]  ( .DIN(\IDinst/n4842 ), .CLK(clk), .CLRB(n864), 
        .SETB(1'b1), .Q(n189) );
  dffascs1 \IDinst/EPC_reg[13]  ( .DIN(\IDinst/n4843 ), .CLK(clk), .CLRB(n876), 
        .SETB(1'b1), .Q(n191) );
  dffascs1 \IDinst/EPC_reg[12]  ( .DIN(\IDinst/n4844 ), .CLK(clk), .CLRB(n831), 
        .SETB(1'b1), .Q(n193) );
  dffascs1 \IDinst/EPC_reg[11]  ( .DIN(\IDinst/n4845 ), .CLK(clk), .CLRB(n856), 
        .SETB(1'b1), .Q(n195) );
  dffascs1 \IDinst/EPC_reg[10]  ( .DIN(\IDinst/n4846 ), .CLK(clk), .CLRB(n856), 
        .SETB(1'b1), .Q(n197) );
  dffascs1 \IDinst/EPC_reg[9]  ( .DIN(\IDinst/n4847 ), .CLK(clk), .CLRB(n844), 
        .SETB(1'b1), .Q(n199) );
  dffascs1 \IDinst/EPC_reg[8]  ( .DIN(\IDinst/n4848 ), .CLK(clk), .CLRB(n845), 
        .SETB(1'b1), .Q(n201) );
  dffascs1 \IDinst/EPC_reg[7]  ( .DIN(\IDinst/n4849 ), .CLK(clk), .CLRB(n849), 
        .SETB(1'b1), .Q(n147) );
  dffascs1 \IDinst/EPC_reg[6]  ( .DIN(\IDinst/n4850 ), .CLK(clk), .CLRB(n845), 
        .SETB(1'b1), .Q(n148) );
  dffascs1 \IDinst/EPC_reg[5]  ( .DIN(\IDinst/n4851 ), .CLK(clk), .CLRB(n832), 
        .SETB(1'b1), .Q(n149) );
  dffascs1 \IDinst/EPC_reg[4]  ( .DIN(\IDinst/n4852 ), .CLK(clk), .CLRB(n832), 
        .SETB(1'b1), .Q(n150) );
  dffascs1 \IDinst/EPC_reg[3]  ( .DIN(\IDinst/n4853 ), .CLK(clk), .CLRB(n833), 
        .SETB(1'b1), .Q(n151) );
  dffascs1 \IDinst/EPC_reg[2]  ( .DIN(\IDinst/n4854 ), .CLK(clk), .CLRB(n830), 
        .SETB(1'b1), .Q(n152) );
  dffascs1 \IDinst/EPC_reg[1]  ( .DIN(\IDinst/n4855 ), .CLK(clk), .CLRB(n830), 
        .SETB(1'b1), .Q(n153) );
  dffascs1 \IDinst/EPC_reg[0]  ( .DIN(\IDinst/n4856 ), .CLK(clk), .CLRB(n926), 
        .SETB(1'b1), .Q(n154) );
  dffascs1 \IDinst/CLI_reg  ( .DIN(\IDinst/n5947 ), .CLK(clk), .CLRB(n951), 
        .SETB(1'b1), .Q(CLI), .QN(\IDinst/n1444 ) );
  dffascs1 \IDinst/RegFile_reg[0][15]  ( .DIN(\IDinst/n5420 ), .CLK(clk), 
        .CLRB(n821), .SETB(1'b1), .Q(\IDinst/RegFile[0][15] ) );
  dffascs1 \IDinst/RegFile_reg[1][15]  ( .DIN(\IDinst/n5419 ), .CLK(clk), 
        .CLRB(n821), .SETB(1'b1), .Q(\IDinst/RegFile[1][15] ) );
  dffascs1 \IDinst/RegFile_reg[2][15]  ( .DIN(\IDinst/n5418 ), .CLK(clk), 
        .CLRB(n821), .SETB(1'b1), .Q(\IDinst/RegFile[2][15] ) );
  dffascs1 \IDinst/RegFile_reg[3][15]  ( .DIN(\IDinst/n5417 ), .CLK(clk), 
        .CLRB(n821), .SETB(1'b1), .Q(\IDinst/RegFile[3][15] ) );
  dffascs1 \IDinst/RegFile_reg[4][15]  ( .DIN(\IDinst/n5416 ), .CLK(clk), 
        .CLRB(n821), .SETB(1'b1), .Q(\IDinst/RegFile[4][15] ) );
  dffascs1 \IDinst/RegFile_reg[5][15]  ( .DIN(\IDinst/n5415 ), .CLK(clk), 
        .CLRB(n821), .SETB(1'b1), .Q(\IDinst/RegFile[5][15] ) );
  dffascs1 \IDinst/RegFile_reg[6][15]  ( .DIN(\IDinst/n5414 ), .CLK(clk), 
        .CLRB(n821), .SETB(1'b1), .Q(\IDinst/RegFile[6][15] ) );
  dffascs1 \IDinst/RegFile_reg[7][15]  ( .DIN(\IDinst/n5413 ), .CLK(clk), 
        .CLRB(n821), .SETB(1'b1), .Q(\IDinst/RegFile[7][15] ) );
  dffascs1 \IDinst/RegFile_reg[8][15]  ( .DIN(\IDinst/n5412 ), .CLK(clk), 
        .CLRB(n822), .SETB(1'b1), .Q(\IDinst/RegFile[8][15] ) );
  dffascs1 \IDinst/RegFile_reg[9][15]  ( .DIN(\IDinst/n5411 ), .CLK(clk), 
        .CLRB(n822), .SETB(1'b1), .Q(\IDinst/RegFile[9][15] ) );
  dffascs1 \IDinst/RegFile_reg[10][15]  ( .DIN(\IDinst/n5410 ), .CLK(clk), 
        .CLRB(n822), .SETB(1'b1), .Q(\IDinst/RegFile[10][15] ) );
  dffascs1 \IDinst/RegFile_reg[11][15]  ( .DIN(\IDinst/n5409 ), .CLK(clk), 
        .CLRB(n822), .SETB(1'b1), .Q(\IDinst/RegFile[11][15] ) );
  dffascs1 \IDinst/RegFile_reg[12][15]  ( .DIN(\IDinst/n5408 ), .CLK(clk), 
        .CLRB(n822), .SETB(1'b1), .Q(\IDinst/RegFile[12][15] ) );
  dffascs1 \IDinst/RegFile_reg[13][15]  ( .DIN(\IDinst/n5407 ), .CLK(clk), 
        .CLRB(n822), .SETB(1'b1), .Q(\IDinst/RegFile[13][15] ) );
  dffascs1 \IDinst/RegFile_reg[14][15]  ( .DIN(\IDinst/n5406 ), .CLK(clk), 
        .CLRB(n822), .SETB(1'b1), .Q(\IDinst/RegFile[14][15] ) );
  dffascs1 \IDinst/RegFile_reg[15][15]  ( .DIN(\IDinst/n5405 ), .CLK(clk), 
        .CLRB(n822), .SETB(1'b1), .Q(\IDinst/RegFile[15][15] ) );
  dffascs1 \IDinst/RegFile_reg[16][15]  ( .DIN(\IDinst/n5404 ), .CLK(clk), 
        .CLRB(n822), .SETB(1'b1), .Q(\IDinst/RegFile[16][15] ) );
  dffascs1 \IDinst/RegFile_reg[17][15]  ( .DIN(\IDinst/n5403 ), .CLK(clk), 
        .CLRB(n822), .SETB(1'b1), .Q(\IDinst/RegFile[17][15] ) );
  dffascs1 \IDinst/RegFile_reg[18][15]  ( .DIN(\IDinst/n5402 ), .CLK(clk), 
        .CLRB(n823), .SETB(1'b1), .Q(\IDinst/RegFile[18][15] ) );
  dffascs1 \IDinst/RegFile_reg[19][15]  ( .DIN(\IDinst/n5401 ), .CLK(clk), 
        .CLRB(n823), .SETB(1'b1), .Q(\IDinst/RegFile[19][15] ) );
  dffascs1 \IDinst/RegFile_reg[20][15]  ( .DIN(\IDinst/n5400 ), .CLK(clk), 
        .CLRB(n823), .SETB(1'b1), .Q(\IDinst/RegFile[20][15] ) );
  dffascs1 \IDinst/RegFile_reg[21][15]  ( .DIN(\IDinst/n5399 ), .CLK(clk), 
        .CLRB(n823), .SETB(1'b1), .Q(\IDinst/RegFile[21][15] ) );
  dffascs1 \IDinst/RegFile_reg[22][15]  ( .DIN(\IDinst/n5398 ), .CLK(clk), 
        .CLRB(n823), .SETB(1'b1), .Q(\IDinst/RegFile[22][15] ) );
  dffascs1 \IDinst/RegFile_reg[23][15]  ( .DIN(\IDinst/n5397 ), .CLK(clk), 
        .CLRB(n823), .SETB(1'b1), .Q(\IDinst/RegFile[23][15] ) );
  dffascs1 \IDinst/RegFile_reg[24][15]  ( .DIN(\IDinst/n5396 ), .CLK(clk), 
        .CLRB(n823), .SETB(1'b1), .Q(\IDinst/RegFile[24][15] ) );
  dffascs1 \IDinst/RegFile_reg[25][15]  ( .DIN(\IDinst/n5395 ), .CLK(clk), 
        .CLRB(n823), .SETB(1'b1), .Q(\IDinst/RegFile[25][15] ) );
  dffascs1 \IDinst/RegFile_reg[26][15]  ( .DIN(\IDinst/n5394 ), .CLK(clk), 
        .CLRB(n823), .SETB(1'b1), .Q(\IDinst/RegFile[26][15] ) );
  dffascs1 \IDinst/RegFile_reg[27][15]  ( .DIN(\IDinst/n5393 ), .CLK(clk), 
        .CLRB(n823), .SETB(1'b1), .Q(\IDinst/RegFile[27][15] ) );
  dffascs1 \IDinst/RegFile_reg[28][15]  ( .DIN(\IDinst/n5392 ), .CLK(clk), 
        .CLRB(n824), .SETB(1'b1), .Q(\IDinst/RegFile[28][15] ) );
  dffascs1 \IDinst/RegFile_reg[29][15]  ( .DIN(\IDinst/n5391 ), .CLK(clk), 
        .CLRB(n824), .SETB(1'b1), .Q(\IDinst/RegFile[29][15] ) );
  dffascs1 \IDinst/RegFile_reg[30][15]  ( .DIN(\IDinst/n5390 ), .CLK(clk), 
        .CLRB(n824), .SETB(1'b1), .Q(\IDinst/RegFile[30][15] ) );
  dffascs1 \IDinst/RegFile_reg[31][15]  ( .DIN(\IDinst/n5389 ), .CLK(clk), 
        .CLRB(n824), .SETB(1'b1), .Q(\IDinst/RegFile[31][15] ) );
  dffascs1 \IDinst/RegFile_reg[0][16]  ( .DIN(\IDinst/n5388 ), .CLK(clk), 
        .CLRB(n922), .SETB(1'b1), .Q(\IDinst/RegFile[0][16] ) );
  dffascs1 \IDinst/RegFile_reg[1][16]  ( .DIN(\IDinst/n5387 ), .CLK(clk), 
        .CLRB(n922), .SETB(1'b1), .Q(\IDinst/RegFile[1][16] ) );
  dffascs1 \IDinst/RegFile_reg[2][16]  ( .DIN(\IDinst/n5386 ), .CLK(clk), 
        .CLRB(n922), .SETB(1'b1), .Q(\IDinst/RegFile[2][16] ) );
  dffascs1 \IDinst/RegFile_reg[3][16]  ( .DIN(\IDinst/n5385 ), .CLK(clk), 
        .CLRB(n922), .SETB(1'b1), .Q(\IDinst/RegFile[3][16] ) );
  dffascs1 \IDinst/RegFile_reg[4][16]  ( .DIN(\IDinst/n5384 ), .CLK(clk), 
        .CLRB(n922), .SETB(1'b1), .Q(\IDinst/RegFile[4][16] ) );
  dffascs1 \IDinst/RegFile_reg[5][16]  ( .DIN(\IDinst/n5383 ), .CLK(clk), 
        .CLRB(n923), .SETB(1'b1), .Q(\IDinst/RegFile[5][16] ) );
  dffascs1 \IDinst/RegFile_reg[6][16]  ( .DIN(\IDinst/n5382 ), .CLK(clk), 
        .CLRB(n923), .SETB(1'b1), .Q(\IDinst/RegFile[6][16] ) );
  dffascs1 \IDinst/RegFile_reg[7][16]  ( .DIN(\IDinst/n5381 ), .CLK(clk), 
        .CLRB(n923), .SETB(1'b1), .Q(\IDinst/RegFile[7][16] ) );
  dffascs1 \IDinst/RegFile_reg[8][16]  ( .DIN(\IDinst/n5380 ), .CLK(clk), 
        .CLRB(n923), .SETB(1'b1), .Q(\IDinst/RegFile[8][16] ) );
  dffascs1 \IDinst/RegFile_reg[9][16]  ( .DIN(\IDinst/n5379 ), .CLK(clk), 
        .CLRB(n923), .SETB(1'b1), .Q(\IDinst/RegFile[9][16] ) );
  dffascs1 \IDinst/RegFile_reg[10][16]  ( .DIN(\IDinst/n5378 ), .CLK(clk), 
        .CLRB(n923), .SETB(1'b1), .Q(\IDinst/RegFile[10][16] ) );
  dffascs1 \IDinst/RegFile_reg[11][16]  ( .DIN(\IDinst/n5377 ), .CLK(clk), 
        .CLRB(n923), .SETB(1'b1), .Q(\IDinst/RegFile[11][16] ) );
  dffascs1 \IDinst/RegFile_reg[12][16]  ( .DIN(\IDinst/n5376 ), .CLK(clk), 
        .CLRB(n923), .SETB(1'b1), .Q(\IDinst/RegFile[12][16] ) );
  dffascs1 \IDinst/RegFile_reg[13][16]  ( .DIN(\IDinst/n5375 ), .CLK(clk), 
        .CLRB(n923), .SETB(1'b1), .Q(\IDinst/RegFile[13][16] ) );
  dffascs1 \IDinst/RegFile_reg[14][16]  ( .DIN(\IDinst/n5374 ), .CLK(clk), 
        .CLRB(n923), .SETB(1'b1), .Q(\IDinst/RegFile[14][16] ) );
  dffascs1 \IDinst/RegFile_reg[15][16]  ( .DIN(\IDinst/n5373 ), .CLK(clk), 
        .CLRB(n924), .SETB(1'b1), .Q(\IDinst/RegFile[15][16] ) );
  dffascs1 \IDinst/RegFile_reg[16][16]  ( .DIN(\IDinst/n5372 ), .CLK(clk), 
        .CLRB(n924), .SETB(1'b1), .Q(\IDinst/RegFile[16][16] ) );
  dffascs1 \IDinst/RegFile_reg[17][16]  ( .DIN(\IDinst/n5371 ), .CLK(clk), 
        .CLRB(n924), .SETB(1'b1), .Q(\IDinst/RegFile[17][16] ) );
  dffascs1 \IDinst/RegFile_reg[18][16]  ( .DIN(\IDinst/n5370 ), .CLK(clk), 
        .CLRB(n924), .SETB(1'b1), .Q(\IDinst/RegFile[18][16] ) );
  dffascs1 \IDinst/RegFile_reg[19][16]  ( .DIN(\IDinst/n5369 ), .CLK(clk), 
        .CLRB(n924), .SETB(1'b1), .Q(\IDinst/RegFile[19][16] ) );
  dffascs1 \IDinst/RegFile_reg[20][16]  ( .DIN(\IDinst/n5368 ), .CLK(clk), 
        .CLRB(n924), .SETB(1'b1), .Q(\IDinst/RegFile[20][16] ) );
  dffascs1 \IDinst/RegFile_reg[21][16]  ( .DIN(\IDinst/n5367 ), .CLK(clk), 
        .CLRB(n924), .SETB(1'b1), .Q(\IDinst/RegFile[21][16] ) );
  dffascs1 \IDinst/RegFile_reg[22][16]  ( .DIN(\IDinst/n5366 ), .CLK(clk), 
        .CLRB(n924), .SETB(1'b1), .Q(\IDinst/RegFile[22][16] ) );
  dffascs1 \IDinst/RegFile_reg[23][16]  ( .DIN(\IDinst/n5365 ), .CLK(clk), 
        .CLRB(n924), .SETB(1'b1), .Q(\IDinst/RegFile[23][16] ) );
  dffascs1 \IDinst/RegFile_reg[24][16]  ( .DIN(\IDinst/n5364 ), .CLK(clk), 
        .CLRB(n924), .SETB(1'b1), .Q(\IDinst/RegFile[24][16] ) );
  dffascs1 \IDinst/RegFile_reg[25][16]  ( .DIN(\IDinst/n5363 ), .CLK(clk), 
        .CLRB(n925), .SETB(1'b1), .Q(\IDinst/RegFile[25][16] ) );
  dffascs1 \IDinst/RegFile_reg[26][16]  ( .DIN(\IDinst/n5362 ), .CLK(clk), 
        .CLRB(n925), .SETB(1'b1), .Q(\IDinst/RegFile[26][16] ) );
  dffascs1 \IDinst/RegFile_reg[27][16]  ( .DIN(\IDinst/n5361 ), .CLK(clk), 
        .CLRB(n925), .SETB(1'b1), .Q(\IDinst/RegFile[27][16] ) );
  dffascs1 \IDinst/RegFile_reg[28][16]  ( .DIN(\IDinst/n5360 ), .CLK(clk), 
        .CLRB(n925), .SETB(1'b1), .Q(\IDinst/RegFile[28][16] ) );
  dffascs1 \IDinst/RegFile_reg[29][16]  ( .DIN(\IDinst/n5359 ), .CLK(clk), 
        .CLRB(n925), .SETB(1'b1), .Q(\IDinst/RegFile[29][16] ) );
  dffascs1 \IDinst/RegFile_reg[30][16]  ( .DIN(\IDinst/n5358 ), .CLK(clk), 
        .CLRB(n925), .SETB(1'b1), .Q(\IDinst/RegFile[30][16] ) );
  dffascs1 \IDinst/RegFile_reg[31][16]  ( .DIN(\IDinst/n5357 ), .CLK(clk), 
        .CLRB(n925), .SETB(1'b1), .Q(\IDinst/RegFile[31][16] ) );
  dffascs1 \IDinst/RegFile_reg[0][17]  ( .DIN(\IDinst/n5356 ), .CLK(clk), 
        .CLRB(n817), .SETB(1'b1), .Q(\IDinst/RegFile[0][17] ) );
  dffascs1 \IDinst/RegFile_reg[1][17]  ( .DIN(\IDinst/n5355 ), .CLK(clk), 
        .CLRB(n817), .SETB(1'b1), .Q(\IDinst/RegFile[1][17] ) );
  dffascs1 \IDinst/RegFile_reg[2][17]  ( .DIN(\IDinst/n5354 ), .CLK(clk), 
        .CLRB(n817), .SETB(1'b1), .Q(\IDinst/RegFile[2][17] ) );
  dffascs1 \IDinst/RegFile_reg[3][17]  ( .DIN(\IDinst/n5353 ), .CLK(clk), 
        .CLRB(n817), .SETB(1'b1), .Q(\IDinst/RegFile[3][17] ) );
  dffascs1 \IDinst/RegFile_reg[4][17]  ( .DIN(\IDinst/n5352 ), .CLK(clk), 
        .CLRB(n817), .SETB(1'b1), .Q(\IDinst/RegFile[4][17] ) );
  dffascs1 \IDinst/RegFile_reg[5][17]  ( .DIN(\IDinst/n5351 ), .CLK(clk), 
        .CLRB(n817), .SETB(1'b1), .Q(\IDinst/RegFile[5][17] ) );
  dffascs1 \IDinst/RegFile_reg[6][17]  ( .DIN(\IDinst/n5350 ), .CLK(clk), 
        .CLRB(n817), .SETB(1'b1), .Q(\IDinst/RegFile[6][17] ) );
  dffascs1 \IDinst/RegFile_reg[7][17]  ( .DIN(\IDinst/n5349 ), .CLK(clk), 
        .CLRB(n817), .SETB(1'b1), .Q(\IDinst/RegFile[7][17] ) );
  dffascs1 \IDinst/RegFile_reg[8][17]  ( .DIN(\IDinst/n5348 ), .CLK(clk), 
        .CLRB(n817), .SETB(1'b1), .Q(\IDinst/RegFile[8][17] ) );
  dffascs1 \IDinst/RegFile_reg[9][17]  ( .DIN(\IDinst/n5347 ), .CLK(clk), 
        .CLRB(n818), .SETB(1'b1), .Q(\IDinst/RegFile[9][17] ) );
  dffascs1 \IDinst/RegFile_reg[10][17]  ( .DIN(\IDinst/n5346 ), .CLK(clk), 
        .CLRB(n818), .SETB(1'b1), .Q(\IDinst/RegFile[10][17] ) );
  dffascs1 \IDinst/RegFile_reg[11][17]  ( .DIN(\IDinst/n5345 ), .CLK(clk), 
        .CLRB(n818), .SETB(1'b1), .Q(\IDinst/RegFile[11][17] ) );
  dffascs1 \IDinst/RegFile_reg[12][17]  ( .DIN(\IDinst/n5344 ), .CLK(clk), 
        .CLRB(n818), .SETB(1'b1), .Q(\IDinst/RegFile[12][17] ) );
  dffascs1 \IDinst/RegFile_reg[13][17]  ( .DIN(\IDinst/n5343 ), .CLK(clk), 
        .CLRB(n818), .SETB(1'b1), .Q(\IDinst/RegFile[13][17] ) );
  dffascs1 \IDinst/RegFile_reg[14][17]  ( .DIN(\IDinst/n5342 ), .CLK(clk), 
        .CLRB(n818), .SETB(1'b1), .Q(\IDinst/RegFile[14][17] ) );
  dffascs1 \IDinst/RegFile_reg[15][17]  ( .DIN(\IDinst/n5341 ), .CLK(clk), 
        .CLRB(n818), .SETB(1'b1), .Q(\IDinst/RegFile[15][17] ) );
  dffascs1 \IDinst/RegFile_reg[16][17]  ( .DIN(\IDinst/n5340 ), .CLK(clk), 
        .CLRB(n818), .SETB(1'b1), .Q(\IDinst/RegFile[16][17] ) );
  dffascs1 \IDinst/RegFile_reg[17][17]  ( .DIN(\IDinst/n5339 ), .CLK(clk), 
        .CLRB(n818), .SETB(1'b1), .Q(\IDinst/RegFile[17][17] ) );
  dffascs1 \IDinst/RegFile_reg[18][17]  ( .DIN(\IDinst/n5338 ), .CLK(clk), 
        .CLRB(n818), .SETB(1'b1), .Q(\IDinst/RegFile[18][17] ) );
  dffascs1 \IDinst/RegFile_reg[19][17]  ( .DIN(\IDinst/n5337 ), .CLK(clk), 
        .CLRB(n819), .SETB(1'b1), .Q(\IDinst/RegFile[19][17] ) );
  dffascs1 \IDinst/RegFile_reg[20][17]  ( .DIN(\IDinst/n5336 ), .CLK(clk), 
        .CLRB(n819), .SETB(1'b1), .Q(\IDinst/RegFile[20][17] ) );
  dffascs1 \IDinst/RegFile_reg[21][17]  ( .DIN(\IDinst/n5335 ), .CLK(clk), 
        .CLRB(n819), .SETB(1'b1), .Q(\IDinst/RegFile[21][17] ) );
  dffascs1 \IDinst/RegFile_reg[22][17]  ( .DIN(\IDinst/n5334 ), .CLK(clk), 
        .CLRB(n819), .SETB(1'b1), .Q(\IDinst/RegFile[22][17] ) );
  dffascs1 \IDinst/RegFile_reg[23][17]  ( .DIN(\IDinst/n5333 ), .CLK(clk), 
        .CLRB(n819), .SETB(1'b1), .Q(\IDinst/RegFile[23][17] ) );
  dffascs1 \IDinst/RegFile_reg[24][17]  ( .DIN(\IDinst/n5332 ), .CLK(clk), 
        .CLRB(n819), .SETB(1'b1), .Q(\IDinst/RegFile[24][17] ) );
  dffascs1 \IDinst/RegFile_reg[25][17]  ( .DIN(\IDinst/n5331 ), .CLK(clk), 
        .CLRB(n819), .SETB(1'b1), .Q(\IDinst/RegFile[25][17] ) );
  dffascs1 \IDinst/RegFile_reg[26][17]  ( .DIN(\IDinst/n5330 ), .CLK(clk), 
        .CLRB(n819), .SETB(1'b1), .Q(\IDinst/RegFile[26][17] ) );
  dffascs1 \IDinst/RegFile_reg[27][17]  ( .DIN(\IDinst/n5329 ), .CLK(clk), 
        .CLRB(n819), .SETB(1'b1), .Q(\IDinst/RegFile[27][17] ) );
  dffascs1 \IDinst/RegFile_reg[28][17]  ( .DIN(\IDinst/n5328 ), .CLK(clk), 
        .CLRB(n819), .SETB(1'b1), .Q(\IDinst/RegFile[28][17] ) );
  dffascs1 \IDinst/RegFile_reg[29][17]  ( .DIN(\IDinst/n5327 ), .CLK(clk), 
        .CLRB(n820), .SETB(1'b1), .Q(\IDinst/RegFile[29][17] ) );
  dffascs1 \IDinst/RegFile_reg[30][17]  ( .DIN(\IDinst/n5326 ), .CLK(clk), 
        .CLRB(n820), .SETB(1'b1), .Q(\IDinst/RegFile[30][17] ) );
  dffascs1 \IDinst/RegFile_reg[31][17]  ( .DIN(\IDinst/n5325 ), .CLK(clk), 
        .CLRB(n820), .SETB(1'b1), .Q(\IDinst/RegFile[31][17] ) );
  dffascs1 \IDinst/RegFile_reg[0][18]  ( .DIN(\IDinst/n5324 ), .CLK(clk), 
        .CLRB(n872), .SETB(1'b1), .Q(\IDinst/RegFile[0][18] ) );
  dffascs1 \IDinst/RegFile_reg[1][18]  ( .DIN(\IDinst/n5323 ), .CLK(clk), 
        .CLRB(n872), .SETB(1'b1), .Q(\IDinst/RegFile[1][18] ) );
  dffascs1 \IDinst/RegFile_reg[2][18]  ( .DIN(\IDinst/n5322 ), .CLK(clk), 
        .CLRB(n872), .SETB(1'b1), .Q(\IDinst/RegFile[2][18] ) );
  dffascs1 \IDinst/RegFile_reg[3][18]  ( .DIN(\IDinst/n5321 ), .CLK(clk), 
        .CLRB(n872), .SETB(1'b1), .Q(\IDinst/RegFile[3][18] ) );
  dffascs1 \IDinst/RegFile_reg[4][18]  ( .DIN(\IDinst/n5320 ), .CLK(clk), 
        .CLRB(n872), .SETB(1'b1), .Q(\IDinst/RegFile[4][18] ) );
  dffascs1 \IDinst/RegFile_reg[5][18]  ( .DIN(\IDinst/n5319 ), .CLK(clk), 
        .CLRB(n873), .SETB(1'b1), .Q(\IDinst/RegFile[5][18] ) );
  dffascs1 \IDinst/RegFile_reg[6][18]  ( .DIN(\IDinst/n5318 ), .CLK(clk), 
        .CLRB(n873), .SETB(1'b1), .Q(\IDinst/RegFile[6][18] ) );
  dffascs1 \IDinst/RegFile_reg[7][18]  ( .DIN(\IDinst/n5317 ), .CLK(clk), 
        .CLRB(n873), .SETB(1'b1), .Q(\IDinst/RegFile[7][18] ) );
  dffascs1 \IDinst/RegFile_reg[8][18]  ( .DIN(\IDinst/n5316 ), .CLK(clk), 
        .CLRB(n873), .SETB(1'b1), .Q(\IDinst/RegFile[8][18] ) );
  dffascs1 \IDinst/RegFile_reg[9][18]  ( .DIN(\IDinst/n5315 ), .CLK(clk), 
        .CLRB(n873), .SETB(1'b1), .Q(\IDinst/RegFile[9][18] ) );
  dffascs1 \IDinst/RegFile_reg[10][18]  ( .DIN(\IDinst/n5314 ), .CLK(clk), 
        .CLRB(n873), .SETB(1'b1), .Q(\IDinst/RegFile[10][18] ) );
  dffascs1 \IDinst/RegFile_reg[11][18]  ( .DIN(\IDinst/n5313 ), .CLK(clk), 
        .CLRB(n873), .SETB(1'b1), .Q(\IDinst/RegFile[11][18] ) );
  dffascs1 \IDinst/RegFile_reg[12][18]  ( .DIN(\IDinst/n5312 ), .CLK(clk), 
        .CLRB(n873), .SETB(1'b1), .Q(\IDinst/RegFile[12][18] ) );
  dffascs1 \IDinst/RegFile_reg[13][18]  ( .DIN(\IDinst/n5311 ), .CLK(clk), 
        .CLRB(n873), .SETB(1'b1), .Q(\IDinst/RegFile[13][18] ) );
  dffascs1 \IDinst/RegFile_reg[14][18]  ( .DIN(\IDinst/n5310 ), .CLK(clk), 
        .CLRB(n873), .SETB(1'b1), .Q(\IDinst/RegFile[14][18] ) );
  dffascs1 \IDinst/RegFile_reg[15][18]  ( .DIN(\IDinst/n5309 ), .CLK(clk), 
        .CLRB(n874), .SETB(1'b1), .Q(\IDinst/RegFile[15][18] ) );
  dffascs1 \IDinst/RegFile_reg[16][18]  ( .DIN(\IDinst/n5308 ), .CLK(clk), 
        .CLRB(n874), .SETB(1'b1), .Q(\IDinst/RegFile[16][18] ) );
  dffascs1 \IDinst/RegFile_reg[17][18]  ( .DIN(\IDinst/n5307 ), .CLK(clk), 
        .CLRB(n874), .SETB(1'b1), .Q(\IDinst/RegFile[17][18] ) );
  dffascs1 \IDinst/RegFile_reg[18][18]  ( .DIN(\IDinst/n5306 ), .CLK(clk), 
        .CLRB(n874), .SETB(1'b1), .Q(\IDinst/RegFile[18][18] ) );
  dffascs1 \IDinst/RegFile_reg[19][18]  ( .DIN(\IDinst/n5305 ), .CLK(clk), 
        .CLRB(n874), .SETB(1'b1), .Q(\IDinst/RegFile[19][18] ) );
  dffascs1 \IDinst/RegFile_reg[20][18]  ( .DIN(\IDinst/n5304 ), .CLK(clk), 
        .CLRB(n874), .SETB(1'b1), .Q(\IDinst/RegFile[20][18] ) );
  dffascs1 \IDinst/RegFile_reg[21][18]  ( .DIN(\IDinst/n5303 ), .CLK(clk), 
        .CLRB(n874), .SETB(1'b1), .Q(\IDinst/RegFile[21][18] ) );
  dffascs1 \IDinst/RegFile_reg[22][18]  ( .DIN(\IDinst/n5302 ), .CLK(clk), 
        .CLRB(n874), .SETB(1'b1), .Q(\IDinst/RegFile[22][18] ) );
  dffascs1 \IDinst/RegFile_reg[23][18]  ( .DIN(\IDinst/n5301 ), .CLK(clk), 
        .CLRB(n874), .SETB(1'b1), .Q(\IDinst/RegFile[23][18] ) );
  dffascs1 \IDinst/RegFile_reg[24][18]  ( .DIN(\IDinst/n5300 ), .CLK(clk), 
        .CLRB(n874), .SETB(1'b1), .Q(\IDinst/RegFile[24][18] ) );
  dffascs1 \IDinst/RegFile_reg[25][18]  ( .DIN(\IDinst/n5299 ), .CLK(clk), 
        .CLRB(n875), .SETB(1'b1), .Q(\IDinst/RegFile[25][18] ) );
  dffascs1 \IDinst/RegFile_reg[26][18]  ( .DIN(\IDinst/n5298 ), .CLK(clk), 
        .CLRB(n875), .SETB(1'b1), .Q(\IDinst/RegFile[26][18] ) );
  dffascs1 \IDinst/RegFile_reg[27][18]  ( .DIN(\IDinst/n5297 ), .CLK(clk), 
        .CLRB(n875), .SETB(1'b1), .Q(\IDinst/RegFile[27][18] ) );
  dffascs1 \IDinst/RegFile_reg[28][18]  ( .DIN(\IDinst/n5296 ), .CLK(clk), 
        .CLRB(n875), .SETB(1'b1), .Q(\IDinst/RegFile[28][18] ) );
  dffascs1 \IDinst/RegFile_reg[29][18]  ( .DIN(\IDinst/n5295 ), .CLK(clk), 
        .CLRB(n875), .SETB(1'b1), .Q(\IDinst/RegFile[29][18] ) );
  dffascs1 \IDinst/RegFile_reg[30][18]  ( .DIN(\IDinst/n5294 ), .CLK(clk), 
        .CLRB(n875), .SETB(1'b1), .Q(\IDinst/RegFile[30][18] ) );
  dffascs1 \IDinst/RegFile_reg[31][18]  ( .DIN(\IDinst/n5293 ), .CLK(clk), 
        .CLRB(n875), .SETB(1'b1), .Q(\IDinst/RegFile[31][18] ) );
  dffascs1 \IDinst/RegFile_reg[0][19]  ( .DIN(\IDinst/n5292 ), .CLK(clk), 
        .CLRB(n813), .SETB(1'b1), .Q(\IDinst/RegFile[0][19] ) );
  dffascs1 \IDinst/RegFile_reg[1][19]  ( .DIN(\IDinst/n5291 ), .CLK(clk), 
        .CLRB(n813), .SETB(1'b1), .Q(\IDinst/RegFile[1][19] ) );
  dffascs1 \IDinst/RegFile_reg[2][19]  ( .DIN(\IDinst/n5290 ), .CLK(clk), 
        .CLRB(n813), .SETB(1'b1), .Q(\IDinst/RegFile[2][19] ) );
  dffascs1 \IDinst/RegFile_reg[3][19]  ( .DIN(\IDinst/n5289 ), .CLK(clk), 
        .CLRB(n813), .SETB(1'b1), .Q(\IDinst/RegFile[3][19] ) );
  dffascs1 \IDinst/RegFile_reg[4][19]  ( .DIN(\IDinst/n5288 ), .CLK(clk), 
        .CLRB(n813), .SETB(1'b1), .Q(\IDinst/RegFile[4][19] ) );
  dffascs1 \IDinst/RegFile_reg[5][19]  ( .DIN(\IDinst/n5287 ), .CLK(clk), 
        .CLRB(n814), .SETB(1'b1), .Q(\IDinst/RegFile[5][19] ) );
  dffascs1 \IDinst/RegFile_reg[6][19]  ( .DIN(\IDinst/n5286 ), .CLK(clk), 
        .CLRB(n814), .SETB(1'b1), .Q(\IDinst/RegFile[6][19] ) );
  dffascs1 \IDinst/RegFile_reg[7][19]  ( .DIN(\IDinst/n5285 ), .CLK(clk), 
        .CLRB(n814), .SETB(1'b1), .Q(\IDinst/RegFile[7][19] ) );
  dffascs1 \IDinst/RegFile_reg[8][19]  ( .DIN(\IDinst/n5284 ), .CLK(clk), 
        .CLRB(n814), .SETB(1'b1), .Q(\IDinst/RegFile[8][19] ) );
  dffascs1 \IDinst/RegFile_reg[9][19]  ( .DIN(\IDinst/n5283 ), .CLK(clk), 
        .CLRB(n814), .SETB(1'b1), .Q(\IDinst/RegFile[9][19] ) );
  dffascs1 \IDinst/RegFile_reg[10][19]  ( .DIN(\IDinst/n5282 ), .CLK(clk), 
        .CLRB(n814), .SETB(1'b1), .Q(\IDinst/RegFile[10][19] ) );
  dffascs1 \IDinst/RegFile_reg[11][19]  ( .DIN(\IDinst/n5281 ), .CLK(clk), 
        .CLRB(n814), .SETB(1'b1), .Q(\IDinst/RegFile[11][19] ) );
  dffascs1 \IDinst/RegFile_reg[12][19]  ( .DIN(\IDinst/n5280 ), .CLK(clk), 
        .CLRB(n814), .SETB(1'b1), .Q(\IDinst/RegFile[12][19] ) );
  dffascs1 \IDinst/RegFile_reg[13][19]  ( .DIN(\IDinst/n5279 ), .CLK(clk), 
        .CLRB(n814), .SETB(1'b1), .Q(\IDinst/RegFile[13][19] ) );
  dffascs1 \IDinst/RegFile_reg[14][19]  ( .DIN(\IDinst/n5278 ), .CLK(clk), 
        .CLRB(n814), .SETB(1'b1), .Q(\IDinst/RegFile[14][19] ) );
  dffascs1 \IDinst/RegFile_reg[15][19]  ( .DIN(\IDinst/n5277 ), .CLK(clk), 
        .CLRB(n815), .SETB(1'b1), .Q(\IDinst/RegFile[15][19] ) );
  dffascs1 \IDinst/RegFile_reg[16][19]  ( .DIN(\IDinst/n5276 ), .CLK(clk), 
        .CLRB(n815), .SETB(1'b1), .Q(\IDinst/RegFile[16][19] ) );
  dffascs1 \IDinst/RegFile_reg[17][19]  ( .DIN(\IDinst/n5275 ), .CLK(clk), 
        .CLRB(n815), .SETB(1'b1), .Q(\IDinst/RegFile[17][19] ) );
  dffascs1 \IDinst/RegFile_reg[18][19]  ( .DIN(\IDinst/n5274 ), .CLK(clk), 
        .CLRB(n815), .SETB(1'b1), .Q(\IDinst/RegFile[18][19] ) );
  dffascs1 \IDinst/RegFile_reg[19][19]  ( .DIN(\IDinst/n5273 ), .CLK(clk), 
        .CLRB(n815), .SETB(1'b1), .Q(\IDinst/RegFile[19][19] ) );
  dffascs1 \IDinst/RegFile_reg[20][19]  ( .DIN(\IDinst/n5272 ), .CLK(clk), 
        .CLRB(n815), .SETB(1'b1), .Q(\IDinst/RegFile[20][19] ) );
  dffascs1 \IDinst/RegFile_reg[21][19]  ( .DIN(\IDinst/n5271 ), .CLK(clk), 
        .CLRB(n815), .SETB(1'b1), .Q(\IDinst/RegFile[21][19] ) );
  dffascs1 \IDinst/RegFile_reg[22][19]  ( .DIN(\IDinst/n5270 ), .CLK(clk), 
        .CLRB(n815), .SETB(1'b1), .Q(\IDinst/RegFile[22][19] ) );
  dffascs1 \IDinst/RegFile_reg[23][19]  ( .DIN(\IDinst/n5269 ), .CLK(clk), 
        .CLRB(n815), .SETB(1'b1), .Q(\IDinst/RegFile[23][19] ) );
  dffascs1 \IDinst/RegFile_reg[24][19]  ( .DIN(\IDinst/n5268 ), .CLK(clk), 
        .CLRB(n815), .SETB(1'b1), .Q(\IDinst/RegFile[24][19] ) );
  dffascs1 \IDinst/RegFile_reg[25][19]  ( .DIN(\IDinst/n5267 ), .CLK(clk), 
        .CLRB(n816), .SETB(1'b1), .Q(\IDinst/RegFile[25][19] ) );
  dffascs1 \IDinst/RegFile_reg[26][19]  ( .DIN(\IDinst/n5266 ), .CLK(clk), 
        .CLRB(n816), .SETB(1'b1), .Q(\IDinst/RegFile[26][19] ) );
  dffascs1 \IDinst/RegFile_reg[27][19]  ( .DIN(\IDinst/n5265 ), .CLK(clk), 
        .CLRB(n816), .SETB(1'b1), .Q(\IDinst/RegFile[27][19] ) );
  dffascs1 \IDinst/RegFile_reg[28][19]  ( .DIN(\IDinst/n5264 ), .CLK(clk), 
        .CLRB(n816), .SETB(1'b1), .Q(\IDinst/RegFile[28][19] ) );
  dffascs1 \IDinst/RegFile_reg[29][19]  ( .DIN(\IDinst/n5263 ), .CLK(clk), 
        .CLRB(n816), .SETB(1'b1), .Q(\IDinst/RegFile[29][19] ) );
  dffascs1 \IDinst/RegFile_reg[30][19]  ( .DIN(\IDinst/n5262 ), .CLK(clk), 
        .CLRB(n816), .SETB(1'b1), .Q(\IDinst/RegFile[30][19] ) );
  dffascs1 \IDinst/RegFile_reg[31][19]  ( .DIN(\IDinst/n5261 ), .CLK(clk), 
        .CLRB(n816), .SETB(1'b1), .Q(\IDinst/RegFile[31][19] ) );
  dffascs1 \IDinst/RegFile_reg[0][20]  ( .DIN(\IDinst/n5260 ), .CLK(clk), 
        .CLRB(n884), .SETB(1'b1), .Q(\IDinst/RegFile[0][20] ) );
  dffascs1 \IDinst/RegFile_reg[1][20]  ( .DIN(\IDinst/n5259 ), .CLK(clk), 
        .CLRB(n884), .SETB(1'b1), .Q(\IDinst/RegFile[1][20] ) );
  dffascs1 \IDinst/RegFile_reg[2][20]  ( .DIN(\IDinst/n5258 ), .CLK(clk), 
        .CLRB(n885), .SETB(1'b1), .Q(\IDinst/RegFile[2][20] ) );
  dffascs1 \IDinst/RegFile_reg[3][20]  ( .DIN(\IDinst/n5257 ), .CLK(clk), 
        .CLRB(n885), .SETB(1'b1), .Q(\IDinst/RegFile[3][20] ) );
  dffascs1 \IDinst/RegFile_reg[4][20]  ( .DIN(\IDinst/n5256 ), .CLK(clk), 
        .CLRB(n885), .SETB(1'b1), .Q(\IDinst/RegFile[4][20] ) );
  dffascs1 \IDinst/RegFile_reg[5][20]  ( .DIN(\IDinst/n5255 ), .CLK(clk), 
        .CLRB(n885), .SETB(1'b1), .Q(\IDinst/RegFile[5][20] ) );
  dffascs1 \IDinst/RegFile_reg[6][20]  ( .DIN(\IDinst/n5254 ), .CLK(clk), 
        .CLRB(n885), .SETB(1'b1), .Q(\IDinst/RegFile[6][20] ) );
  dffascs1 \IDinst/RegFile_reg[7][20]  ( .DIN(\IDinst/n5253 ), .CLK(clk), 
        .CLRB(n885), .SETB(1'b1), .Q(\IDinst/RegFile[7][20] ) );
  dffascs1 \IDinst/RegFile_reg[8][20]  ( .DIN(\IDinst/n5252 ), .CLK(clk), 
        .CLRB(n885), .SETB(1'b1), .Q(\IDinst/RegFile[8][20] ) );
  dffascs1 \IDinst/RegFile_reg[9][20]  ( .DIN(\IDinst/n5251 ), .CLK(clk), 
        .CLRB(n885), .SETB(1'b1), .Q(\IDinst/RegFile[9][20] ) );
  dffascs1 \IDinst/RegFile_reg[10][20]  ( .DIN(\IDinst/n5250 ), .CLK(clk), 
        .CLRB(n885), .SETB(1'b1), .Q(\IDinst/RegFile[10][20] ) );
  dffascs1 \IDinst/RegFile_reg[11][20]  ( .DIN(\IDinst/n5249 ), .CLK(clk), 
        .CLRB(n885), .SETB(1'b1), .Q(\IDinst/RegFile[11][20] ) );
  dffascs1 \IDinst/RegFile_reg[12][20]  ( .DIN(\IDinst/n5248 ), .CLK(clk), 
        .CLRB(n886), .SETB(1'b1), .Q(\IDinst/RegFile[12][20] ) );
  dffascs1 \IDinst/RegFile_reg[13][20]  ( .DIN(\IDinst/n5247 ), .CLK(clk), 
        .CLRB(n886), .SETB(1'b1), .Q(\IDinst/RegFile[13][20] ) );
  dffascs1 \IDinst/RegFile_reg[14][20]  ( .DIN(\IDinst/n5246 ), .CLK(clk), 
        .CLRB(n886), .SETB(1'b1), .Q(\IDinst/RegFile[14][20] ) );
  dffascs1 \IDinst/RegFile_reg[15][20]  ( .DIN(\IDinst/n5245 ), .CLK(clk), 
        .CLRB(n886), .SETB(1'b1), .Q(\IDinst/RegFile[15][20] ) );
  dffascs1 \IDinst/RegFile_reg[16][20]  ( .DIN(\IDinst/n5244 ), .CLK(clk), 
        .CLRB(n886), .SETB(1'b1), .Q(\IDinst/RegFile[16][20] ) );
  dffascs1 \IDinst/RegFile_reg[17][20]  ( .DIN(\IDinst/n5243 ), .CLK(clk), 
        .CLRB(n886), .SETB(1'b1), .Q(\IDinst/RegFile[17][20] ) );
  dffascs1 \IDinst/RegFile_reg[18][20]  ( .DIN(\IDinst/n5242 ), .CLK(clk), 
        .CLRB(n886), .SETB(1'b1), .Q(\IDinst/RegFile[18][20] ) );
  dffascs1 \IDinst/RegFile_reg[19][20]  ( .DIN(\IDinst/n5241 ), .CLK(clk), 
        .CLRB(n886), .SETB(1'b1), .Q(\IDinst/RegFile[19][20] ) );
  dffascs1 \IDinst/RegFile_reg[20][20]  ( .DIN(\IDinst/n5240 ), .CLK(clk), 
        .CLRB(n886), .SETB(1'b1), .Q(\IDinst/RegFile[20][20] ) );
  dffascs1 \IDinst/RegFile_reg[21][20]  ( .DIN(\IDinst/n5239 ), .CLK(clk), 
        .CLRB(n886), .SETB(1'b1), .Q(\IDinst/RegFile[21][20] ) );
  dffascs1 \IDinst/RegFile_reg[22][20]  ( .DIN(\IDinst/n5238 ), .CLK(clk), 
        .CLRB(n887), .SETB(1'b1), .Q(\IDinst/RegFile[22][20] ) );
  dffascs1 \IDinst/RegFile_reg[23][20]  ( .DIN(\IDinst/n5237 ), .CLK(clk), 
        .CLRB(n887), .SETB(1'b1), .Q(\IDinst/RegFile[23][20] ) );
  dffascs1 \IDinst/RegFile_reg[24][20]  ( .DIN(\IDinst/n5236 ), .CLK(clk), 
        .CLRB(n887), .SETB(1'b1), .Q(\IDinst/RegFile[24][20] ) );
  dffascs1 \IDinst/RegFile_reg[25][20]  ( .DIN(\IDinst/n5235 ), .CLK(clk), 
        .CLRB(n887), .SETB(1'b1), .Q(\IDinst/RegFile[25][20] ) );
  dffascs1 \IDinst/RegFile_reg[26][20]  ( .DIN(\IDinst/n5234 ), .CLK(clk), 
        .CLRB(n887), .SETB(1'b1), .Q(\IDinst/RegFile[26][20] ) );
  dffascs1 \IDinst/RegFile_reg[27][20]  ( .DIN(\IDinst/n5233 ), .CLK(clk), 
        .CLRB(n887), .SETB(1'b1), .Q(\IDinst/RegFile[27][20] ) );
  dffascs1 \IDinst/RegFile_reg[28][20]  ( .DIN(\IDinst/n5232 ), .CLK(clk), 
        .CLRB(n887), .SETB(1'b1), .Q(\IDinst/RegFile[28][20] ) );
  dffascs1 \IDinst/RegFile_reg[29][20]  ( .DIN(\IDinst/n5231 ), .CLK(clk), 
        .CLRB(n887), .SETB(1'b1), .Q(\IDinst/RegFile[29][20] ) );
  dffascs1 \IDinst/RegFile_reg[30][20]  ( .DIN(\IDinst/n5230 ), .CLK(clk), 
        .CLRB(n887), .SETB(1'b1), .Q(\IDinst/RegFile[30][20] ) );
  dffascs1 \IDinst/RegFile_reg[31][20]  ( .DIN(\IDinst/n5229 ), .CLK(clk), 
        .CLRB(n887), .SETB(1'b1), .Q(\IDinst/RegFile[31][20] ) );
  dffascs1 \IDinst/RegFile_reg[0][21]  ( .DIN(\IDinst/n5228 ), .CLK(clk), 
        .CLRB(n824), .SETB(1'b1), .Q(\IDinst/RegFile[0][21] ) );
  dffascs1 \IDinst/RegFile_reg[1][21]  ( .DIN(\IDinst/n5227 ), .CLK(clk), 
        .CLRB(n824), .SETB(1'b1), .Q(\IDinst/RegFile[1][21] ) );
  dffascs1 \IDinst/RegFile_reg[2][21]  ( .DIN(\IDinst/n5226 ), .CLK(clk), 
        .CLRB(n825), .SETB(1'b1), .Q(\IDinst/RegFile[2][21] ) );
  dffascs1 \IDinst/RegFile_reg[3][21]  ( .DIN(\IDinst/n5225 ), .CLK(clk), 
        .CLRB(n825), .SETB(1'b1), .Q(\IDinst/RegFile[3][21] ) );
  dffascs1 \IDinst/RegFile_reg[4][21]  ( .DIN(\IDinst/n5224 ), .CLK(clk), 
        .CLRB(n825), .SETB(1'b1), .Q(\IDinst/RegFile[4][21] ) );
  dffascs1 \IDinst/RegFile_reg[5][21]  ( .DIN(\IDinst/n5223 ), .CLK(clk), 
        .CLRB(n825), .SETB(1'b1), .Q(\IDinst/RegFile[5][21] ) );
  dffascs1 \IDinst/RegFile_reg[6][21]  ( .DIN(\IDinst/n5222 ), .CLK(clk), 
        .CLRB(n825), .SETB(1'b1), .Q(\IDinst/RegFile[6][21] ) );
  dffascs1 \IDinst/RegFile_reg[7][21]  ( .DIN(\IDinst/n5221 ), .CLK(clk), 
        .CLRB(n825), .SETB(1'b1), .Q(\IDinst/RegFile[7][21] ) );
  dffascs1 \IDinst/RegFile_reg[8][21]  ( .DIN(\IDinst/n5220 ), .CLK(clk), 
        .CLRB(n825), .SETB(1'b1), .Q(\IDinst/RegFile[8][21] ) );
  dffascs1 \IDinst/RegFile_reg[9][21]  ( .DIN(\IDinst/n5219 ), .CLK(clk), 
        .CLRB(n825), .SETB(1'b1), .Q(\IDinst/RegFile[9][21] ) );
  dffascs1 \IDinst/RegFile_reg[10][21]  ( .DIN(\IDinst/n5218 ), .CLK(clk), 
        .CLRB(n825), .SETB(1'b1), .Q(\IDinst/RegFile[10][21] ) );
  dffascs1 \IDinst/RegFile_reg[11][21]  ( .DIN(\IDinst/n5217 ), .CLK(clk), 
        .CLRB(n825), .SETB(1'b1), .Q(\IDinst/RegFile[11][21] ) );
  dffascs1 \IDinst/RegFile_reg[12][21]  ( .DIN(\IDinst/n5216 ), .CLK(clk), 
        .CLRB(n826), .SETB(1'b1), .Q(\IDinst/RegFile[12][21] ) );
  dffascs1 \IDinst/RegFile_reg[13][21]  ( .DIN(\IDinst/n5215 ), .CLK(clk), 
        .CLRB(n826), .SETB(1'b1), .Q(\IDinst/RegFile[13][21] ) );
  dffascs1 \IDinst/RegFile_reg[14][21]  ( .DIN(\IDinst/n5214 ), .CLK(clk), 
        .CLRB(n826), .SETB(1'b1), .Q(\IDinst/RegFile[14][21] ) );
  dffascs1 \IDinst/RegFile_reg[15][21]  ( .DIN(\IDinst/n5213 ), .CLK(clk), 
        .CLRB(n826), .SETB(1'b1), .Q(\IDinst/RegFile[15][21] ) );
  dffascs1 \IDinst/RegFile_reg[16][21]  ( .DIN(\IDinst/n5212 ), .CLK(clk), 
        .CLRB(n826), .SETB(1'b1), .Q(\IDinst/RegFile[16][21] ) );
  dffascs1 \IDinst/RegFile_reg[17][21]  ( .DIN(\IDinst/n5211 ), .CLK(clk), 
        .CLRB(n826), .SETB(1'b1), .Q(\IDinst/RegFile[17][21] ) );
  dffascs1 \IDinst/RegFile_reg[18][21]  ( .DIN(\IDinst/n5210 ), .CLK(clk), 
        .CLRB(n826), .SETB(1'b1), .Q(\IDinst/RegFile[18][21] ) );
  dffascs1 \IDinst/RegFile_reg[19][21]  ( .DIN(\IDinst/n5209 ), .CLK(clk), 
        .CLRB(n826), .SETB(1'b1), .Q(\IDinst/RegFile[19][21] ) );
  dffascs1 \IDinst/RegFile_reg[20][21]  ( .DIN(\IDinst/n5208 ), .CLK(clk), 
        .CLRB(n826), .SETB(1'b1), .Q(\IDinst/RegFile[20][21] ) );
  dffascs1 \IDinst/RegFile_reg[21][21]  ( .DIN(\IDinst/n5207 ), .CLK(clk), 
        .CLRB(n826), .SETB(1'b1), .Q(\IDinst/RegFile[21][21] ) );
  dffascs1 \IDinst/RegFile_reg[22][21]  ( .DIN(\IDinst/n5206 ), .CLK(clk), 
        .CLRB(n827), .SETB(1'b1), .Q(\IDinst/RegFile[22][21] ) );
  dffascs1 \IDinst/RegFile_reg[23][21]  ( .DIN(\IDinst/n5205 ), .CLK(clk), 
        .CLRB(n827), .SETB(1'b1), .Q(\IDinst/RegFile[23][21] ) );
  dffascs1 \IDinst/RegFile_reg[24][21]  ( .DIN(\IDinst/n5204 ), .CLK(clk), 
        .CLRB(n827), .SETB(1'b1), .Q(\IDinst/RegFile[24][21] ) );
  dffascs1 \IDinst/RegFile_reg[25][21]  ( .DIN(\IDinst/n5203 ), .CLK(clk), 
        .CLRB(n827), .SETB(1'b1), .Q(\IDinst/RegFile[25][21] ) );
  dffascs1 \IDinst/RegFile_reg[26][21]  ( .DIN(\IDinst/n5202 ), .CLK(clk), 
        .CLRB(n827), .SETB(1'b1), .Q(\IDinst/RegFile[26][21] ) );
  dffascs1 \IDinst/RegFile_reg[27][21]  ( .DIN(\IDinst/n5201 ), .CLK(clk), 
        .CLRB(n827), .SETB(1'b1), .Q(\IDinst/RegFile[27][21] ) );
  dffascs1 \IDinst/RegFile_reg[28][21]  ( .DIN(\IDinst/n5200 ), .CLK(clk), 
        .CLRB(n827), .SETB(1'b1), .Q(\IDinst/RegFile[28][21] ) );
  dffascs1 \IDinst/RegFile_reg[29][21]  ( .DIN(\IDinst/n5199 ), .CLK(clk), 
        .CLRB(n827), .SETB(1'b1), .Q(\IDinst/RegFile[29][21] ) );
  dffascs1 \IDinst/RegFile_reg[30][21]  ( .DIN(\IDinst/n5198 ), .CLK(clk), 
        .CLRB(n827), .SETB(1'b1), .Q(\IDinst/RegFile[30][21] ) );
  dffascs1 \IDinst/RegFile_reg[31][21]  ( .DIN(\IDinst/n5197 ), .CLK(clk), 
        .CLRB(n827), .SETB(1'b1), .Q(\IDinst/RegFile[31][21] ) );
  dffascs1 \IDinst/RegFile_reg[0][22]  ( .DIN(\IDinst/n5196 ), .CLK(clk), 
        .CLRB(n880), .SETB(1'b1), .Q(\IDinst/RegFile[0][22] ) );
  dffascs1 \IDinst/RegFile_reg[1][22]  ( .DIN(\IDinst/n5195 ), .CLK(clk), 
        .CLRB(n880), .SETB(1'b1), .Q(\IDinst/RegFile[1][22] ) );
  dffascs1 \IDinst/RegFile_reg[2][22]  ( .DIN(\IDinst/n5194 ), .CLK(clk), 
        .CLRB(n880), .SETB(1'b1), .Q(\IDinst/RegFile[2][22] ) );
  dffascs1 \IDinst/RegFile_reg[3][22]  ( .DIN(\IDinst/n5193 ), .CLK(clk), 
        .CLRB(n881), .SETB(1'b1), .Q(\IDinst/RegFile[3][22] ) );
  dffascs1 \IDinst/RegFile_reg[4][22]  ( .DIN(\IDinst/n5192 ), .CLK(clk), 
        .CLRB(n881), .SETB(1'b1), .Q(\IDinst/RegFile[4][22] ) );
  dffascs1 \IDinst/RegFile_reg[5][22]  ( .DIN(\IDinst/n5191 ), .CLK(clk), 
        .CLRB(n881), .SETB(1'b1), .Q(\IDinst/RegFile[5][22] ) );
  dffascs1 \IDinst/RegFile_reg[6][22]  ( .DIN(\IDinst/n5190 ), .CLK(clk), 
        .CLRB(n881), .SETB(1'b1), .Q(\IDinst/RegFile[6][22] ) );
  dffascs1 \IDinst/RegFile_reg[7][22]  ( .DIN(\IDinst/n5189 ), .CLK(clk), 
        .CLRB(n881), .SETB(1'b1), .Q(\IDinst/RegFile[7][22] ) );
  dffascs1 \IDinst/RegFile_reg[8][22]  ( .DIN(\IDinst/n5188 ), .CLK(clk), 
        .CLRB(n881), .SETB(1'b1), .Q(\IDinst/RegFile[8][22] ) );
  dffascs1 \IDinst/RegFile_reg[9][22]  ( .DIN(\IDinst/n5187 ), .CLK(clk), 
        .CLRB(n881), .SETB(1'b1), .Q(\IDinst/RegFile[9][22] ) );
  dffascs1 \IDinst/RegFile_reg[10][22]  ( .DIN(\IDinst/n5186 ), .CLK(clk), 
        .CLRB(n881), .SETB(1'b1), .Q(\IDinst/RegFile[10][22] ) );
  dffascs1 \IDinst/RegFile_reg[11][22]  ( .DIN(\IDinst/n5185 ), .CLK(clk), 
        .CLRB(n881), .SETB(1'b1), .Q(\IDinst/RegFile[11][22] ) );
  dffascs1 \IDinst/RegFile_reg[12][22]  ( .DIN(\IDinst/n5184 ), .CLK(clk), 
        .CLRB(n881), .SETB(1'b1), .Q(\IDinst/RegFile[12][22] ) );
  dffascs1 \IDinst/RegFile_reg[13][22]  ( .DIN(\IDinst/n5183 ), .CLK(clk), 
        .CLRB(n882), .SETB(1'b1), .Q(\IDinst/RegFile[13][22] ) );
  dffascs1 \IDinst/RegFile_reg[14][22]  ( .DIN(\IDinst/n5182 ), .CLK(clk), 
        .CLRB(n882), .SETB(1'b1), .Q(\IDinst/RegFile[14][22] ) );
  dffascs1 \IDinst/RegFile_reg[15][22]  ( .DIN(\IDinst/n5181 ), .CLK(clk), 
        .CLRB(n882), .SETB(1'b1), .Q(\IDinst/RegFile[15][22] ) );
  dffascs1 \IDinst/RegFile_reg[16][22]  ( .DIN(\IDinst/n5180 ), .CLK(clk), 
        .CLRB(n882), .SETB(1'b1), .Q(\IDinst/RegFile[16][22] ) );
  dffascs1 \IDinst/RegFile_reg[17][22]  ( .DIN(\IDinst/n5179 ), .CLK(clk), 
        .CLRB(n882), .SETB(1'b1), .Q(\IDinst/RegFile[17][22] ) );
  dffascs1 \IDinst/RegFile_reg[18][22]  ( .DIN(\IDinst/n5178 ), .CLK(clk), 
        .CLRB(n882), .SETB(1'b1), .Q(\IDinst/RegFile[18][22] ) );
  dffascs1 \IDinst/RegFile_reg[19][22]  ( .DIN(\IDinst/n5177 ), .CLK(clk), 
        .CLRB(n882), .SETB(1'b1), .Q(\IDinst/RegFile[19][22] ) );
  dffascs1 \IDinst/RegFile_reg[20][22]  ( .DIN(\IDinst/n5176 ), .CLK(clk), 
        .CLRB(n882), .SETB(1'b1), .Q(\IDinst/RegFile[20][22] ) );
  dffascs1 \IDinst/RegFile_reg[21][22]  ( .DIN(\IDinst/n5175 ), .CLK(clk), 
        .CLRB(n882), .SETB(1'b1), .Q(\IDinst/RegFile[21][22] ) );
  dffascs1 \IDinst/RegFile_reg[22][22]  ( .DIN(\IDinst/n5174 ), .CLK(clk), 
        .CLRB(n882), .SETB(1'b1), .Q(\IDinst/RegFile[22][22] ) );
  dffascs1 \IDinst/RegFile_reg[23][22]  ( .DIN(\IDinst/n5173 ), .CLK(clk), 
        .CLRB(n883), .SETB(1'b1), .Q(\IDinst/RegFile[23][22] ) );
  dffascs1 \IDinst/RegFile_reg[24][22]  ( .DIN(\IDinst/n5172 ), .CLK(clk), 
        .CLRB(n883), .SETB(1'b1), .Q(\IDinst/RegFile[24][22] ) );
  dffascs1 \IDinst/RegFile_reg[25][22]  ( .DIN(\IDinst/n5171 ), .CLK(clk), 
        .CLRB(n883), .SETB(1'b1), .Q(\IDinst/RegFile[25][22] ) );
  dffascs1 \IDinst/RegFile_reg[26][22]  ( .DIN(\IDinst/n5170 ), .CLK(clk), 
        .CLRB(n883), .SETB(1'b1), .Q(\IDinst/RegFile[26][22] ) );
  dffascs1 \IDinst/RegFile_reg[27][22]  ( .DIN(\IDinst/n5169 ), .CLK(clk), 
        .CLRB(n883), .SETB(1'b1), .Q(\IDinst/RegFile[27][22] ) );
  dffascs1 \IDinst/RegFile_reg[28][22]  ( .DIN(\IDinst/n5168 ), .CLK(clk), 
        .CLRB(n883), .SETB(1'b1), .Q(\IDinst/RegFile[28][22] ) );
  dffascs1 \IDinst/RegFile_reg[29][22]  ( .DIN(\IDinst/n5167 ), .CLK(clk), 
        .CLRB(n883), .SETB(1'b1), .Q(\IDinst/RegFile[29][22] ) );
  dffascs1 \IDinst/RegFile_reg[30][22]  ( .DIN(\IDinst/n5166 ), .CLK(clk), 
        .CLRB(n883), .SETB(1'b1), .Q(\IDinst/RegFile[30][22] ) );
  dffascs1 \IDinst/RegFile_reg[31][22]  ( .DIN(\IDinst/n5165 ), .CLK(clk), 
        .CLRB(n883), .SETB(1'b1), .Q(\IDinst/RegFile[31][22] ) );
  dffascs1 \IDinst/RegFile_reg[0][23]  ( .DIN(\IDinst/n5164 ), .CLK(clk), 
        .CLRB(n888), .SETB(1'b1), .Q(\IDinst/RegFile[0][23] ) );
  dffascs1 \IDinst/RegFile_reg[1][23]  ( .DIN(\IDinst/n5163 ), .CLK(clk), 
        .CLRB(n888), .SETB(1'b1), .Q(\IDinst/RegFile[1][23] ) );
  dffascs1 \IDinst/RegFile_reg[2][23]  ( .DIN(\IDinst/n5162 ), .CLK(clk), 
        .CLRB(n888), .SETB(1'b1), .Q(\IDinst/RegFile[2][23] ) );
  dffascs1 \IDinst/RegFile_reg[3][23]  ( .DIN(\IDinst/n5161 ), .CLK(clk), 
        .CLRB(n888), .SETB(1'b1), .Q(\IDinst/RegFile[3][23] ) );
  dffascs1 \IDinst/RegFile_reg[4][23]  ( .DIN(\IDinst/n5160 ), .CLK(clk), 
        .CLRB(n889), .SETB(1'b1), .Q(\IDinst/RegFile[4][23] ) );
  dffascs1 \IDinst/RegFile_reg[5][23]  ( .DIN(\IDinst/n5159 ), .CLK(clk), 
        .CLRB(n889), .SETB(1'b1), .Q(\IDinst/RegFile[5][23] ) );
  dffascs1 \IDinst/RegFile_reg[6][23]  ( .DIN(\IDinst/n5158 ), .CLK(clk), 
        .CLRB(n889), .SETB(1'b1), .Q(\IDinst/RegFile[6][23] ) );
  dffascs1 \IDinst/RegFile_reg[7][23]  ( .DIN(\IDinst/n5157 ), .CLK(clk), 
        .CLRB(n889), .SETB(1'b1), .Q(\IDinst/RegFile[7][23] ) );
  dffascs1 \IDinst/RegFile_reg[8][23]  ( .DIN(\IDinst/n5156 ), .CLK(clk), 
        .CLRB(n889), .SETB(1'b1), .Q(\IDinst/RegFile[8][23] ) );
  dffascs1 \IDinst/RegFile_reg[9][23]  ( .DIN(\IDinst/n5155 ), .CLK(clk), 
        .CLRB(n889), .SETB(1'b1), .Q(\IDinst/RegFile[9][23] ) );
  dffascs1 \IDinst/RegFile_reg[10][23]  ( .DIN(\IDinst/n5154 ), .CLK(clk), 
        .CLRB(n889), .SETB(1'b1), .Q(\IDinst/RegFile[10][23] ) );
  dffascs1 \IDinst/RegFile_reg[11][23]  ( .DIN(\IDinst/n5153 ), .CLK(clk), 
        .CLRB(n889), .SETB(1'b1), .Q(\IDinst/RegFile[11][23] ) );
  dffascs1 \IDinst/RegFile_reg[12][23]  ( .DIN(\IDinst/n5152 ), .CLK(clk), 
        .CLRB(n889), .SETB(1'b1), .Q(\IDinst/RegFile[12][23] ) );
  dffascs1 \IDinst/RegFile_reg[13][23]  ( .DIN(\IDinst/n5151 ), .CLK(clk), 
        .CLRB(n889), .SETB(1'b1), .Q(\IDinst/RegFile[13][23] ) );
  dffascs1 \IDinst/RegFile_reg[14][23]  ( .DIN(\IDinst/n5150 ), .CLK(clk), 
        .CLRB(n890), .SETB(1'b1), .Q(\IDinst/RegFile[14][23] ) );
  dffascs1 \IDinst/RegFile_reg[15][23]  ( .DIN(\IDinst/n5149 ), .CLK(clk), 
        .CLRB(n890), .SETB(1'b1), .Q(\IDinst/RegFile[15][23] ) );
  dffascs1 \IDinst/RegFile_reg[16][23]  ( .DIN(\IDinst/n5148 ), .CLK(clk), 
        .CLRB(n890), .SETB(1'b1), .Q(\IDinst/RegFile[16][23] ) );
  dffascs1 \IDinst/RegFile_reg[17][23]  ( .DIN(\IDinst/n5147 ), .CLK(clk), 
        .CLRB(n890), .SETB(1'b1), .Q(\IDinst/RegFile[17][23] ) );
  dffascs1 \IDinst/RegFile_reg[18][23]  ( .DIN(\IDinst/n5146 ), .CLK(clk), 
        .CLRB(n890), .SETB(1'b1), .Q(\IDinst/RegFile[18][23] ) );
  dffascs1 \IDinst/RegFile_reg[19][23]  ( .DIN(\IDinst/n5145 ), .CLK(clk), 
        .CLRB(n890), .SETB(1'b1), .Q(\IDinst/RegFile[19][23] ) );
  dffascs1 \IDinst/RegFile_reg[20][23]  ( .DIN(\IDinst/n5144 ), .CLK(clk), 
        .CLRB(n890), .SETB(1'b1), .Q(\IDinst/RegFile[20][23] ) );
  dffascs1 \IDinst/RegFile_reg[21][23]  ( .DIN(\IDinst/n5143 ), .CLK(clk), 
        .CLRB(n890), .SETB(1'b1), .Q(\IDinst/RegFile[21][23] ) );
  dffascs1 \IDinst/RegFile_reg[22][23]  ( .DIN(\IDinst/n5142 ), .CLK(clk), 
        .CLRB(n890), .SETB(1'b1), .Q(\IDinst/RegFile[22][23] ) );
  dffascs1 \IDinst/RegFile_reg[23][23]  ( .DIN(\IDinst/n5141 ), .CLK(clk), 
        .CLRB(n890), .SETB(1'b1), .Q(\IDinst/RegFile[23][23] ) );
  dffascs1 \IDinst/RegFile_reg[24][23]  ( .DIN(\IDinst/n5140 ), .CLK(clk), 
        .CLRB(n891), .SETB(1'b1), .Q(\IDinst/RegFile[24][23] ) );
  dffascs1 \IDinst/RegFile_reg[25][23]  ( .DIN(\IDinst/n5139 ), .CLK(clk), 
        .CLRB(n891), .SETB(1'b1), .Q(\IDinst/RegFile[25][23] ) );
  dffascs1 \IDinst/RegFile_reg[26][23]  ( .DIN(\IDinst/n5138 ), .CLK(clk), 
        .CLRB(n891), .SETB(1'b1), .Q(\IDinst/RegFile[26][23] ) );
  dffascs1 \IDinst/RegFile_reg[27][23]  ( .DIN(\IDinst/n5137 ), .CLK(clk), 
        .CLRB(n891), .SETB(1'b1), .Q(\IDinst/RegFile[27][23] ) );
  dffascs1 \IDinst/RegFile_reg[28][23]  ( .DIN(\IDinst/n5136 ), .CLK(clk), 
        .CLRB(n891), .SETB(1'b1), .Q(\IDinst/RegFile[28][23] ) );
  dffascs1 \IDinst/RegFile_reg[29][23]  ( .DIN(\IDinst/n5135 ), .CLK(clk), 
        .CLRB(n891), .SETB(1'b1), .Q(\IDinst/RegFile[29][23] ) );
  dffascs1 \IDinst/RegFile_reg[30][23]  ( .DIN(\IDinst/n5134 ), .CLK(clk), 
        .CLRB(n891), .SETB(1'b1), .Q(\IDinst/RegFile[30][23] ) );
  dffascs1 \IDinst/RegFile_reg[31][23]  ( .DIN(\IDinst/n5133 ), .CLK(clk), 
        .CLRB(n891), .SETB(1'b1), .Q(\IDinst/RegFile[31][23] ) );
  dffascs1 \IDinst/RegFile_reg[0][24]  ( .DIN(\IDinst/n5132 ), .CLK(clk), 
        .CLRB(n903), .SETB(1'b1), .Q(\IDinst/RegFile[0][24] ) );
  dffascs1 \IDinst/RegFile_reg[1][24]  ( .DIN(\IDinst/n5131 ), .CLK(clk), 
        .CLRB(n903), .SETB(1'b1), .Q(\IDinst/RegFile[1][24] ) );
  dffascs1 \IDinst/RegFile_reg[2][24]  ( .DIN(\IDinst/n5130 ), .CLK(clk), 
        .CLRB(n903), .SETB(1'b1), .Q(\IDinst/RegFile[2][24] ) );
  dffascs1 \IDinst/RegFile_reg[3][24]  ( .DIN(\IDinst/n5129 ), .CLK(clk), 
        .CLRB(n903), .SETB(1'b1), .Q(\IDinst/RegFile[3][24] ) );
  dffascs1 \IDinst/RegFile_reg[4][24]  ( .DIN(\IDinst/n5128 ), .CLK(clk), 
        .CLRB(n903), .SETB(1'b1), .Q(\IDinst/RegFile[4][24] ) );
  dffascs1 \IDinst/RegFile_reg[5][24]  ( .DIN(\IDinst/n5127 ), .CLK(clk), 
        .CLRB(n903), .SETB(1'b1), .Q(\IDinst/RegFile[5][24] ) );
  dffascs1 \IDinst/RegFile_reg[6][24]  ( .DIN(\IDinst/n5126 ), .CLK(clk), 
        .CLRB(n903), .SETB(1'b1), .Q(\IDinst/RegFile[6][24] ) );
  dffascs1 \IDinst/RegFile_reg[7][24]  ( .DIN(\IDinst/n5125 ), .CLK(clk), 
        .CLRB(n903), .SETB(1'b1), .Q(\IDinst/RegFile[7][24] ) );
  dffascs1 \IDinst/RegFile_reg[8][24]  ( .DIN(\IDinst/n5124 ), .CLK(clk), 
        .CLRB(n903), .SETB(1'b1), .Q(\IDinst/RegFile[8][24] ) );
  dffascs1 \IDinst/RegFile_reg[9][24]  ( .DIN(\IDinst/n5123 ), .CLK(clk), 
        .CLRB(n903), .SETB(1'b1), .Q(\IDinst/RegFile[9][24] ) );
  dffascs1 \IDinst/RegFile_reg[10][24]  ( .DIN(\IDinst/n5122 ), .CLK(clk), 
        .CLRB(n904), .SETB(1'b1), .Q(\IDinst/RegFile[10][24] ) );
  dffascs1 \IDinst/RegFile_reg[11][24]  ( .DIN(\IDinst/n5121 ), .CLK(clk), 
        .CLRB(n904), .SETB(1'b1), .Q(\IDinst/RegFile[11][24] ) );
  dffascs1 \IDinst/RegFile_reg[12][24]  ( .DIN(\IDinst/n5120 ), .CLK(clk), 
        .CLRB(n904), .SETB(1'b1), .Q(\IDinst/RegFile[12][24] ) );
  dffascs1 \IDinst/RegFile_reg[13][24]  ( .DIN(\IDinst/n5119 ), .CLK(clk), 
        .CLRB(n904), .SETB(1'b1), .Q(\IDinst/RegFile[13][24] ) );
  dffascs1 \IDinst/RegFile_reg[14][24]  ( .DIN(\IDinst/n5118 ), .CLK(clk), 
        .CLRB(n904), .SETB(1'b1), .Q(\IDinst/RegFile[14][24] ) );
  dffascs1 \IDinst/RegFile_reg[15][24]  ( .DIN(\IDinst/n5117 ), .CLK(clk), 
        .CLRB(n904), .SETB(1'b1), .Q(\IDinst/RegFile[15][24] ) );
  dffascs1 \IDinst/RegFile_reg[16][24]  ( .DIN(\IDinst/n5116 ), .CLK(clk), 
        .CLRB(n904), .SETB(1'b1), .Q(\IDinst/RegFile[16][24] ) );
  dffascs1 \IDinst/RegFile_reg[17][24]  ( .DIN(\IDinst/n5115 ), .CLK(clk), 
        .CLRB(n904), .SETB(1'b1), .Q(\IDinst/RegFile[17][24] ) );
  dffascs1 \IDinst/RegFile_reg[18][24]  ( .DIN(\IDinst/n5114 ), .CLK(clk), 
        .CLRB(n904), .SETB(1'b1), .Q(\IDinst/RegFile[18][24] ) );
  dffascs1 \IDinst/RegFile_reg[19][24]  ( .DIN(\IDinst/n5113 ), .CLK(clk), 
        .CLRB(n904), .SETB(1'b1), .Q(\IDinst/RegFile[19][24] ) );
  dffascs1 \IDinst/RegFile_reg[20][24]  ( .DIN(\IDinst/n5112 ), .CLK(clk), 
        .CLRB(n905), .SETB(1'b1), .Q(\IDinst/RegFile[20][24] ) );
  dffascs1 \IDinst/RegFile_reg[21][24]  ( .DIN(\IDinst/n5111 ), .CLK(clk), 
        .CLRB(n905), .SETB(1'b1), .Q(\IDinst/RegFile[21][24] ) );
  dffascs1 \IDinst/RegFile_reg[22][24]  ( .DIN(\IDinst/n5110 ), .CLK(clk), 
        .CLRB(n905), .SETB(1'b1), .Q(\IDinst/RegFile[22][24] ) );
  dffascs1 \IDinst/RegFile_reg[23][24]  ( .DIN(\IDinst/n5109 ), .CLK(clk), 
        .CLRB(n905), .SETB(1'b1), .Q(\IDinst/RegFile[23][24] ) );
  dffascs1 \IDinst/RegFile_reg[24][24]  ( .DIN(\IDinst/n5108 ), .CLK(clk), 
        .CLRB(n905), .SETB(1'b1), .Q(\IDinst/RegFile[24][24] ) );
  dffascs1 \IDinst/RegFile_reg[25][24]  ( .DIN(\IDinst/n5107 ), .CLK(clk), 
        .CLRB(n905), .SETB(1'b1), .Q(\IDinst/RegFile[25][24] ) );
  dffascs1 \IDinst/RegFile_reg[26][24]  ( .DIN(\IDinst/n5106 ), .CLK(clk), 
        .CLRB(n905), .SETB(1'b1), .Q(\IDinst/RegFile[26][24] ) );
  dffascs1 \IDinst/RegFile_reg[27][24]  ( .DIN(\IDinst/n5105 ), .CLK(clk), 
        .CLRB(n905), .SETB(1'b1), .Q(\IDinst/RegFile[27][24] ) );
  dffascs1 \IDinst/RegFile_reg[28][24]  ( .DIN(\IDinst/n5104 ), .CLK(clk), 
        .CLRB(n905), .SETB(1'b1), .Q(\IDinst/RegFile[28][24] ) );
  dffascs1 \IDinst/RegFile_reg[29][24]  ( .DIN(\IDinst/n5103 ), .CLK(clk), 
        .CLRB(n905), .SETB(1'b1), .Q(\IDinst/RegFile[29][24] ) );
  dffascs1 \IDinst/RegFile_reg[30][24]  ( .DIN(\IDinst/n5102 ), .CLK(clk), 
        .CLRB(n906), .SETB(1'b1), .Q(\IDinst/RegFile[30][24] ) );
  dffascs1 \IDinst/RegFile_reg[31][24]  ( .DIN(\IDinst/n5101 ), .CLK(clk), 
        .CLRB(n906), .SETB(1'b1), .Q(\IDinst/RegFile[31][24] ) );
  dffascs1 \IDinst/RegFile_reg[0][25]  ( .DIN(\IDinst/n5100 ), .CLK(clk), 
        .CLRB(n899), .SETB(1'b1), .Q(\IDinst/RegFile[0][25] ) );
  dffascs1 \IDinst/RegFile_reg[1][25]  ( .DIN(\IDinst/n5099 ), .CLK(clk), 
        .CLRB(n899), .SETB(1'b1), .Q(\IDinst/RegFile[1][25] ) );
  dffascs1 \IDinst/RegFile_reg[2][25]  ( .DIN(\IDinst/n5098 ), .CLK(clk), 
        .CLRB(n899), .SETB(1'b1), .Q(\IDinst/RegFile[2][25] ) );
  dffascs1 \IDinst/RegFile_reg[3][25]  ( .DIN(\IDinst/n5097 ), .CLK(clk), 
        .CLRB(n899), .SETB(1'b1), .Q(\IDinst/RegFile[3][25] ) );
  dffascs1 \IDinst/RegFile_reg[4][25]  ( .DIN(\IDinst/n5096 ), .CLK(clk), 
        .CLRB(n899), .SETB(1'b1), .Q(\IDinst/RegFile[4][25] ) );
  dffascs1 \IDinst/RegFile_reg[5][25]  ( .DIN(\IDinst/n5095 ), .CLK(clk), 
        .CLRB(n900), .SETB(1'b1), .Q(\IDinst/RegFile[5][25] ) );
  dffascs1 \IDinst/RegFile_reg[6][25]  ( .DIN(\IDinst/n5094 ), .CLK(clk), 
        .CLRB(n900), .SETB(1'b1), .Q(\IDinst/RegFile[6][25] ) );
  dffascs1 \IDinst/RegFile_reg[7][25]  ( .DIN(\IDinst/n5093 ), .CLK(clk), 
        .CLRB(n900), .SETB(1'b1), .Q(\IDinst/RegFile[7][25] ) );
  dffascs1 \IDinst/RegFile_reg[8][25]  ( .DIN(\IDinst/n5092 ), .CLK(clk), 
        .CLRB(n900), .SETB(1'b1), .Q(\IDinst/RegFile[8][25] ) );
  dffascs1 \IDinst/RegFile_reg[9][25]  ( .DIN(\IDinst/n5091 ), .CLK(clk), 
        .CLRB(n900), .SETB(1'b1), .Q(\IDinst/RegFile[9][25] ) );
  dffascs1 \IDinst/RegFile_reg[10][25]  ( .DIN(\IDinst/n5090 ), .CLK(clk), 
        .CLRB(n900), .SETB(1'b1), .Q(\IDinst/RegFile[10][25] ) );
  dffascs1 \IDinst/RegFile_reg[11][25]  ( .DIN(\IDinst/n5089 ), .CLK(clk), 
        .CLRB(n900), .SETB(1'b1), .Q(\IDinst/RegFile[11][25] ) );
  dffascs1 \IDinst/RegFile_reg[12][25]  ( .DIN(\IDinst/n5088 ), .CLK(clk), 
        .CLRB(n900), .SETB(1'b1), .Q(\IDinst/RegFile[12][25] ) );
  dffascs1 \IDinst/RegFile_reg[13][25]  ( .DIN(\IDinst/n5087 ), .CLK(clk), 
        .CLRB(n900), .SETB(1'b1), .Q(\IDinst/RegFile[13][25] ) );
  dffascs1 \IDinst/RegFile_reg[14][25]  ( .DIN(\IDinst/n5086 ), .CLK(clk), 
        .CLRB(n900), .SETB(1'b1), .Q(\IDinst/RegFile[14][25] ) );
  dffascs1 \IDinst/RegFile_reg[15][25]  ( .DIN(\IDinst/n5085 ), .CLK(clk), 
        .CLRB(n901), .SETB(1'b1), .Q(\IDinst/RegFile[15][25] ) );
  dffascs1 \IDinst/RegFile_reg[16][25]  ( .DIN(\IDinst/n5084 ), .CLK(clk), 
        .CLRB(n901), .SETB(1'b1), .Q(\IDinst/RegFile[16][25] ) );
  dffascs1 \IDinst/RegFile_reg[17][25]  ( .DIN(\IDinst/n5083 ), .CLK(clk), 
        .CLRB(n901), .SETB(1'b1), .Q(\IDinst/RegFile[17][25] ) );
  dffascs1 \IDinst/RegFile_reg[18][25]  ( .DIN(\IDinst/n5082 ), .CLK(clk), 
        .CLRB(n901), .SETB(1'b1), .Q(\IDinst/RegFile[18][25] ) );
  dffascs1 \IDinst/RegFile_reg[19][25]  ( .DIN(\IDinst/n5081 ), .CLK(clk), 
        .CLRB(n901), .SETB(1'b1), .Q(\IDinst/RegFile[19][25] ) );
  dffascs1 \IDinst/RegFile_reg[20][25]  ( .DIN(\IDinst/n5080 ), .CLK(clk), 
        .CLRB(n901), .SETB(1'b1), .Q(\IDinst/RegFile[20][25] ) );
  dffascs1 \IDinst/RegFile_reg[21][25]  ( .DIN(\IDinst/n5079 ), .CLK(clk), 
        .CLRB(n901), .SETB(1'b1), .Q(\IDinst/RegFile[21][25] ) );
  dffascs1 \IDinst/RegFile_reg[22][25]  ( .DIN(\IDinst/n5078 ), .CLK(clk), 
        .CLRB(n901), .SETB(1'b1), .Q(\IDinst/RegFile[22][25] ) );
  dffascs1 \IDinst/RegFile_reg[23][25]  ( .DIN(\IDinst/n5077 ), .CLK(clk), 
        .CLRB(n901), .SETB(1'b1), .Q(\IDinst/RegFile[23][25] ) );
  dffascs1 \IDinst/RegFile_reg[24][25]  ( .DIN(\IDinst/n5076 ), .CLK(clk), 
        .CLRB(n901), .SETB(1'b1), .Q(\IDinst/RegFile[24][25] ) );
  dffascs1 \IDinst/RegFile_reg[25][25]  ( .DIN(\IDinst/n5075 ), .CLK(clk), 
        .CLRB(n902), .SETB(1'b1), .Q(\IDinst/RegFile[25][25] ) );
  dffascs1 \IDinst/RegFile_reg[26][25]  ( .DIN(\IDinst/n5074 ), .CLK(clk), 
        .CLRB(n902), .SETB(1'b1), .Q(\IDinst/RegFile[26][25] ) );
  dffascs1 \IDinst/RegFile_reg[27][25]  ( .DIN(\IDinst/n5073 ), .CLK(clk), 
        .CLRB(n902), .SETB(1'b1), .Q(\IDinst/RegFile[27][25] ) );
  dffascs1 \IDinst/RegFile_reg[28][25]  ( .DIN(\IDinst/n5072 ), .CLK(clk), 
        .CLRB(n902), .SETB(1'b1), .Q(\IDinst/RegFile[28][25] ) );
  dffascs1 \IDinst/RegFile_reg[29][25]  ( .DIN(\IDinst/n5071 ), .CLK(clk), 
        .CLRB(n902), .SETB(1'b1), .Q(\IDinst/RegFile[29][25] ) );
  dffascs1 \IDinst/RegFile_reg[30][25]  ( .DIN(\IDinst/n5070 ), .CLK(clk), 
        .CLRB(n902), .SETB(1'b1), .Q(\IDinst/RegFile[30][25] ) );
  dffascs1 \IDinst/RegFile_reg[31][25]  ( .DIN(\IDinst/n5069 ), .CLK(clk), 
        .CLRB(n902), .SETB(1'b1), .Q(\IDinst/RegFile[31][25] ) );
  dffascs1 \IDinst/RegFile_reg[0][26]  ( .DIN(\IDinst/n5068 ), .CLK(clk), 
        .CLRB(n910), .SETB(1'b1), .Q(\IDinst/RegFile[0][26] ) );
  dffascs1 \IDinst/RegFile_reg[1][26]  ( .DIN(\IDinst/n5067 ), .CLK(clk), 
        .CLRB(n910), .SETB(1'b1), .Q(\IDinst/RegFile[1][26] ) );
  dffascs1 \IDinst/RegFile_reg[2][26]  ( .DIN(\IDinst/n5066 ), .CLK(clk), 
        .CLRB(n910), .SETB(1'b1), .Q(\IDinst/RegFile[2][26] ) );
  dffascs1 \IDinst/RegFile_reg[3][26]  ( .DIN(\IDinst/n5065 ), .CLK(clk), 
        .CLRB(n910), .SETB(1'b1), .Q(\IDinst/RegFile[3][26] ) );
  dffascs1 \IDinst/RegFile_reg[4][26]  ( .DIN(\IDinst/n5064 ), .CLK(clk), 
        .CLRB(n910), .SETB(1'b1), .Q(\IDinst/RegFile[4][26] ) );
  dffascs1 \IDinst/RegFile_reg[5][26]  ( .DIN(\IDinst/n5063 ), .CLK(clk), 
        .CLRB(n910), .SETB(1'b1), .Q(\IDinst/RegFile[5][26] ) );
  dffascs1 \IDinst/RegFile_reg[6][26]  ( .DIN(\IDinst/n5062 ), .CLK(clk), 
        .CLRB(n910), .SETB(1'b1), .Q(\IDinst/RegFile[6][26] ) );
  dffascs1 \IDinst/RegFile_reg[7][26]  ( .DIN(\IDinst/n5061 ), .CLK(clk), 
        .CLRB(n911), .SETB(1'b1), .Q(\IDinst/RegFile[7][26] ) );
  dffascs1 \IDinst/RegFile_reg[8][26]  ( .DIN(\IDinst/n5060 ), .CLK(clk), 
        .CLRB(n911), .SETB(1'b1), .Q(\IDinst/RegFile[8][26] ) );
  dffascs1 \IDinst/RegFile_reg[9][26]  ( .DIN(\IDinst/n5059 ), .CLK(clk), 
        .CLRB(n911), .SETB(1'b1), .Q(\IDinst/RegFile[9][26] ) );
  dffascs1 \IDinst/RegFile_reg[10][26]  ( .DIN(\IDinst/n5058 ), .CLK(clk), 
        .CLRB(n911), .SETB(1'b1), .Q(\IDinst/RegFile[10][26] ) );
  dffascs1 \IDinst/RegFile_reg[11][26]  ( .DIN(\IDinst/n5057 ), .CLK(clk), 
        .CLRB(n911), .SETB(1'b1), .Q(\IDinst/RegFile[11][26] ) );
  dffascs1 \IDinst/RegFile_reg[12][26]  ( .DIN(\IDinst/n5056 ), .CLK(clk), 
        .CLRB(n911), .SETB(1'b1), .Q(\IDinst/RegFile[12][26] ) );
  dffascs1 \IDinst/RegFile_reg[13][26]  ( .DIN(\IDinst/n5055 ), .CLK(clk), 
        .CLRB(n911), .SETB(1'b1), .Q(\IDinst/RegFile[13][26] ) );
  dffascs1 \IDinst/RegFile_reg[14][26]  ( .DIN(\IDinst/n5054 ), .CLK(clk), 
        .CLRB(n911), .SETB(1'b1), .Q(\IDinst/RegFile[14][26] ) );
  dffascs1 \IDinst/RegFile_reg[15][26]  ( .DIN(\IDinst/n5053 ), .CLK(clk), 
        .CLRB(n911), .SETB(1'b1), .Q(\IDinst/RegFile[15][26] ) );
  dffascs1 \IDinst/RegFile_reg[16][26]  ( .DIN(\IDinst/n5052 ), .CLK(clk), 
        .CLRB(n911), .SETB(1'b1), .Q(\IDinst/RegFile[16][26] ) );
  dffascs1 \IDinst/RegFile_reg[17][26]  ( .DIN(\IDinst/n5051 ), .CLK(clk), 
        .CLRB(n912), .SETB(1'b1), .Q(\IDinst/RegFile[17][26] ) );
  dffascs1 \IDinst/RegFile_reg[18][26]  ( .DIN(\IDinst/n5050 ), .CLK(clk), 
        .CLRB(n912), .SETB(1'b1), .Q(\IDinst/RegFile[18][26] ) );
  dffascs1 \IDinst/RegFile_reg[19][26]  ( .DIN(\IDinst/n5049 ), .CLK(clk), 
        .CLRB(n912), .SETB(1'b1), .Q(\IDinst/RegFile[19][26] ) );
  dffascs1 \IDinst/RegFile_reg[20][26]  ( .DIN(\IDinst/n5048 ), .CLK(clk), 
        .CLRB(n912), .SETB(1'b1), .Q(\IDinst/RegFile[20][26] ) );
  dffascs1 \IDinst/RegFile_reg[21][26]  ( .DIN(\IDinst/n5047 ), .CLK(clk), 
        .CLRB(n912), .SETB(1'b1), .Q(\IDinst/RegFile[21][26] ) );
  dffascs1 \IDinst/RegFile_reg[22][26]  ( .DIN(\IDinst/n5046 ), .CLK(clk), 
        .CLRB(n912), .SETB(1'b1), .Q(\IDinst/RegFile[22][26] ) );
  dffascs1 \IDinst/RegFile_reg[23][26]  ( .DIN(\IDinst/n5045 ), .CLK(clk), 
        .CLRB(n912), .SETB(1'b1), .Q(\IDinst/RegFile[23][26] ) );
  dffascs1 \IDinst/RegFile_reg[24][26]  ( .DIN(\IDinst/n5044 ), .CLK(clk), 
        .CLRB(n912), .SETB(1'b1), .Q(\IDinst/RegFile[24][26] ) );
  dffascs1 \IDinst/RegFile_reg[25][26]  ( .DIN(\IDinst/n5043 ), .CLK(clk), 
        .CLRB(n912), .SETB(1'b1), .Q(\IDinst/RegFile[25][26] ) );
  dffascs1 \IDinst/RegFile_reg[26][26]  ( .DIN(\IDinst/n5042 ), .CLK(clk), 
        .CLRB(n912), .SETB(1'b1), .Q(\IDinst/RegFile[26][26] ) );
  dffascs1 \IDinst/RegFile_reg[27][26]  ( .DIN(\IDinst/n5041 ), .CLK(clk), 
        .CLRB(n913), .SETB(1'b1), .Q(\IDinst/RegFile[27][26] ) );
  dffascs1 \IDinst/RegFile_reg[28][26]  ( .DIN(\IDinst/n5040 ), .CLK(clk), 
        .CLRB(n913), .SETB(1'b1), .Q(\IDinst/RegFile[28][26] ) );
  dffascs1 \IDinst/RegFile_reg[29][26]  ( .DIN(\IDinst/n5039 ), .CLK(clk), 
        .CLRB(n913), .SETB(1'b1), .Q(\IDinst/RegFile[29][26] ) );
  dffascs1 \IDinst/RegFile_reg[30][26]  ( .DIN(\IDinst/n5038 ), .CLK(clk), 
        .CLRB(n913), .SETB(1'b1), .Q(\IDinst/RegFile[30][26] ) );
  dffascs1 \IDinst/RegFile_reg[31][26]  ( .DIN(\IDinst/n5037 ), .CLK(clk), 
        .CLRB(n913), .SETB(1'b1), .Q(\IDinst/RegFile[31][26] ) );
  dffascs1 \IDinst/RegFile_reg[0][27]  ( .DIN(\IDinst/n5036 ), .CLK(clk), 
        .CLRB(n906), .SETB(1'b1), .Q(\IDinst/RegFile[0][27] ) );
  dffascs1 \IDinst/RegFile_reg[1][27]  ( .DIN(\IDinst/n5035 ), .CLK(clk), 
        .CLRB(n906), .SETB(1'b1), .Q(\IDinst/RegFile[1][27] ) );
  dffascs1 \IDinst/RegFile_reg[2][27]  ( .DIN(\IDinst/n5034 ), .CLK(clk), 
        .CLRB(n907), .SETB(1'b1), .Q(\IDinst/RegFile[2][27] ) );
  dffascs1 \IDinst/RegFile_reg[3][27]  ( .DIN(\IDinst/n5033 ), .CLK(clk), 
        .CLRB(n907), .SETB(1'b1), .Q(\IDinst/RegFile[3][27] ) );
  dffascs1 \IDinst/RegFile_reg[4][27]  ( .DIN(\IDinst/n5032 ), .CLK(clk), 
        .CLRB(n907), .SETB(1'b1), .Q(\IDinst/RegFile[4][27] ) );
  dffascs1 \IDinst/RegFile_reg[5][27]  ( .DIN(\IDinst/n5031 ), .CLK(clk), 
        .CLRB(n907), .SETB(1'b1), .Q(\IDinst/RegFile[5][27] ) );
  dffascs1 \IDinst/RegFile_reg[6][27]  ( .DIN(\IDinst/n5030 ), .CLK(clk), 
        .CLRB(n907), .SETB(1'b1), .Q(\IDinst/RegFile[6][27] ) );
  dffascs1 \IDinst/RegFile_reg[7][27]  ( .DIN(\IDinst/n5029 ), .CLK(clk), 
        .CLRB(n907), .SETB(1'b1), .Q(\IDinst/RegFile[7][27] ) );
  dffascs1 \IDinst/RegFile_reg[8][27]  ( .DIN(\IDinst/n5028 ), .CLK(clk), 
        .CLRB(n907), .SETB(1'b1), .Q(\IDinst/RegFile[8][27] ) );
  dffascs1 \IDinst/RegFile_reg[9][27]  ( .DIN(\IDinst/n5027 ), .CLK(clk), 
        .CLRB(n907), .SETB(1'b1), .Q(\IDinst/RegFile[9][27] ) );
  dffascs1 \IDinst/RegFile_reg[10][27]  ( .DIN(\IDinst/n5026 ), .CLK(clk), 
        .CLRB(n907), .SETB(1'b1), .Q(\IDinst/RegFile[10][27] ) );
  dffascs1 \IDinst/RegFile_reg[11][27]  ( .DIN(\IDinst/n5025 ), .CLK(clk), 
        .CLRB(n907), .SETB(1'b1), .Q(\IDinst/RegFile[11][27] ) );
  dffascs1 \IDinst/RegFile_reg[12][27]  ( .DIN(\IDinst/n5024 ), .CLK(clk), 
        .CLRB(n908), .SETB(1'b1), .Q(\IDinst/RegFile[12][27] ) );
  dffascs1 \IDinst/RegFile_reg[13][27]  ( .DIN(\IDinst/n5023 ), .CLK(clk), 
        .CLRB(n908), .SETB(1'b1), .Q(\IDinst/RegFile[13][27] ) );
  dffascs1 \IDinst/RegFile_reg[14][27]  ( .DIN(\IDinst/n5022 ), .CLK(clk), 
        .CLRB(n908), .SETB(1'b1), .Q(\IDinst/RegFile[14][27] ) );
  dffascs1 \IDinst/RegFile_reg[15][27]  ( .DIN(\IDinst/n5021 ), .CLK(clk), 
        .CLRB(n908), .SETB(1'b1), .Q(\IDinst/RegFile[15][27] ) );
  dffascs1 \IDinst/RegFile_reg[16][27]  ( .DIN(\IDinst/n5020 ), .CLK(clk), 
        .CLRB(n908), .SETB(1'b1), .Q(\IDinst/RegFile[16][27] ) );
  dffascs1 \IDinst/RegFile_reg[17][27]  ( .DIN(\IDinst/n5019 ), .CLK(clk), 
        .CLRB(n908), .SETB(1'b1), .Q(\IDinst/RegFile[17][27] ) );
  dffascs1 \IDinst/RegFile_reg[18][27]  ( .DIN(\IDinst/n5018 ), .CLK(clk), 
        .CLRB(n908), .SETB(1'b1), .Q(\IDinst/RegFile[18][27] ) );
  dffascs1 \IDinst/RegFile_reg[19][27]  ( .DIN(\IDinst/n5017 ), .CLK(clk), 
        .CLRB(n908), .SETB(1'b1), .Q(\IDinst/RegFile[19][27] ) );
  dffascs1 \IDinst/RegFile_reg[20][27]  ( .DIN(\IDinst/n5016 ), .CLK(clk), 
        .CLRB(n908), .SETB(1'b1), .Q(\IDinst/RegFile[20][27] ) );
  dffascs1 \IDinst/RegFile_reg[21][27]  ( .DIN(\IDinst/n5015 ), .CLK(clk), 
        .CLRB(n908), .SETB(1'b1), .Q(\IDinst/RegFile[21][27] ) );
  dffascs1 \IDinst/RegFile_reg[22][27]  ( .DIN(\IDinst/n5014 ), .CLK(clk), 
        .CLRB(n909), .SETB(1'b1), .Q(\IDinst/RegFile[22][27] ) );
  dffascs1 \IDinst/RegFile_reg[23][27]  ( .DIN(\IDinst/n5013 ), .CLK(clk), 
        .CLRB(n909), .SETB(1'b1), .Q(\IDinst/RegFile[23][27] ) );
  dffascs1 \IDinst/RegFile_reg[24][27]  ( .DIN(\IDinst/n5012 ), .CLK(clk), 
        .CLRB(n909), .SETB(1'b1), .Q(\IDinst/RegFile[24][27] ) );
  dffascs1 \IDinst/RegFile_reg[25][27]  ( .DIN(\IDinst/n5011 ), .CLK(clk), 
        .CLRB(n909), .SETB(1'b1), .Q(\IDinst/RegFile[25][27] ) );
  dffascs1 \IDinst/RegFile_reg[26][27]  ( .DIN(\IDinst/n5010 ), .CLK(clk), 
        .CLRB(n909), .SETB(1'b1), .Q(\IDinst/RegFile[26][27] ) );
  dffascs1 \IDinst/RegFile_reg[27][27]  ( .DIN(\IDinst/n5009 ), .CLK(clk), 
        .CLRB(n909), .SETB(1'b1), .Q(\IDinst/RegFile[27][27] ) );
  dffascs1 \IDinst/RegFile_reg[28][27]  ( .DIN(\IDinst/n5008 ), .CLK(clk), 
        .CLRB(n909), .SETB(1'b1), .Q(\IDinst/RegFile[28][27] ) );
  dffascs1 \IDinst/RegFile_reg[29][27]  ( .DIN(\IDinst/n5007 ), .CLK(clk), 
        .CLRB(n909), .SETB(1'b1), .Q(\IDinst/RegFile[29][27] ) );
  dffascs1 \IDinst/RegFile_reg[30][27]  ( .DIN(\IDinst/n5006 ), .CLK(clk), 
        .CLRB(n909), .SETB(1'b1), .Q(\IDinst/RegFile[30][27] ) );
  dffascs1 \IDinst/RegFile_reg[31][27]  ( .DIN(\IDinst/n5005 ), .CLK(clk), 
        .CLRB(n909), .SETB(1'b1), .Q(\IDinst/RegFile[31][27] ) );
  dffascs1 \IDinst/RegFile_reg[0][28]  ( .DIN(\IDinst/n5004 ), .CLK(clk), 
        .CLRB(n918), .SETB(1'b1), .Q(\IDinst/RegFile[0][28] ) );
  dffascs1 \IDinst/RegFile_reg[1][28]  ( .DIN(\IDinst/n5003 ), .CLK(clk), 
        .CLRB(n919), .SETB(1'b1), .Q(\IDinst/RegFile[1][28] ) );
  dffascs1 \IDinst/RegFile_reg[2][28]  ( .DIN(\IDinst/n5002 ), .CLK(clk), 
        .CLRB(n919), .SETB(1'b1), .Q(\IDinst/RegFile[2][28] ) );
  dffascs1 \IDinst/RegFile_reg[3][28]  ( .DIN(\IDinst/n5001 ), .CLK(clk), 
        .CLRB(n919), .SETB(1'b1), .Q(\IDinst/RegFile[3][28] ) );
  dffascs1 \IDinst/RegFile_reg[4][28]  ( .DIN(\IDinst/n5000 ), .CLK(clk), 
        .CLRB(n919), .SETB(1'b1), .Q(\IDinst/RegFile[4][28] ) );
  dffascs1 \IDinst/RegFile_reg[5][28]  ( .DIN(\IDinst/n4999 ), .CLK(clk), 
        .CLRB(n919), .SETB(1'b1), .Q(\IDinst/RegFile[5][28] ) );
  dffascs1 \IDinst/RegFile_reg[6][28]  ( .DIN(\IDinst/n4998 ), .CLK(clk), 
        .CLRB(n919), .SETB(1'b1), .Q(\IDinst/RegFile[6][28] ) );
  dffascs1 \IDinst/RegFile_reg[7][28]  ( .DIN(\IDinst/n4997 ), .CLK(clk), 
        .CLRB(n919), .SETB(1'b1), .Q(\IDinst/RegFile[7][28] ) );
  dffascs1 \IDinst/RegFile_reg[8][28]  ( .DIN(\IDinst/n4996 ), .CLK(clk), 
        .CLRB(n919), .SETB(1'b1), .Q(\IDinst/RegFile[8][28] ) );
  dffascs1 \IDinst/RegFile_reg[9][28]  ( .DIN(\IDinst/n4995 ), .CLK(clk), 
        .CLRB(n919), .SETB(1'b1), .Q(\IDinst/RegFile[9][28] ) );
  dffascs1 \IDinst/RegFile_reg[10][28]  ( .DIN(\IDinst/n4994 ), .CLK(clk), 
        .CLRB(n919), .SETB(1'b1), .Q(\IDinst/RegFile[10][28] ) );
  dffascs1 \IDinst/RegFile_reg[11][28]  ( .DIN(\IDinst/n4993 ), .CLK(clk), 
        .CLRB(n920), .SETB(1'b1), .Q(\IDinst/RegFile[11][28] ) );
  dffascs1 \IDinst/RegFile_reg[12][28]  ( .DIN(\IDinst/n4992 ), .CLK(clk), 
        .CLRB(n920), .SETB(1'b1), .Q(\IDinst/RegFile[12][28] ) );
  dffascs1 \IDinst/RegFile_reg[13][28]  ( .DIN(\IDinst/n4991 ), .CLK(clk), 
        .CLRB(n920), .SETB(1'b1), .Q(\IDinst/RegFile[13][28] ) );
  dffascs1 \IDinst/RegFile_reg[14][28]  ( .DIN(\IDinst/n4990 ), .CLK(clk), 
        .CLRB(n920), .SETB(1'b1), .Q(\IDinst/RegFile[14][28] ) );
  dffascs1 \IDinst/RegFile_reg[15][28]  ( .DIN(\IDinst/n4989 ), .CLK(clk), 
        .CLRB(n920), .SETB(1'b1), .Q(\IDinst/RegFile[15][28] ) );
  dffascs1 \IDinst/RegFile_reg[16][28]  ( .DIN(\IDinst/n4988 ), .CLK(clk), 
        .CLRB(n920), .SETB(1'b1), .Q(\IDinst/RegFile[16][28] ) );
  dffascs1 \IDinst/RegFile_reg[17][28]  ( .DIN(\IDinst/n4987 ), .CLK(clk), 
        .CLRB(n920), .SETB(1'b1), .Q(\IDinst/RegFile[17][28] ) );
  dffascs1 \IDinst/RegFile_reg[18][28]  ( .DIN(\IDinst/n4986 ), .CLK(clk), 
        .CLRB(n920), .SETB(1'b1), .Q(\IDinst/RegFile[18][28] ) );
  dffascs1 \IDinst/RegFile_reg[19][28]  ( .DIN(\IDinst/n4985 ), .CLK(clk), 
        .CLRB(n920), .SETB(1'b1), .Q(\IDinst/RegFile[19][28] ) );
  dffascs1 \IDinst/RegFile_reg[20][28]  ( .DIN(\IDinst/n4984 ), .CLK(clk), 
        .CLRB(n920), .SETB(1'b1), .Q(\IDinst/RegFile[20][28] ) );
  dffascs1 \IDinst/RegFile_reg[21][28]  ( .DIN(\IDinst/n4983 ), .CLK(clk), 
        .CLRB(n921), .SETB(1'b1), .Q(\IDinst/RegFile[21][28] ) );
  dffascs1 \IDinst/RegFile_reg[22][28]  ( .DIN(\IDinst/n4982 ), .CLK(clk), 
        .CLRB(n921), .SETB(1'b1), .Q(\IDinst/RegFile[22][28] ) );
  dffascs1 \IDinst/RegFile_reg[23][28]  ( .DIN(\IDinst/n4981 ), .CLK(clk), 
        .CLRB(n921), .SETB(1'b1), .Q(\IDinst/RegFile[23][28] ) );
  dffascs1 \IDinst/RegFile_reg[24][28]  ( .DIN(\IDinst/n4980 ), .CLK(clk), 
        .CLRB(n921), .SETB(1'b1), .Q(\IDinst/RegFile[24][28] ) );
  dffascs1 \IDinst/RegFile_reg[25][28]  ( .DIN(\IDinst/n4979 ), .CLK(clk), 
        .CLRB(n921), .SETB(1'b1), .Q(\IDinst/RegFile[25][28] ) );
  dffascs1 \IDinst/RegFile_reg[26][28]  ( .DIN(\IDinst/n4978 ), .CLK(clk), 
        .CLRB(n921), .SETB(1'b1), .Q(\IDinst/RegFile[26][28] ) );
  dffascs1 \IDinst/RegFile_reg[27][28]  ( .DIN(\IDinst/n4977 ), .CLK(clk), 
        .CLRB(n921), .SETB(1'b1), .Q(\IDinst/RegFile[27][28] ) );
  dffascs1 \IDinst/RegFile_reg[28][28]  ( .DIN(\IDinst/n4976 ), .CLK(clk), 
        .CLRB(n921), .SETB(1'b1), .Q(\IDinst/RegFile[28][28] ) );
  dffascs1 \IDinst/RegFile_reg[29][28]  ( .DIN(\IDinst/n4975 ), .CLK(clk), 
        .CLRB(n921), .SETB(1'b1), .Q(\IDinst/RegFile[29][28] ) );
  dffascs1 \IDinst/RegFile_reg[30][28]  ( .DIN(\IDinst/n4974 ), .CLK(clk), 
        .CLRB(n921), .SETB(1'b1), .Q(\IDinst/RegFile[30][28] ) );
  dffascs1 \IDinst/RegFile_reg[31][28]  ( .DIN(\IDinst/n4973 ), .CLK(clk), 
        .CLRB(n922), .SETB(1'b1), .Q(\IDinst/RegFile[31][28] ) );
  dffascs1 \IDinst/RegFile_reg[0][29]  ( .DIN(\IDinst/n4972 ), .CLK(clk), 
        .CLRB(n962), .SETB(1'b1), .Q(\IDinst/RegFile[0][29] ) );
  dffascs1 \IDinst/RegFile_reg[1][29]  ( .DIN(\IDinst/n4971 ), .CLK(clk), 
        .CLRB(n936), .SETB(1'b1), .Q(\IDinst/RegFile[1][29] ) );
  dffascs1 \IDinst/RegFile_reg[2][29]  ( .DIN(\IDinst/n4970 ), .CLK(clk), 
        .CLRB(n937), .SETB(1'b1), .Q(\IDinst/RegFile[2][29] ) );
  dffascs1 \IDinst/RegFile_reg[3][29]  ( .DIN(\IDinst/n4969 ), .CLK(clk), 
        .CLRB(n937), .SETB(1'b1), .Q(\IDinst/RegFile[3][29] ) );
  dffascs1 \IDinst/RegFile_reg[4][29]  ( .DIN(\IDinst/n4968 ), .CLK(clk), 
        .CLRB(n937), .SETB(1'b1), .Q(\IDinst/RegFile[4][29] ) );
  dffascs1 \IDinst/RegFile_reg[5][29]  ( .DIN(\IDinst/n4967 ), .CLK(clk), 
        .CLRB(n938), .SETB(1'b1), .Q(\IDinst/RegFile[5][29] ) );
  dffascs1 \IDinst/RegFile_reg[6][29]  ( .DIN(\IDinst/n4966 ), .CLK(clk), 
        .CLRB(n938), .SETB(1'b1), .Q(\IDinst/RegFile[6][29] ) );
  dffascs1 \IDinst/RegFile_reg[7][29]  ( .DIN(\IDinst/n4965 ), .CLK(clk), 
        .CLRB(n939), .SETB(1'b1), .Q(\IDinst/RegFile[7][29] ) );
  dffascs1 \IDinst/RegFile_reg[8][29]  ( .DIN(\IDinst/n4964 ), .CLK(clk), 
        .CLRB(n933), .SETB(1'b1), .Q(\IDinst/RegFile[8][29] ) );
  dffascs1 \IDinst/RegFile_reg[9][29]  ( .DIN(\IDinst/n4963 ), .CLK(clk), 
        .CLRB(n933), .SETB(1'b1), .Q(\IDinst/RegFile[9][29] ) );
  dffascs1 \IDinst/RegFile_reg[10][29]  ( .DIN(\IDinst/n4962 ), .CLK(clk), 
        .CLRB(n934), .SETB(1'b1), .Q(\IDinst/RegFile[10][29] ) );
  dffascs1 \IDinst/RegFile_reg[11][29]  ( .DIN(\IDinst/n4961 ), .CLK(clk), 
        .CLRB(n934), .SETB(1'b1), .Q(\IDinst/RegFile[11][29] ) );
  dffascs1 \IDinst/RegFile_reg[12][29]  ( .DIN(\IDinst/n4960 ), .CLK(clk), 
        .CLRB(n935), .SETB(1'b1), .Q(\IDinst/RegFile[12][29] ) );
  dffascs1 \IDinst/RegFile_reg[13][29]  ( .DIN(\IDinst/n4959 ), .CLK(clk), 
        .CLRB(n935), .SETB(1'b1), .Q(\IDinst/RegFile[13][29] ) );
  dffascs1 \IDinst/RegFile_reg[14][29]  ( .DIN(\IDinst/n4958 ), .CLK(clk), 
        .CLRB(n935), .SETB(1'b1), .Q(\IDinst/RegFile[14][29] ) );
  dffascs1 \IDinst/RegFile_reg[15][29]  ( .DIN(\IDinst/n4957 ), .CLK(clk), 
        .CLRB(n936), .SETB(1'b1), .Q(\IDinst/RegFile[15][29] ) );
  dffascs1 \IDinst/RegFile_reg[16][29]  ( .DIN(\IDinst/n4956 ), .CLK(clk), 
        .CLRB(n930), .SETB(1'b1), .Q(\IDinst/RegFile[16][29] ) );
  dffascs1 \IDinst/RegFile_reg[17][29]  ( .DIN(\IDinst/n4955 ), .CLK(clk), 
        .CLRB(n930), .SETB(1'b1), .Q(\IDinst/RegFile[17][29] ) );
  dffascs1 \IDinst/RegFile_reg[18][29]  ( .DIN(\IDinst/n4954 ), .CLK(clk), 
        .CLRB(n931), .SETB(1'b1), .Q(\IDinst/RegFile[18][29] ) );
  dffascs1 \IDinst/RegFile_reg[19][29]  ( .DIN(\IDinst/n4953 ), .CLK(clk), 
        .CLRB(n931), .SETB(1'b1), .Q(\IDinst/RegFile[19][29] ) );
  dffascs1 \IDinst/RegFile_reg[20][29]  ( .DIN(\IDinst/n4952 ), .CLK(clk), 
        .CLRB(n931), .SETB(1'b1), .Q(\IDinst/RegFile[20][29] ) );
  dffascs1 \IDinst/RegFile_reg[21][29]  ( .DIN(\IDinst/n4951 ), .CLK(clk), 
        .CLRB(n932), .SETB(1'b1), .Q(\IDinst/RegFile[21][29] ) );
  dffascs1 \IDinst/RegFile_reg[22][29]  ( .DIN(\IDinst/n4950 ), .CLK(clk), 
        .CLRB(n932), .SETB(1'b1), .Q(\IDinst/RegFile[22][29] ) );
  dffascs1 \IDinst/RegFile_reg[23][29]  ( .DIN(\IDinst/n4949 ), .CLK(clk), 
        .CLRB(n933), .SETB(1'b1), .Q(\IDinst/RegFile[23][29] ) );
  dffascs1 \IDinst/RegFile_reg[24][29]  ( .DIN(\IDinst/n4948 ), .CLK(clk), 
        .CLRB(n927), .SETB(1'b1), .Q(\IDinst/RegFile[24][29] ) );
  dffascs1 \IDinst/RegFile_reg[25][29]  ( .DIN(\IDinst/n4947 ), .CLK(clk), 
        .CLRB(n927), .SETB(1'b1), .Q(\IDinst/RegFile[25][29] ) );
  dffascs1 \IDinst/RegFile_reg[26][29]  ( .DIN(\IDinst/n4946 ), .CLK(clk), 
        .CLRB(n927), .SETB(1'b1), .Q(\IDinst/RegFile[26][29] ) );
  dffascs1 \IDinst/RegFile_reg[27][29]  ( .DIN(\IDinst/n4945 ), .CLK(clk), 
        .CLRB(n928), .SETB(1'b1), .Q(\IDinst/RegFile[27][29] ) );
  dffascs1 \IDinst/RegFile_reg[28][29]  ( .DIN(\IDinst/n4944 ), .CLK(clk), 
        .CLRB(n928), .SETB(1'b1), .Q(\IDinst/RegFile[28][29] ) );
  dffascs1 \IDinst/RegFile_reg[29][29]  ( .DIN(\IDinst/n4943 ), .CLK(clk), 
        .CLRB(n929), .SETB(1'b1), .Q(\IDinst/RegFile[29][29] ) );
  dffascs1 \IDinst/RegFile_reg[30][29]  ( .DIN(\IDinst/n4942 ), .CLK(clk), 
        .CLRB(n929), .SETB(1'b1), .Q(\IDinst/RegFile[30][29] ) );
  dffascs1 \IDinst/RegFile_reg[31][29]  ( .DIN(\IDinst/n4941 ), .CLK(clk), 
        .CLRB(n929), .SETB(1'b1), .Q(\IDinst/RegFile[31][29] ) );
  dffascs1 \IDinst/RegFile_reg[0][30]  ( .DIN(\IDinst/n4940 ), .CLK(clk), 
        .CLRB(n963), .SETB(1'b1), .Q(\IDinst/RegFile[0][30] ) );
  dffascs1 \IDinst/RegFile_reg[1][30]  ( .DIN(\IDinst/n4939 ), .CLK(clk), 
        .CLRB(n936), .SETB(1'b1), .Q(\IDinst/RegFile[1][30] ) );
  dffascs1 \IDinst/RegFile_reg[2][30]  ( .DIN(\IDinst/n4938 ), .CLK(clk), 
        .CLRB(n937), .SETB(1'b1), .Q(\IDinst/RegFile[2][30] ) );
  dffascs1 \IDinst/RegFile_reg[3][30]  ( .DIN(\IDinst/n4937 ), .CLK(clk), 
        .CLRB(n937), .SETB(1'b1), .Q(\IDinst/RegFile[3][30] ) );
  dffascs1 \IDinst/RegFile_reg[4][30]  ( .DIN(\IDinst/n4936 ), .CLK(clk), 
        .CLRB(n938), .SETB(1'b1), .Q(\IDinst/RegFile[4][30] ) );
  dffascs1 \IDinst/RegFile_reg[5][30]  ( .DIN(\IDinst/n4935 ), .CLK(clk), 
        .CLRB(n938), .SETB(1'b1), .Q(\IDinst/RegFile[5][30] ) );
  dffascs1 \IDinst/RegFile_reg[6][30]  ( .DIN(\IDinst/n4934 ), .CLK(clk), 
        .CLRB(n938), .SETB(1'b1), .Q(\IDinst/RegFile[6][30] ) );
  dffascs1 \IDinst/RegFile_reg[7][30]  ( .DIN(\IDinst/n4933 ), .CLK(clk), 
        .CLRB(n939), .SETB(1'b1), .Q(\IDinst/RegFile[7][30] ) );
  dffascs1 \IDinst/RegFile_reg[8][30]  ( .DIN(\IDinst/n4932 ), .CLK(clk), 
        .CLRB(n933), .SETB(1'b1), .Q(\IDinst/RegFile[8][30] ) );
  dffascs1 \IDinst/RegFile_reg[9][30]  ( .DIN(\IDinst/n4931 ), .CLK(clk), 
        .CLRB(n933), .SETB(1'b1), .Q(\IDinst/RegFile[9][30] ) );
  dffascs1 \IDinst/RegFile_reg[10][30]  ( .DIN(\IDinst/n4930 ), .CLK(clk), 
        .CLRB(n934), .SETB(1'b1), .Q(\IDinst/RegFile[10][30] ) );
  dffascs1 \IDinst/RegFile_reg[11][30]  ( .DIN(\IDinst/n4929 ), .CLK(clk), 
        .CLRB(n934), .SETB(1'b1), .Q(\IDinst/RegFile[11][30] ) );
  dffascs1 \IDinst/RegFile_reg[12][30]  ( .DIN(\IDinst/n4928 ), .CLK(clk), 
        .CLRB(n935), .SETB(1'b1), .Q(\IDinst/RegFile[12][30] ) );
  dffascs1 \IDinst/RegFile_reg[13][30]  ( .DIN(\IDinst/n4927 ), .CLK(clk), 
        .CLRB(n935), .SETB(1'b1), .Q(\IDinst/RegFile[13][30] ) );
  dffascs1 \IDinst/RegFile_reg[14][30]  ( .DIN(\IDinst/n4926 ), .CLK(clk), 
        .CLRB(n935), .SETB(1'b1), .Q(\IDinst/RegFile[14][30] ) );
  dffascs1 \IDinst/RegFile_reg[15][30]  ( .DIN(\IDinst/n4925 ), .CLK(clk), 
        .CLRB(n936), .SETB(1'b1), .Q(\IDinst/RegFile[15][30] ) );
  dffascs1 \IDinst/RegFile_reg[16][30]  ( .DIN(\IDinst/n4924 ), .CLK(clk), 
        .CLRB(n930), .SETB(1'b1), .Q(\IDinst/RegFile[16][30] ) );
  dffascs1 \IDinst/RegFile_reg[17][30]  ( .DIN(\IDinst/n4923 ), .CLK(clk), 
        .CLRB(n930), .SETB(1'b1), .Q(\IDinst/RegFile[17][30] ) );
  dffascs1 \IDinst/RegFile_reg[18][30]  ( .DIN(\IDinst/n4922 ), .CLK(clk), 
        .CLRB(n931), .SETB(1'b1), .Q(\IDinst/RegFile[18][30] ) );
  dffascs1 \IDinst/RegFile_reg[19][30]  ( .DIN(\IDinst/n4921 ), .CLK(clk), 
        .CLRB(n931), .SETB(1'b1), .Q(\IDinst/RegFile[19][30] ) );
  dffascs1 \IDinst/RegFile_reg[20][30]  ( .DIN(\IDinst/n4920 ), .CLK(clk), 
        .CLRB(n931), .SETB(1'b1), .Q(\IDinst/RegFile[20][30] ) );
  dffascs1 \IDinst/RegFile_reg[21][30]  ( .DIN(\IDinst/n4919 ), .CLK(clk), 
        .CLRB(n932), .SETB(1'b1), .Q(\IDinst/RegFile[21][30] ) );
  dffascs1 \IDinst/RegFile_reg[22][30]  ( .DIN(\IDinst/n4918 ), .CLK(clk), 
        .CLRB(n932), .SETB(1'b1), .Q(\IDinst/RegFile[22][30] ) );
  dffascs1 \IDinst/RegFile_reg[23][30]  ( .DIN(\IDinst/n4917 ), .CLK(clk), 
        .CLRB(n933), .SETB(1'b1), .Q(\IDinst/RegFile[23][30] ) );
  dffascs1 \IDinst/RegFile_reg[24][30]  ( .DIN(\IDinst/n4916 ), .CLK(clk), 
        .CLRB(n927), .SETB(1'b1), .Q(\IDinst/RegFile[24][30] ) );
  dffascs1 \IDinst/RegFile_reg[25][30]  ( .DIN(\IDinst/n4915 ), .CLK(clk), 
        .CLRB(n927), .SETB(1'b1), .Q(\IDinst/RegFile[25][30] ) );
  dffascs1 \IDinst/RegFile_reg[26][30]  ( .DIN(\IDinst/n4914 ), .CLK(clk), 
        .CLRB(n928), .SETB(1'b1), .Q(\IDinst/RegFile[26][30] ) );
  dffascs1 \IDinst/RegFile_reg[27][30]  ( .DIN(\IDinst/n4913 ), .CLK(clk), 
        .CLRB(n928), .SETB(1'b1), .Q(\IDinst/RegFile[27][30] ) );
  dffascs1 \IDinst/RegFile_reg[28][30]  ( .DIN(\IDinst/n4912 ), .CLK(clk), 
        .CLRB(n928), .SETB(1'b1), .Q(\IDinst/RegFile[28][30] ) );
  dffascs1 \IDinst/RegFile_reg[29][30]  ( .DIN(\IDinst/n4911 ), .CLK(clk), 
        .CLRB(n929), .SETB(1'b1), .Q(\IDinst/RegFile[29][30] ) );
  dffascs1 \IDinst/RegFile_reg[30][30]  ( .DIN(\IDinst/n4910 ), .CLK(clk), 
        .CLRB(n929), .SETB(1'b1), .Q(\IDinst/RegFile[30][30] ) );
  dffascs1 \IDinst/RegFile_reg[31][30]  ( .DIN(\IDinst/n4909 ), .CLK(clk), 
        .CLRB(n929), .SETB(1'b1), .Q(\IDinst/RegFile[31][30] ) );
  dffascs1 \IDinst/RegFile_reg[0][31]  ( .DIN(\IDinst/n4908 ), .CLK(clk), 
        .CLRB(n963), .SETB(1'b1), .Q(\IDinst/RegFile[0][31] ) );
  dffascs1 \IDinst/RegFile_reg[1][31]  ( .DIN(\IDinst/n4907 ), .CLK(clk), 
        .CLRB(n936), .SETB(1'b1), .Q(\IDinst/RegFile[1][31] ) );
  dffascs1 \IDinst/RegFile_reg[2][31]  ( .DIN(\IDinst/n4906 ), .CLK(clk), 
        .CLRB(n937), .SETB(1'b1), .Q(\IDinst/RegFile[2][31] ) );
  dffascs1 \IDinst/RegFile_reg[3][31]  ( .DIN(\IDinst/n4905 ), .CLK(clk), 
        .CLRB(n937), .SETB(1'b1), .Q(\IDinst/RegFile[3][31] ) );
  dffascs1 \IDinst/RegFile_reg[4][31]  ( .DIN(\IDinst/n4904 ), .CLK(clk), 
        .CLRB(n938), .SETB(1'b1), .Q(\IDinst/RegFile[4][31] ) );
  dffascs1 \IDinst/RegFile_reg[5][31]  ( .DIN(\IDinst/n4903 ), .CLK(clk), 
        .CLRB(n938), .SETB(1'b1), .Q(\IDinst/RegFile[5][31] ) );
  dffascs1 \IDinst/RegFile_reg[6][31]  ( .DIN(\IDinst/n4902 ), .CLK(clk), 
        .CLRB(n938), .SETB(1'b1), .Q(\IDinst/RegFile[6][31] ) );
  dffascs1 \IDinst/RegFile_reg[7][31]  ( .DIN(\IDinst/n4901 ), .CLK(clk), 
        .CLRB(n939), .SETB(1'b1), .Q(\IDinst/RegFile[7][31] ) );
  dffascs1 \IDinst/RegFile_reg[8][31]  ( .DIN(\IDinst/n4900 ), .CLK(clk), 
        .CLRB(n933), .SETB(1'b1), .Q(\IDinst/RegFile[8][31] ) );
  dffascs1 \IDinst/RegFile_reg[9][31]  ( .DIN(\IDinst/n4899 ), .CLK(clk), 
        .CLRB(n934), .SETB(1'b1), .Q(\IDinst/RegFile[9][31] ) );
  dffascs1 \IDinst/RegFile_reg[10][31]  ( .DIN(\IDinst/n4898 ), .CLK(clk), 
        .CLRB(n934), .SETB(1'b1), .Q(\IDinst/RegFile[10][31] ) );
  dffascs1 \IDinst/RegFile_reg[11][31]  ( .DIN(\IDinst/n4897 ), .CLK(clk), 
        .CLRB(n934), .SETB(1'b1), .Q(\IDinst/RegFile[11][31] ) );
  dffascs1 \IDinst/RegFile_reg[12][31]  ( .DIN(\IDinst/n4896 ), .CLK(clk), 
        .CLRB(n935), .SETB(1'b1), .Q(\IDinst/RegFile[12][31] ) );
  dffascs1 \IDinst/RegFile_reg[13][31]  ( .DIN(\IDinst/n4895 ), .CLK(clk), 
        .CLRB(n935), .SETB(1'b1), .Q(\IDinst/RegFile[13][31] ) );
  dffascs1 \IDinst/RegFile_reg[14][31]  ( .DIN(\IDinst/n4894 ), .CLK(clk), 
        .CLRB(n936), .SETB(1'b1), .Q(\IDinst/RegFile[14][31] ) );
  dffascs1 \IDinst/RegFile_reg[15][31]  ( .DIN(\IDinst/n4893 ), .CLK(clk), 
        .CLRB(n936), .SETB(1'b1), .Q(\IDinst/RegFile[15][31] ) );
  dffascs1 \IDinst/RegFile_reg[16][31]  ( .DIN(\IDinst/n4892 ), .CLK(clk), 
        .CLRB(n930), .SETB(1'b1), .Q(\IDinst/RegFile[16][31] ) );
  dffascs1 \IDinst/RegFile_reg[17][31]  ( .DIN(\IDinst/n4891 ), .CLK(clk), 
        .CLRB(n930), .SETB(1'b1), .Q(\IDinst/RegFile[17][31] ) );
  dffascs1 \IDinst/RegFile_reg[18][31]  ( .DIN(\IDinst/n4890 ), .CLK(clk), 
        .CLRB(n931), .SETB(1'b1), .Q(\IDinst/RegFile[18][31] ) );
  dffascs1 \IDinst/RegFile_reg[19][31]  ( .DIN(\IDinst/n4889 ), .CLK(clk), 
        .CLRB(n931), .SETB(1'b1), .Q(\IDinst/RegFile[19][31] ) );
  dffascs1 \IDinst/RegFile_reg[20][31]  ( .DIN(\IDinst/n4888 ), .CLK(clk), 
        .CLRB(n932), .SETB(1'b1), .Q(\IDinst/RegFile[20][31] ) );
  dffascs1 \IDinst/RegFile_reg[21][31]  ( .DIN(\IDinst/n4887 ), .CLK(clk), 
        .CLRB(n932), .SETB(1'b1), .Q(\IDinst/RegFile[21][31] ) );
  dffascs1 \IDinst/RegFile_reg[22][31]  ( .DIN(\IDinst/n4886 ), .CLK(clk), 
        .CLRB(n932), .SETB(1'b1), .Q(\IDinst/RegFile[22][31] ) );
  dffascs1 \IDinst/RegFile_reg[23][31]  ( .DIN(\IDinst/n4885 ), .CLK(clk), 
        .CLRB(n933), .SETB(1'b1), .Q(\IDinst/RegFile[23][31] ) );
  dffascs1 \IDinst/RegFile_reg[24][31]  ( .DIN(\IDinst/n4884 ), .CLK(clk), 
        .CLRB(n927), .SETB(1'b1), .Q(\IDinst/RegFile[24][31] ) );
  dffascs1 \IDinst/RegFile_reg[25][31]  ( .DIN(\IDinst/n4883 ), .CLK(clk), 
        .CLRB(n927), .SETB(1'b1), .Q(\IDinst/RegFile[25][31] ) );
  dffascs1 \IDinst/RegFile_reg[26][31]  ( .DIN(\IDinst/n4882 ), .CLK(clk), 
        .CLRB(n928), .SETB(1'b1), .Q(\IDinst/RegFile[26][31] ) );
  dffascs1 \IDinst/RegFile_reg[27][31]  ( .DIN(\IDinst/n4881 ), .CLK(clk), 
        .CLRB(n928), .SETB(1'b1), .Q(\IDinst/RegFile[27][31] ) );
  dffascs1 \IDinst/RegFile_reg[28][31]  ( .DIN(\IDinst/n4880 ), .CLK(clk), 
        .CLRB(n928), .SETB(1'b1), .Q(\IDinst/RegFile[28][31] ) );
  dffascs1 \IDinst/RegFile_reg[29][31]  ( .DIN(\IDinst/n4879 ), .CLK(clk), 
        .CLRB(n929), .SETB(1'b1), .Q(\IDinst/RegFile[29][31] ) );
  dffascs1 \IDinst/RegFile_reg[30][31]  ( .DIN(\IDinst/n4878 ), .CLK(clk), 
        .CLRB(n929), .SETB(1'b1), .Q(\IDinst/RegFile[30][31] ) );
  dffascs1 \IDinst/RegFile_reg[31][31]  ( .DIN(\IDinst/n4877 ), .CLK(clk), 
        .CLRB(n930), .SETB(1'b1), .Q(\IDinst/RegFile[31][31] ) );
  dffascs1 \IDinst/RegFile_reg[0][8]  ( .DIN(\IDinst/n5644 ), .CLK(clk), 
        .CLRB(n895), .SETB(1'b1), .Q(\IDinst/RegFile[0][8] ) );
  dffascs1 \IDinst/RegFile_reg[1][8]  ( .DIN(\IDinst/n5643 ), .CLK(clk), 
        .CLRB(n895), .SETB(1'b1), .Q(\IDinst/RegFile[1][8] ) );
  dffascs1 \IDinst/RegFile_reg[2][8]  ( .DIN(\IDinst/n5642 ), .CLK(clk), 
        .CLRB(n895), .SETB(1'b1), .Q(\IDinst/RegFile[2][8] ) );
  dffascs1 \IDinst/RegFile_reg[3][8]  ( .DIN(\IDinst/n5641 ), .CLK(clk), 
        .CLRB(n896), .SETB(1'b1), .Q(\IDinst/RegFile[3][8] ) );
  dffascs1 \IDinst/RegFile_reg[4][8]  ( .DIN(\IDinst/n5640 ), .CLK(clk), 
        .CLRB(n896), .SETB(1'b1), .Q(\IDinst/RegFile[4][8] ) );
  dffascs1 \IDinst/RegFile_reg[5][8]  ( .DIN(\IDinst/n5639 ), .CLK(clk), 
        .CLRB(n896), .SETB(1'b1), .Q(\IDinst/RegFile[5][8] ) );
  dffascs1 \IDinst/RegFile_reg[6][8]  ( .DIN(\IDinst/n5638 ), .CLK(clk), 
        .CLRB(n896), .SETB(1'b1), .Q(\IDinst/RegFile[6][8] ) );
  dffascs1 \IDinst/RegFile_reg[7][8]  ( .DIN(\IDinst/n5637 ), .CLK(clk), 
        .CLRB(n896), .SETB(1'b1), .Q(\IDinst/RegFile[7][8] ) );
  dffascs1 \IDinst/RegFile_reg[8][8]  ( .DIN(\IDinst/n5636 ), .CLK(clk), 
        .CLRB(n896), .SETB(1'b1), .Q(\IDinst/RegFile[8][8] ) );
  dffascs1 \IDinst/RegFile_reg[9][8]  ( .DIN(\IDinst/n5635 ), .CLK(clk), 
        .CLRB(n896), .SETB(1'b1), .Q(\IDinst/RegFile[9][8] ) );
  dffascs1 \IDinst/RegFile_reg[10][8]  ( .DIN(\IDinst/n5634 ), .CLK(clk), 
        .CLRB(n896), .SETB(1'b1), .Q(\IDinst/RegFile[10][8] ) );
  dffascs1 \IDinst/RegFile_reg[11][8]  ( .DIN(\IDinst/n5633 ), .CLK(clk), 
        .CLRB(n896), .SETB(1'b1), .Q(\IDinst/RegFile[11][8] ) );
  dffascs1 \IDinst/RegFile_reg[12][8]  ( .DIN(\IDinst/n5632 ), .CLK(clk), 
        .CLRB(n896), .SETB(1'b1), .Q(\IDinst/RegFile[12][8] ) );
  dffascs1 \IDinst/RegFile_reg[13][8]  ( .DIN(\IDinst/n5631 ), .CLK(clk), 
        .CLRB(n897), .SETB(1'b1), .Q(\IDinst/RegFile[13][8] ) );
  dffascs1 \IDinst/RegFile_reg[14][8]  ( .DIN(\IDinst/n5630 ), .CLK(clk), 
        .CLRB(n897), .SETB(1'b1), .Q(\IDinst/RegFile[14][8] ) );
  dffascs1 \IDinst/RegFile_reg[15][8]  ( .DIN(\IDinst/n5629 ), .CLK(clk), 
        .CLRB(n897), .SETB(1'b1), .Q(\IDinst/RegFile[15][8] ) );
  dffascs1 \IDinst/RegFile_reg[16][8]  ( .DIN(\IDinst/n5628 ), .CLK(clk), 
        .CLRB(n897), .SETB(1'b1), .Q(\IDinst/RegFile[16][8] ) );
  dffascs1 \IDinst/RegFile_reg[17][8]  ( .DIN(\IDinst/n5627 ), .CLK(clk), 
        .CLRB(n897), .SETB(1'b1), .Q(\IDinst/RegFile[17][8] ) );
  dffascs1 \IDinst/RegFile_reg[18][8]  ( .DIN(\IDinst/n5626 ), .CLK(clk), 
        .CLRB(n897), .SETB(1'b1), .Q(\IDinst/RegFile[18][8] ) );
  dffascs1 \IDinst/RegFile_reg[19][8]  ( .DIN(\IDinst/n5625 ), .CLK(clk), 
        .CLRB(n897), .SETB(1'b1), .Q(\IDinst/RegFile[19][8] ) );
  dffascs1 \IDinst/RegFile_reg[20][8]  ( .DIN(\IDinst/n5624 ), .CLK(clk), 
        .CLRB(n897), .SETB(1'b1), .Q(\IDinst/RegFile[20][8] ) );
  dffascs1 \IDinst/RegFile_reg[21][8]  ( .DIN(\IDinst/n5623 ), .CLK(clk), 
        .CLRB(n897), .SETB(1'b1), .Q(\IDinst/RegFile[21][8] ) );
  dffascs1 \IDinst/RegFile_reg[22][8]  ( .DIN(\IDinst/n5622 ), .CLK(clk), 
        .CLRB(n897), .SETB(1'b1), .Q(\IDinst/RegFile[22][8] ) );
  dffascs1 \IDinst/RegFile_reg[23][8]  ( .DIN(\IDinst/n5621 ), .CLK(clk), 
        .CLRB(n898), .SETB(1'b1), .Q(\IDinst/RegFile[23][8] ) );
  dffascs1 \IDinst/RegFile_reg[24][8]  ( .DIN(\IDinst/n5620 ), .CLK(clk), 
        .CLRB(n898), .SETB(1'b1), .Q(\IDinst/RegFile[24][8] ) );
  dffascs1 \IDinst/RegFile_reg[25][8]  ( .DIN(\IDinst/n5619 ), .CLK(clk), 
        .CLRB(n898), .SETB(1'b1), .Q(\IDinst/RegFile[25][8] ) );
  dffascs1 \IDinst/RegFile_reg[26][8]  ( .DIN(\IDinst/n5618 ), .CLK(clk), 
        .CLRB(n898), .SETB(1'b1), .Q(\IDinst/RegFile[26][8] ) );
  dffascs1 \IDinst/RegFile_reg[27][8]  ( .DIN(\IDinst/n5617 ), .CLK(clk), 
        .CLRB(n898), .SETB(1'b1), .Q(\IDinst/RegFile[27][8] ) );
  dffascs1 \IDinst/RegFile_reg[28][8]  ( .DIN(\IDinst/n5616 ), .CLK(clk), 
        .CLRB(n898), .SETB(1'b1), .Q(\IDinst/RegFile[28][8] ) );
  dffascs1 \IDinst/RegFile_reg[29][8]  ( .DIN(\IDinst/n5615 ), .CLK(clk), 
        .CLRB(n898), .SETB(1'b1), .Q(\IDinst/RegFile[29][8] ) );
  dffascs1 \IDinst/RegFile_reg[30][8]  ( .DIN(\IDinst/n5614 ), .CLK(clk), 
        .CLRB(n898), .SETB(1'b1), .Q(\IDinst/RegFile[30][8] ) );
  dffascs1 \IDinst/RegFile_reg[31][8]  ( .DIN(\IDinst/n5613 ), .CLK(clk), 
        .CLRB(n898), .SETB(1'b1), .Q(\IDinst/RegFile[31][8] ) );
  dffascs1 \IDinst/RegFile_reg[0][9]  ( .DIN(\IDinst/n5612 ), .CLK(clk), 
        .CLRB(n860), .SETB(1'b1), .Q(\IDinst/RegFile[0][9] ) );
  dffascs1 \IDinst/RegFile_reg[1][9]  ( .DIN(\IDinst/n5611 ), .CLK(clk), 
        .CLRB(n860), .SETB(1'b1), .Q(\IDinst/RegFile[1][9] ) );
  dffascs1 \IDinst/RegFile_reg[2][9]  ( .DIN(\IDinst/n5610 ), .CLK(clk), 
        .CLRB(n860), .SETB(1'b1), .Q(\IDinst/RegFile[2][9] ) );
  dffascs1 \IDinst/RegFile_reg[3][9]  ( .DIN(\IDinst/n5609 ), .CLK(clk), 
        .CLRB(n861), .SETB(1'b1), .Q(\IDinst/RegFile[3][9] ) );
  dffascs1 \IDinst/RegFile_reg[4][9]  ( .DIN(\IDinst/n5608 ), .CLK(clk), 
        .CLRB(n861), .SETB(1'b1), .Q(\IDinst/RegFile[4][9] ) );
  dffascs1 \IDinst/RegFile_reg[5][9]  ( .DIN(\IDinst/n5607 ), .CLK(clk), 
        .CLRB(n861), .SETB(1'b1), .Q(\IDinst/RegFile[5][9] ) );
  dffascs1 \IDinst/RegFile_reg[6][9]  ( .DIN(\IDinst/n5606 ), .CLK(clk), 
        .CLRB(n861), .SETB(1'b1), .Q(\IDinst/RegFile[6][9] ) );
  dffascs1 \IDinst/RegFile_reg[7][9]  ( .DIN(\IDinst/n5605 ), .CLK(clk), 
        .CLRB(n861), .SETB(1'b1), .Q(\IDinst/RegFile[7][9] ) );
  dffascs1 \IDinst/RegFile_reg[8][9]  ( .DIN(\IDinst/n5604 ), .CLK(clk), 
        .CLRB(n861), .SETB(1'b1), .Q(\IDinst/RegFile[8][9] ) );
  dffascs1 \IDinst/RegFile_reg[9][9]  ( .DIN(\IDinst/n5603 ), .CLK(clk), 
        .CLRB(n861), .SETB(1'b1), .Q(\IDinst/RegFile[9][9] ) );
  dffascs1 \IDinst/RegFile_reg[10][9]  ( .DIN(\IDinst/n5602 ), .CLK(clk), 
        .CLRB(n861), .SETB(1'b1), .Q(\IDinst/RegFile[10][9] ) );
  dffascs1 \IDinst/RegFile_reg[11][9]  ( .DIN(\IDinst/n5601 ), .CLK(clk), 
        .CLRB(n861), .SETB(1'b1), .Q(\IDinst/RegFile[11][9] ) );
  dffascs1 \IDinst/RegFile_reg[12][9]  ( .DIN(\IDinst/n5600 ), .CLK(clk), 
        .CLRB(n861), .SETB(1'b1), .Q(\IDinst/RegFile[12][9] ) );
  dffascs1 \IDinst/RegFile_reg[13][9]  ( .DIN(\IDinst/n5599 ), .CLK(clk), 
        .CLRB(n862), .SETB(1'b1), .Q(\IDinst/RegFile[13][9] ) );
  dffascs1 \IDinst/RegFile_reg[14][9]  ( .DIN(\IDinst/n5598 ), .CLK(clk), 
        .CLRB(n862), .SETB(1'b1), .Q(\IDinst/RegFile[14][9] ) );
  dffascs1 \IDinst/RegFile_reg[15][9]  ( .DIN(\IDinst/n5597 ), .CLK(clk), 
        .CLRB(n862), .SETB(1'b1), .Q(\IDinst/RegFile[15][9] ) );
  dffascs1 \IDinst/RegFile_reg[16][9]  ( .DIN(\IDinst/n5596 ), .CLK(clk), 
        .CLRB(n862), .SETB(1'b1), .Q(\IDinst/RegFile[16][9] ) );
  dffascs1 \IDinst/RegFile_reg[17][9]  ( .DIN(\IDinst/n5595 ), .CLK(clk), 
        .CLRB(n862), .SETB(1'b1), .Q(\IDinst/RegFile[17][9] ) );
  dffascs1 \IDinst/RegFile_reg[18][9]  ( .DIN(\IDinst/n5594 ), .CLK(clk), 
        .CLRB(n862), .SETB(1'b1), .Q(\IDinst/RegFile[18][9] ) );
  dffascs1 \IDinst/RegFile_reg[19][9]  ( .DIN(\IDinst/n5593 ), .CLK(clk), 
        .CLRB(n862), .SETB(1'b1), .Q(\IDinst/RegFile[19][9] ) );
  dffascs1 \IDinst/RegFile_reg[20][9]  ( .DIN(\IDinst/n5592 ), .CLK(clk), 
        .CLRB(n862), .SETB(1'b1), .Q(\IDinst/RegFile[20][9] ) );
  dffascs1 \IDinst/RegFile_reg[21][9]  ( .DIN(\IDinst/n5591 ), .CLK(clk), 
        .CLRB(n862), .SETB(1'b1), .Q(\IDinst/RegFile[21][9] ) );
  dffascs1 \IDinst/RegFile_reg[22][9]  ( .DIN(\IDinst/n5590 ), .CLK(clk), 
        .CLRB(n862), .SETB(1'b1), .Q(\IDinst/RegFile[22][9] ) );
  dffascs1 \IDinst/RegFile_reg[23][9]  ( .DIN(\IDinst/n5589 ), .CLK(clk), 
        .CLRB(n863), .SETB(1'b1), .Q(\IDinst/RegFile[23][9] ) );
  dffascs1 \IDinst/RegFile_reg[24][9]  ( .DIN(\IDinst/n5588 ), .CLK(clk), 
        .CLRB(n863), .SETB(1'b1), .Q(\IDinst/RegFile[24][9] ) );
  dffascs1 \IDinst/RegFile_reg[25][9]  ( .DIN(\IDinst/n5587 ), .CLK(clk), 
        .CLRB(n863), .SETB(1'b1), .Q(\IDinst/RegFile[25][9] ) );
  dffascs1 \IDinst/RegFile_reg[26][9]  ( .DIN(\IDinst/n5586 ), .CLK(clk), 
        .CLRB(n863), .SETB(1'b1), .Q(\IDinst/RegFile[26][9] ) );
  dffascs1 \IDinst/RegFile_reg[27][9]  ( .DIN(\IDinst/n5585 ), .CLK(clk), 
        .CLRB(n863), .SETB(1'b1), .Q(\IDinst/RegFile[27][9] ) );
  dffascs1 \IDinst/RegFile_reg[28][9]  ( .DIN(\IDinst/n5584 ), .CLK(clk), 
        .CLRB(n863), .SETB(1'b1), .Q(\IDinst/RegFile[28][9] ) );
  dffascs1 \IDinst/RegFile_reg[29][9]  ( .DIN(\IDinst/n5583 ), .CLK(clk), 
        .CLRB(n863), .SETB(1'b1), .Q(\IDinst/RegFile[29][9] ) );
  dffascs1 \IDinst/RegFile_reg[30][9]  ( .DIN(\IDinst/n5582 ), .CLK(clk), 
        .CLRB(n863), .SETB(1'b1), .Q(\IDinst/RegFile[30][9] ) );
  dffascs1 \IDinst/RegFile_reg[31][9]  ( .DIN(\IDinst/n5581 ), .CLK(clk), 
        .CLRB(n863), .SETB(1'b1), .Q(\IDinst/RegFile[31][9] ) );
  dffascs1 \IDinst/RegFile_reg[0][10]  ( .DIN(\IDinst/n5580 ), .CLK(clk), 
        .CLRB(n857), .SETB(1'b1), .Q(\IDinst/RegFile[0][10] ) );
  dffascs1 \IDinst/RegFile_reg[1][10]  ( .DIN(\IDinst/n5579 ), .CLK(clk), 
        .CLRB(n857), .SETB(1'b1), .Q(\IDinst/RegFile[1][10] ) );
  dffascs1 \IDinst/RegFile_reg[2][10]  ( .DIN(\IDinst/n5578 ), .CLK(clk), 
        .CLRB(n857), .SETB(1'b1), .Q(\IDinst/RegFile[2][10] ) );
  dffascs1 \IDinst/RegFile_reg[3][10]  ( .DIN(\IDinst/n5577 ), .CLK(clk), 
        .CLRB(n857), .SETB(1'b1), .Q(\IDinst/RegFile[3][10] ) );
  dffascs1 \IDinst/RegFile_reg[4][10]  ( .DIN(\IDinst/n5576 ), .CLK(clk), 
        .CLRB(n857), .SETB(1'b1), .Q(\IDinst/RegFile[4][10] ) );
  dffascs1 \IDinst/RegFile_reg[5][10]  ( .DIN(\IDinst/n5575 ), .CLK(clk), 
        .CLRB(n857), .SETB(1'b1), .Q(\IDinst/RegFile[5][10] ) );
  dffascs1 \IDinst/RegFile_reg[6][10]  ( .DIN(\IDinst/n5574 ), .CLK(clk), 
        .CLRB(n857), .SETB(1'b1), .Q(\IDinst/RegFile[6][10] ) );
  dffascs1 \IDinst/RegFile_reg[7][10]  ( .DIN(\IDinst/n5573 ), .CLK(clk), 
        .CLRB(n857), .SETB(1'b1), .Q(\IDinst/RegFile[7][10] ) );
  dffascs1 \IDinst/RegFile_reg[8][10]  ( .DIN(\IDinst/n5572 ), .CLK(clk), 
        .CLRB(n858), .SETB(1'b1), .Q(\IDinst/RegFile[8][10] ) );
  dffascs1 \IDinst/RegFile_reg[9][10]  ( .DIN(\IDinst/n5571 ), .CLK(clk), 
        .CLRB(n858), .SETB(1'b1), .Q(\IDinst/RegFile[9][10] ) );
  dffascs1 \IDinst/RegFile_reg[10][10]  ( .DIN(\IDinst/n5570 ), .CLK(clk), 
        .CLRB(n858), .SETB(1'b1), .Q(\IDinst/RegFile[10][10] ) );
  dffascs1 \IDinst/RegFile_reg[11][10]  ( .DIN(\IDinst/n5569 ), .CLK(clk), 
        .CLRB(n858), .SETB(1'b1), .Q(\IDinst/RegFile[11][10] ) );
  dffascs1 \IDinst/RegFile_reg[12][10]  ( .DIN(\IDinst/n5568 ), .CLK(clk), 
        .CLRB(n858), .SETB(1'b1), .Q(\IDinst/RegFile[12][10] ) );
  dffascs1 \IDinst/RegFile_reg[13][10]  ( .DIN(\IDinst/n5567 ), .CLK(clk), 
        .CLRB(n858), .SETB(1'b1), .Q(\IDinst/RegFile[13][10] ) );
  dffascs1 \IDinst/RegFile_reg[14][10]  ( .DIN(\IDinst/n5566 ), .CLK(clk), 
        .CLRB(n858), .SETB(1'b1), .Q(\IDinst/RegFile[14][10] ) );
  dffascs1 \IDinst/RegFile_reg[15][10]  ( .DIN(\IDinst/n5565 ), .CLK(clk), 
        .CLRB(n858), .SETB(1'b1), .Q(\IDinst/RegFile[15][10] ) );
  dffascs1 \IDinst/RegFile_reg[16][10]  ( .DIN(\IDinst/n5564 ), .CLK(clk), 
        .CLRB(n858), .SETB(1'b1), .Q(\IDinst/RegFile[16][10] ) );
  dffascs1 \IDinst/RegFile_reg[17][10]  ( .DIN(\IDinst/n5563 ), .CLK(clk), 
        .CLRB(n858), .SETB(1'b1), .Q(\IDinst/RegFile[17][10] ) );
  dffascs1 \IDinst/RegFile_reg[18][10]  ( .DIN(\IDinst/n5562 ), .CLK(clk), 
        .CLRB(n859), .SETB(1'b1), .Q(\IDinst/RegFile[18][10] ) );
  dffascs1 \IDinst/RegFile_reg[19][10]  ( .DIN(\IDinst/n5561 ), .CLK(clk), 
        .CLRB(n859), .SETB(1'b1), .Q(\IDinst/RegFile[19][10] ) );
  dffascs1 \IDinst/RegFile_reg[20][10]  ( .DIN(\IDinst/n5560 ), .CLK(clk), 
        .CLRB(n859), .SETB(1'b1), .Q(\IDinst/RegFile[20][10] ) );
  dffascs1 \IDinst/RegFile_reg[21][10]  ( .DIN(\IDinst/n5559 ), .CLK(clk), 
        .CLRB(n859), .SETB(1'b1), .Q(\IDinst/RegFile[21][10] ) );
  dffascs1 \IDinst/RegFile_reg[22][10]  ( .DIN(\IDinst/n5558 ), .CLK(clk), 
        .CLRB(n859), .SETB(1'b1), .Q(\IDinst/RegFile[22][10] ) );
  dffascs1 \IDinst/RegFile_reg[23][10]  ( .DIN(\IDinst/n5557 ), .CLK(clk), 
        .CLRB(n859), .SETB(1'b1), .Q(\IDinst/RegFile[23][10] ) );
  dffascs1 \IDinst/RegFile_reg[24][10]  ( .DIN(\IDinst/n5556 ), .CLK(clk), 
        .CLRB(n859), .SETB(1'b1), .Q(\IDinst/RegFile[24][10] ) );
  dffascs1 \IDinst/RegFile_reg[25][10]  ( .DIN(\IDinst/n5555 ), .CLK(clk), 
        .CLRB(n859), .SETB(1'b1), .Q(\IDinst/RegFile[25][10] ) );
  dffascs1 \IDinst/RegFile_reg[26][10]  ( .DIN(\IDinst/n5554 ), .CLK(clk), 
        .CLRB(n859), .SETB(1'b1), .Q(\IDinst/RegFile[26][10] ) );
  dffascs1 \IDinst/RegFile_reg[27][10]  ( .DIN(\IDinst/n5553 ), .CLK(clk), 
        .CLRB(n859), .SETB(1'b1), .Q(\IDinst/RegFile[27][10] ) );
  dffascs1 \IDinst/RegFile_reg[28][10]  ( .DIN(\IDinst/n5552 ), .CLK(clk), 
        .CLRB(n860), .SETB(1'b1), .Q(\IDinst/RegFile[28][10] ) );
  dffascs1 \IDinst/RegFile_reg[29][10]  ( .DIN(\IDinst/n5551 ), .CLK(clk), 
        .CLRB(n860), .SETB(1'b1), .Q(\IDinst/RegFile[29][10] ) );
  dffascs1 \IDinst/RegFile_reg[30][10]  ( .DIN(\IDinst/n5550 ), .CLK(clk), 
        .CLRB(n860), .SETB(1'b1), .Q(\IDinst/RegFile[30][10] ) );
  dffascs1 \IDinst/RegFile_reg[31][10]  ( .DIN(\IDinst/n5549 ), .CLK(clk), 
        .CLRB(n860), .SETB(1'b1), .Q(\IDinst/RegFile[31][10] ) );
  dffascs1 \IDinst/RegFile_reg[0][11]  ( .DIN(\IDinst/n5548 ), .CLK(clk), 
        .CLRB(n892), .SETB(1'b1), .Q(\IDinst/RegFile[0][11] ) );
  dffascs1 \IDinst/RegFile_reg[1][11]  ( .DIN(\IDinst/n5547 ), .CLK(clk), 
        .CLRB(n892), .SETB(1'b1), .Q(\IDinst/RegFile[1][11] ) );
  dffascs1 \IDinst/RegFile_reg[2][11]  ( .DIN(\IDinst/n5546 ), .CLK(clk), 
        .CLRB(n892), .SETB(1'b1), .Q(\IDinst/RegFile[2][11] ) );
  dffascs1 \IDinst/RegFile_reg[3][11]  ( .DIN(\IDinst/n5545 ), .CLK(clk), 
        .CLRB(n892), .SETB(1'b1), .Q(\IDinst/RegFile[3][11] ) );
  dffascs1 \IDinst/RegFile_reg[4][11]  ( .DIN(\IDinst/n5544 ), .CLK(clk), 
        .CLRB(n892), .SETB(1'b1), .Q(\IDinst/RegFile[4][11] ) );
  dffascs1 \IDinst/RegFile_reg[5][11]  ( .DIN(\IDinst/n5543 ), .CLK(clk), 
        .CLRB(n892), .SETB(1'b1), .Q(\IDinst/RegFile[5][11] ) );
  dffascs1 \IDinst/RegFile_reg[6][11]  ( .DIN(\IDinst/n5542 ), .CLK(clk), 
        .CLRB(n892), .SETB(1'b1), .Q(\IDinst/RegFile[6][11] ) );
  dffascs1 \IDinst/RegFile_reg[7][11]  ( .DIN(\IDinst/n5541 ), .CLK(clk), 
        .CLRB(n892), .SETB(1'b1), .Q(\IDinst/RegFile[7][11] ) );
  dffascs1 \IDinst/RegFile_reg[8][11]  ( .DIN(\IDinst/n5540 ), .CLK(clk), 
        .CLRB(n892), .SETB(1'b1), .Q(\IDinst/RegFile[8][11] ) );
  dffascs1 \IDinst/RegFile_reg[9][11]  ( .DIN(\IDinst/n5539 ), .CLK(clk), 
        .CLRB(n893), .SETB(1'b1), .Q(\IDinst/RegFile[9][11] ) );
  dffascs1 \IDinst/RegFile_reg[10][11]  ( .DIN(\IDinst/n5538 ), .CLK(clk), 
        .CLRB(n893), .SETB(1'b1), .Q(\IDinst/RegFile[10][11] ) );
  dffascs1 \IDinst/RegFile_reg[11][11]  ( .DIN(\IDinst/n5537 ), .CLK(clk), 
        .CLRB(n893), .SETB(1'b1), .Q(\IDinst/RegFile[11][11] ) );
  dffascs1 \IDinst/RegFile_reg[12][11]  ( .DIN(\IDinst/n5536 ), .CLK(clk), 
        .CLRB(n893), .SETB(1'b1), .Q(\IDinst/RegFile[12][11] ) );
  dffascs1 \IDinst/RegFile_reg[13][11]  ( .DIN(\IDinst/n5535 ), .CLK(clk), 
        .CLRB(n893), .SETB(1'b1), .Q(\IDinst/RegFile[13][11] ) );
  dffascs1 \IDinst/RegFile_reg[14][11]  ( .DIN(\IDinst/n5534 ), .CLK(clk), 
        .CLRB(n893), .SETB(1'b1), .Q(\IDinst/RegFile[14][11] ) );
  dffascs1 \IDinst/RegFile_reg[15][11]  ( .DIN(\IDinst/n5533 ), .CLK(clk), 
        .CLRB(n893), .SETB(1'b1), .Q(\IDinst/RegFile[15][11] ) );
  dffascs1 \IDinst/RegFile_reg[16][11]  ( .DIN(\IDinst/n5532 ), .CLK(clk), 
        .CLRB(n893), .SETB(1'b1), .Q(\IDinst/RegFile[16][11] ) );
  dffascs1 \IDinst/RegFile_reg[17][11]  ( .DIN(\IDinst/n5531 ), .CLK(clk), 
        .CLRB(n893), .SETB(1'b1), .Q(\IDinst/RegFile[17][11] ) );
  dffascs1 \IDinst/RegFile_reg[18][11]  ( .DIN(\IDinst/n5530 ), .CLK(clk), 
        .CLRB(n893), .SETB(1'b1), .Q(\IDinst/RegFile[18][11] ) );
  dffascs1 \IDinst/RegFile_reg[19][11]  ( .DIN(\IDinst/n5529 ), .CLK(clk), 
        .CLRB(n894), .SETB(1'b1), .Q(\IDinst/RegFile[19][11] ) );
  dffascs1 \IDinst/RegFile_reg[20][11]  ( .DIN(\IDinst/n5528 ), .CLK(clk), 
        .CLRB(n894), .SETB(1'b1), .Q(\IDinst/RegFile[20][11] ) );
  dffascs1 \IDinst/RegFile_reg[21][11]  ( .DIN(\IDinst/n5527 ), .CLK(clk), 
        .CLRB(n894), .SETB(1'b1), .Q(\IDinst/RegFile[21][11] ) );
  dffascs1 \IDinst/RegFile_reg[22][11]  ( .DIN(\IDinst/n5526 ), .CLK(clk), 
        .CLRB(n894), .SETB(1'b1), .Q(\IDinst/RegFile[22][11] ) );
  dffascs1 \IDinst/RegFile_reg[23][11]  ( .DIN(\IDinst/n5525 ), .CLK(clk), 
        .CLRB(n894), .SETB(1'b1), .Q(\IDinst/RegFile[23][11] ) );
  dffascs1 \IDinst/RegFile_reg[24][11]  ( .DIN(\IDinst/n5524 ), .CLK(clk), 
        .CLRB(n894), .SETB(1'b1), .Q(\IDinst/RegFile[24][11] ) );
  dffascs1 \IDinst/RegFile_reg[25][11]  ( .DIN(\IDinst/n5523 ), .CLK(clk), 
        .CLRB(n894), .SETB(1'b1), .Q(\IDinst/RegFile[25][11] ) );
  dffascs1 \IDinst/RegFile_reg[26][11]  ( .DIN(\IDinst/n5522 ), .CLK(clk), 
        .CLRB(n894), .SETB(1'b1), .Q(\IDinst/RegFile[26][11] ) );
  dffascs1 \IDinst/RegFile_reg[27][11]  ( .DIN(\IDinst/n5521 ), .CLK(clk), 
        .CLRB(n894), .SETB(1'b1), .Q(\IDinst/RegFile[27][11] ) );
  dffascs1 \IDinst/RegFile_reg[28][11]  ( .DIN(\IDinst/n5520 ), .CLK(clk), 
        .CLRB(n894), .SETB(1'b1), .Q(\IDinst/RegFile[28][11] ) );
  dffascs1 \IDinst/RegFile_reg[29][11]  ( .DIN(\IDinst/n5519 ), .CLK(clk), 
        .CLRB(n895), .SETB(1'b1), .Q(\IDinst/RegFile[29][11] ) );
  dffascs1 \IDinst/RegFile_reg[30][11]  ( .DIN(\IDinst/n5518 ), .CLK(clk), 
        .CLRB(n895), .SETB(1'b1), .Q(\IDinst/RegFile[30][11] ) );
  dffascs1 \IDinst/RegFile_reg[31][11]  ( .DIN(\IDinst/n5517 ), .CLK(clk), 
        .CLRB(n895), .SETB(1'b1), .Q(\IDinst/RegFile[31][11] ) );
  dffascs1 \IDinst/RegFile_reg[0][12]  ( .DIN(\IDinst/n5516 ), .CLK(clk), 
        .CLRB(n914), .SETB(1'b1), .Q(\IDinst/RegFile[0][12] ) );
  dffascs1 \IDinst/RegFile_reg[1][12]  ( .DIN(\IDinst/n5515 ), .CLK(clk), 
        .CLRB(n914), .SETB(1'b1), .Q(\IDinst/RegFile[1][12] ) );
  dffascs1 \IDinst/RegFile_reg[2][12]  ( .DIN(\IDinst/n5514 ), .CLK(clk), 
        .CLRB(n915), .SETB(1'b1), .Q(\IDinst/RegFile[2][12] ) );
  dffascs1 \IDinst/RegFile_reg[3][12]  ( .DIN(\IDinst/n5513 ), .CLK(clk), 
        .CLRB(n915), .SETB(1'b1), .Q(\IDinst/RegFile[3][12] ) );
  dffascs1 \IDinst/RegFile_reg[4][12]  ( .DIN(\IDinst/n5512 ), .CLK(clk), 
        .CLRB(n915), .SETB(1'b1), .Q(\IDinst/RegFile[4][12] ) );
  dffascs1 \IDinst/RegFile_reg[5][12]  ( .DIN(\IDinst/n5511 ), .CLK(clk), 
        .CLRB(n915), .SETB(1'b1), .Q(\IDinst/RegFile[5][12] ) );
  dffascs1 \IDinst/RegFile_reg[6][12]  ( .DIN(\IDinst/n5510 ), .CLK(clk), 
        .CLRB(n915), .SETB(1'b1), .Q(\IDinst/RegFile[6][12] ) );
  dffascs1 \IDinst/RegFile_reg[7][12]  ( .DIN(\IDinst/n5509 ), .CLK(clk), 
        .CLRB(n915), .SETB(1'b1), .Q(\IDinst/RegFile[7][12] ) );
  dffascs1 \IDinst/RegFile_reg[8][12]  ( .DIN(\IDinst/n5508 ), .CLK(clk), 
        .CLRB(n915), .SETB(1'b1), .Q(\IDinst/RegFile[8][12] ) );
  dffascs1 \IDinst/RegFile_reg[9][12]  ( .DIN(\IDinst/n5507 ), .CLK(clk), 
        .CLRB(n915), .SETB(1'b1), .Q(\IDinst/RegFile[9][12] ) );
  dffascs1 \IDinst/RegFile_reg[10][12]  ( .DIN(\IDinst/n5506 ), .CLK(clk), 
        .CLRB(n915), .SETB(1'b1), .Q(\IDinst/RegFile[10][12] ) );
  dffascs1 \IDinst/RegFile_reg[11][12]  ( .DIN(\IDinst/n5505 ), .CLK(clk), 
        .CLRB(n915), .SETB(1'b1), .Q(\IDinst/RegFile[11][12] ) );
  dffascs1 \IDinst/RegFile_reg[12][12]  ( .DIN(\IDinst/n5504 ), .CLK(clk), 
        .CLRB(n916), .SETB(1'b1), .Q(\IDinst/RegFile[12][12] ) );
  dffascs1 \IDinst/RegFile_reg[13][12]  ( .DIN(\IDinst/n5503 ), .CLK(clk), 
        .CLRB(n916), .SETB(1'b1), .Q(\IDinst/RegFile[13][12] ) );
  dffascs1 \IDinst/RegFile_reg[14][12]  ( .DIN(\IDinst/n5502 ), .CLK(clk), 
        .CLRB(n916), .SETB(1'b1), .Q(\IDinst/RegFile[14][12] ) );
  dffascs1 \IDinst/RegFile_reg[15][12]  ( .DIN(\IDinst/n5501 ), .CLK(clk), 
        .CLRB(n916), .SETB(1'b1), .Q(\IDinst/RegFile[15][12] ) );
  dffascs1 \IDinst/RegFile_reg[16][12]  ( .DIN(\IDinst/n5500 ), .CLK(clk), 
        .CLRB(n916), .SETB(1'b1), .Q(\IDinst/RegFile[16][12] ) );
  dffascs1 \IDinst/RegFile_reg[17][12]  ( .DIN(\IDinst/n5499 ), .CLK(clk), 
        .CLRB(n916), .SETB(1'b1), .Q(\IDinst/RegFile[17][12] ) );
  dffascs1 \IDinst/RegFile_reg[18][12]  ( .DIN(\IDinst/n5498 ), .CLK(clk), 
        .CLRB(n916), .SETB(1'b1), .Q(\IDinst/RegFile[18][12] ) );
  dffascs1 \IDinst/RegFile_reg[19][12]  ( .DIN(\IDinst/n5497 ), .CLK(clk), 
        .CLRB(n916), .SETB(1'b1), .Q(\IDinst/RegFile[19][12] ) );
  dffascs1 \IDinst/RegFile_reg[20][12]  ( .DIN(\IDinst/n5496 ), .CLK(clk), 
        .CLRB(n916), .SETB(1'b1), .Q(\IDinst/RegFile[20][12] ) );
  dffascs1 \IDinst/RegFile_reg[21][12]  ( .DIN(\IDinst/n5495 ), .CLK(clk), 
        .CLRB(n916), .SETB(1'b1), .Q(\IDinst/RegFile[21][12] ) );
  dffascs1 \IDinst/RegFile_reg[22][12]  ( .DIN(\IDinst/n5494 ), .CLK(clk), 
        .CLRB(n917), .SETB(1'b1), .Q(\IDinst/RegFile[22][12] ) );
  dffascs1 \IDinst/RegFile_reg[23][12]  ( .DIN(\IDinst/n5493 ), .CLK(clk), 
        .CLRB(n917), .SETB(1'b1), .Q(\IDinst/RegFile[23][12] ) );
  dffascs1 \IDinst/RegFile_reg[24][12]  ( .DIN(\IDinst/n5492 ), .CLK(clk), 
        .CLRB(n917), .SETB(1'b1), .Q(\IDinst/RegFile[24][12] ) );
  dffascs1 \IDinst/RegFile_reg[25][12]  ( .DIN(\IDinst/n5491 ), .CLK(clk), 
        .CLRB(n917), .SETB(1'b1), .Q(\IDinst/RegFile[25][12] ) );
  dffascs1 \IDinst/RegFile_reg[26][12]  ( .DIN(\IDinst/n5490 ), .CLK(clk), 
        .CLRB(n917), .SETB(1'b1), .Q(\IDinst/RegFile[26][12] ) );
  dffascs1 \IDinst/RegFile_reg[27][12]  ( .DIN(\IDinst/n5489 ), .CLK(clk), 
        .CLRB(n917), .SETB(1'b1), .Q(\IDinst/RegFile[27][12] ) );
  dffascs1 \IDinst/RegFile_reg[28][12]  ( .DIN(\IDinst/n5488 ), .CLK(clk), 
        .CLRB(n917), .SETB(1'b1), .Q(\IDinst/RegFile[28][12] ) );
  dffascs1 \IDinst/RegFile_reg[29][12]  ( .DIN(\IDinst/n5487 ), .CLK(clk), 
        .CLRB(n917), .SETB(1'b1), .Q(\IDinst/RegFile[29][12] ) );
  dffascs1 \IDinst/RegFile_reg[30][12]  ( .DIN(\IDinst/n5486 ), .CLK(clk), 
        .CLRB(n917), .SETB(1'b1), .Q(\IDinst/RegFile[30][12] ) );
  dffascs1 \IDinst/RegFile_reg[31][12]  ( .DIN(\IDinst/n5485 ), .CLK(clk), 
        .CLRB(n917), .SETB(1'b1), .Q(\IDinst/RegFile[31][12] ) );
  dffascs1 \IDinst/RegFile_reg[0][13]  ( .DIN(\IDinst/n5484 ), .CLK(clk), 
        .CLRB(n876), .SETB(1'b1), .Q(\IDinst/RegFile[0][13] ) );
  dffascs1 \IDinst/RegFile_reg[1][13]  ( .DIN(\IDinst/n5483 ), .CLK(clk), 
        .CLRB(n876), .SETB(1'b1), .Q(\IDinst/RegFile[1][13] ) );
  dffascs1 \IDinst/RegFile_reg[2][13]  ( .DIN(\IDinst/n5482 ), .CLK(clk), 
        .CLRB(n876), .SETB(1'b1), .Q(\IDinst/RegFile[2][13] ) );
  dffascs1 \IDinst/RegFile_reg[3][13]  ( .DIN(\IDinst/n5481 ), .CLK(clk), 
        .CLRB(n876), .SETB(1'b1), .Q(\IDinst/RegFile[3][13] ) );
  dffascs1 \IDinst/RegFile_reg[4][13]  ( .DIN(\IDinst/n5480 ), .CLK(clk), 
        .CLRB(n876), .SETB(1'b1), .Q(\IDinst/RegFile[4][13] ) );
  dffascs1 \IDinst/RegFile_reg[5][13]  ( .DIN(\IDinst/n5479 ), .CLK(clk), 
        .CLRB(n876), .SETB(1'b1), .Q(\IDinst/RegFile[5][13] ) );
  dffascs1 \IDinst/RegFile_reg[6][13]  ( .DIN(\IDinst/n5478 ), .CLK(clk), 
        .CLRB(n876), .SETB(1'b1), .Q(\IDinst/RegFile[6][13] ) );
  dffascs1 \IDinst/RegFile_reg[7][13]  ( .DIN(\IDinst/n5477 ), .CLK(clk), 
        .CLRB(n877), .SETB(1'b1), .Q(\IDinst/RegFile[7][13] ) );
  dffascs1 \IDinst/RegFile_reg[8][13]  ( .DIN(\IDinst/n5476 ), .CLK(clk), 
        .CLRB(n877), .SETB(1'b1), .Q(\IDinst/RegFile[8][13] ) );
  dffascs1 \IDinst/RegFile_reg[9][13]  ( .DIN(\IDinst/n5475 ), .CLK(clk), 
        .CLRB(n877), .SETB(1'b1), .Q(\IDinst/RegFile[9][13] ) );
  dffascs1 \IDinst/RegFile_reg[10][13]  ( .DIN(\IDinst/n5474 ), .CLK(clk), 
        .CLRB(n877), .SETB(1'b1), .Q(\IDinst/RegFile[10][13] ) );
  dffascs1 \IDinst/RegFile_reg[11][13]  ( .DIN(\IDinst/n5473 ), .CLK(clk), 
        .CLRB(n877), .SETB(1'b1), .Q(\IDinst/RegFile[11][13] ) );
  dffascs1 \IDinst/RegFile_reg[12][13]  ( .DIN(\IDinst/n5472 ), .CLK(clk), 
        .CLRB(n877), .SETB(1'b1), .Q(\IDinst/RegFile[12][13] ) );
  dffascs1 \IDinst/RegFile_reg[13][13]  ( .DIN(\IDinst/n5471 ), .CLK(clk), 
        .CLRB(n877), .SETB(1'b1), .Q(\IDinst/RegFile[13][13] ) );
  dffascs1 \IDinst/RegFile_reg[14][13]  ( .DIN(\IDinst/n5470 ), .CLK(clk), 
        .CLRB(n877), .SETB(1'b1), .Q(\IDinst/RegFile[14][13] ) );
  dffascs1 \IDinst/RegFile_reg[15][13]  ( .DIN(\IDinst/n5469 ), .CLK(clk), 
        .CLRB(n877), .SETB(1'b1), .Q(\IDinst/RegFile[15][13] ) );
  dffascs1 \IDinst/RegFile_reg[16][13]  ( .DIN(\IDinst/n5468 ), .CLK(clk), 
        .CLRB(n877), .SETB(1'b1), .Q(\IDinst/RegFile[16][13] ) );
  dffascs1 \IDinst/RegFile_reg[17][13]  ( .DIN(\IDinst/n5467 ), .CLK(clk), 
        .CLRB(n878), .SETB(1'b1), .Q(\IDinst/RegFile[17][13] ) );
  dffascs1 \IDinst/RegFile_reg[18][13]  ( .DIN(\IDinst/n5466 ), .CLK(clk), 
        .CLRB(n878), .SETB(1'b1), .Q(\IDinst/RegFile[18][13] ) );
  dffascs1 \IDinst/RegFile_reg[19][13]  ( .DIN(\IDinst/n5465 ), .CLK(clk), 
        .CLRB(n878), .SETB(1'b1), .Q(\IDinst/RegFile[19][13] ) );
  dffascs1 \IDinst/RegFile_reg[20][13]  ( .DIN(\IDinst/n5464 ), .CLK(clk), 
        .CLRB(n878), .SETB(1'b1), .Q(\IDinst/RegFile[20][13] ) );
  dffascs1 \IDinst/RegFile_reg[21][13]  ( .DIN(\IDinst/n5463 ), .CLK(clk), 
        .CLRB(n878), .SETB(1'b1), .Q(\IDinst/RegFile[21][13] ) );
  dffascs1 \IDinst/RegFile_reg[22][13]  ( .DIN(\IDinst/n5462 ), .CLK(clk), 
        .CLRB(n878), .SETB(1'b1), .Q(\IDinst/RegFile[22][13] ) );
  dffascs1 \IDinst/RegFile_reg[23][13]  ( .DIN(\IDinst/n5461 ), .CLK(clk), 
        .CLRB(n878), .SETB(1'b1), .Q(\IDinst/RegFile[23][13] ) );
  dffascs1 \IDinst/RegFile_reg[24][13]  ( .DIN(\IDinst/n5460 ), .CLK(clk), 
        .CLRB(n878), .SETB(1'b1), .Q(\IDinst/RegFile[24][13] ) );
  dffascs1 \IDinst/RegFile_reg[25][13]  ( .DIN(\IDinst/n5459 ), .CLK(clk), 
        .CLRB(n878), .SETB(1'b1), .Q(\IDinst/RegFile[25][13] ) );
  dffascs1 \IDinst/RegFile_reg[26][13]  ( .DIN(\IDinst/n5458 ), .CLK(clk), 
        .CLRB(n878), .SETB(1'b1), .Q(\IDinst/RegFile[26][13] ) );
  dffascs1 \IDinst/RegFile_reg[27][13]  ( .DIN(\IDinst/n5457 ), .CLK(clk), 
        .CLRB(n879), .SETB(1'b1), .Q(\IDinst/RegFile[27][13] ) );
  dffascs1 \IDinst/RegFile_reg[28][13]  ( .DIN(\IDinst/n5456 ), .CLK(clk), 
        .CLRB(n879), .SETB(1'b1), .Q(\IDinst/RegFile[28][13] ) );
  dffascs1 \IDinst/RegFile_reg[29][13]  ( .DIN(\IDinst/n5455 ), .CLK(clk), 
        .CLRB(n879), .SETB(1'b1), .Q(\IDinst/RegFile[29][13] ) );
  dffascs1 \IDinst/RegFile_reg[30][13]  ( .DIN(\IDinst/n5454 ), .CLK(clk), 
        .CLRB(n879), .SETB(1'b1), .Q(\IDinst/RegFile[30][13] ) );
  dffascs1 \IDinst/RegFile_reg[31][13]  ( .DIN(\IDinst/n5453 ), .CLK(clk), 
        .CLRB(n879), .SETB(1'b1), .Q(\IDinst/RegFile[31][13] ) );
  dffascs1 \IDinst/RegFile_reg[0][14]  ( .DIN(\IDinst/n5452 ), .CLK(clk), 
        .CLRB(n864), .SETB(1'b1), .Q(\IDinst/RegFile[0][14] ) );
  dffascs1 \IDinst/RegFile_reg[1][14]  ( .DIN(\IDinst/n5451 ), .CLK(clk), 
        .CLRB(n864), .SETB(1'b1), .Q(\IDinst/RegFile[1][14] ) );
  dffascs1 \IDinst/RegFile_reg[2][14]  ( .DIN(\IDinst/n5450 ), .CLK(clk), 
        .CLRB(n865), .SETB(1'b1), .Q(\IDinst/RegFile[2][14] ) );
  dffascs1 \IDinst/RegFile_reg[3][14]  ( .DIN(\IDinst/n5449 ), .CLK(clk), 
        .CLRB(n865), .SETB(1'b1), .Q(\IDinst/RegFile[3][14] ) );
  dffascs1 \IDinst/RegFile_reg[4][14]  ( .DIN(\IDinst/n5448 ), .CLK(clk), 
        .CLRB(n865), .SETB(1'b1), .Q(\IDinst/RegFile[4][14] ) );
  dffascs1 \IDinst/RegFile_reg[5][14]  ( .DIN(\IDinst/n5447 ), .CLK(clk), 
        .CLRB(n865), .SETB(1'b1), .Q(\IDinst/RegFile[5][14] ) );
  dffascs1 \IDinst/RegFile_reg[6][14]  ( .DIN(\IDinst/n5446 ), .CLK(clk), 
        .CLRB(n865), .SETB(1'b1), .Q(\IDinst/RegFile[6][14] ) );
  dffascs1 \IDinst/RegFile_reg[7][14]  ( .DIN(\IDinst/n5445 ), .CLK(clk), 
        .CLRB(n865), .SETB(1'b1), .Q(\IDinst/RegFile[7][14] ) );
  dffascs1 \IDinst/RegFile_reg[8][14]  ( .DIN(\IDinst/n5444 ), .CLK(clk), 
        .CLRB(n865), .SETB(1'b1), .Q(\IDinst/RegFile[8][14] ) );
  dffascs1 \IDinst/RegFile_reg[9][14]  ( .DIN(\IDinst/n5443 ), .CLK(clk), 
        .CLRB(n865), .SETB(1'b1), .Q(\IDinst/RegFile[9][14] ) );
  dffascs1 \IDinst/RegFile_reg[10][14]  ( .DIN(\IDinst/n5442 ), .CLK(clk), 
        .CLRB(n865), .SETB(1'b1), .Q(\IDinst/RegFile[10][14] ) );
  dffascs1 \IDinst/RegFile_reg[11][14]  ( .DIN(\IDinst/n5441 ), .CLK(clk), 
        .CLRB(n865), .SETB(1'b1), .Q(\IDinst/RegFile[11][14] ) );
  dffascs1 \IDinst/RegFile_reg[12][14]  ( .DIN(\IDinst/n5440 ), .CLK(clk), 
        .CLRB(n866), .SETB(1'b1), .Q(\IDinst/RegFile[12][14] ) );
  dffascs1 \IDinst/RegFile_reg[13][14]  ( .DIN(\IDinst/n5439 ), .CLK(clk), 
        .CLRB(n866), .SETB(1'b1), .Q(\IDinst/RegFile[13][14] ) );
  dffascs1 \IDinst/RegFile_reg[14][14]  ( .DIN(\IDinst/n5438 ), .CLK(clk), 
        .CLRB(n866), .SETB(1'b1), .Q(\IDinst/RegFile[14][14] ) );
  dffascs1 \IDinst/RegFile_reg[15][14]  ( .DIN(\IDinst/n5437 ), .CLK(clk), 
        .CLRB(n866), .SETB(1'b1), .Q(\IDinst/RegFile[15][14] ) );
  dffascs1 \IDinst/RegFile_reg[16][14]  ( .DIN(\IDinst/n5436 ), .CLK(clk), 
        .CLRB(n866), .SETB(1'b1), .Q(\IDinst/RegFile[16][14] ) );
  dffascs1 \IDinst/RegFile_reg[17][14]  ( .DIN(\IDinst/n5435 ), .CLK(clk), 
        .CLRB(n866), .SETB(1'b1), .Q(\IDinst/RegFile[17][14] ) );
  dffascs1 \IDinst/RegFile_reg[18][14]  ( .DIN(\IDinst/n5434 ), .CLK(clk), 
        .CLRB(n866), .SETB(1'b1), .Q(\IDinst/RegFile[18][14] ) );
  dffascs1 \IDinst/RegFile_reg[19][14]  ( .DIN(\IDinst/n5433 ), .CLK(clk), 
        .CLRB(n866), .SETB(1'b1), .Q(\IDinst/RegFile[19][14] ) );
  dffascs1 \IDinst/RegFile_reg[20][14]  ( .DIN(\IDinst/n5432 ), .CLK(clk), 
        .CLRB(n866), .SETB(1'b1), .Q(\IDinst/RegFile[20][14] ) );
  dffascs1 \IDinst/RegFile_reg[21][14]  ( .DIN(\IDinst/n5431 ), .CLK(clk), 
        .CLRB(n866), .SETB(1'b1), .Q(\IDinst/RegFile[21][14] ) );
  dffascs1 \IDinst/RegFile_reg[22][14]  ( .DIN(\IDinst/n5430 ), .CLK(clk), 
        .CLRB(n867), .SETB(1'b1), .Q(\IDinst/RegFile[22][14] ) );
  dffascs1 \IDinst/RegFile_reg[23][14]  ( .DIN(\IDinst/n5429 ), .CLK(clk), 
        .CLRB(n867), .SETB(1'b1), .Q(\IDinst/RegFile[23][14] ) );
  dffascs1 \IDinst/RegFile_reg[24][14]  ( .DIN(\IDinst/n5428 ), .CLK(clk), 
        .CLRB(n867), .SETB(1'b1), .Q(\IDinst/RegFile[24][14] ) );
  dffascs1 \IDinst/RegFile_reg[25][14]  ( .DIN(\IDinst/n5427 ), .CLK(clk), 
        .CLRB(n867), .SETB(1'b1), .Q(\IDinst/RegFile[25][14] ) );
  dffascs1 \IDinst/RegFile_reg[26][14]  ( .DIN(\IDinst/n5426 ), .CLK(clk), 
        .CLRB(n867), .SETB(1'b1), .Q(\IDinst/RegFile[26][14] ) );
  dffascs1 \IDinst/RegFile_reg[27][14]  ( .DIN(\IDinst/n5425 ), .CLK(clk), 
        .CLRB(n867), .SETB(1'b1), .Q(\IDinst/RegFile[27][14] ) );
  dffascs1 \IDinst/RegFile_reg[28][14]  ( .DIN(\IDinst/n5424 ), .CLK(clk), 
        .CLRB(n867), .SETB(1'b1), .Q(\IDinst/RegFile[28][14] ) );
  dffascs1 \IDinst/RegFile_reg[29][14]  ( .DIN(\IDinst/n5423 ), .CLK(clk), 
        .CLRB(n867), .SETB(1'b1), .Q(\IDinst/RegFile[29][14] ) );
  dffascs1 \IDinst/RegFile_reg[30][14]  ( .DIN(\IDinst/n5422 ), .CLK(clk), 
        .CLRB(n867), .SETB(1'b1), .Q(\IDinst/RegFile[30][14] ) );
  dffascs1 \IDinst/RegFile_reg[31][14]  ( .DIN(\IDinst/n5421 ), .CLK(clk), 
        .CLRB(n867), .SETB(1'b1), .Q(\IDinst/RegFile[31][14] ) );
  dffascs1 \IDinst/opcode_of_WB_reg[0]  ( .DIN(\IDinst/opcode_of_MEM[0]), 
        .CLK(clk), .CLRB(n939), .SETB(1'b1), .QN(n9405) );
  dffascs1 \IDinst/opcode_of_MEM_reg[0]  ( .DIN(IR_opcode_field[0]), .CLK(clk), 
        .CLRB(n939), .SETB(1'b1), .Q(\IDinst/opcode_of_MEM[0]) );
  dffascs1 \IDinst/IR_opcode_field_reg[0]  ( .DIN(\IDinst/n5650 ), .CLK(clk), 
        .CLRB(n940), .SETB(1'b1), .Q(IR_opcode_field[0]), .QN(n132) );
  dffascs1 \IDinst/opcode_of_WB_reg[1]  ( .DIN(\IDinst/opcode_of_MEM[1]), 
        .CLK(clk), .CLRB(n940), .SETB(1'b1), .QN(n9403) );
  dffascs1 \IDinst/opcode_of_MEM_reg[1]  ( .DIN(IR_opcode_field[1]), .CLK(clk), 
        .CLRB(n940), .SETB(1'b1), .Q(\IDinst/opcode_of_MEM[1]), .QN(n225) );
  dffascs1 \IDinst/IR_opcode_field_reg[1]  ( .DIN(\IDinst/n5649 ), .CLK(clk), 
        .CLRB(n940), .SETB(1'b1), .Q(IR_opcode_field[1]), .QN(n40) );
  dffascs1 \IDinst/opcode_of_WB_reg[2]  ( .DIN(\IDinst/opcode_of_MEM[2]), 
        .CLK(clk), .CLRB(n940), .SETB(1'b1), .Q(\IDinst/opcode_of_WB[2] ), 
        .QN(n379) );
  dffascs1 \IDinst/opcode_of_MEM_reg[2]  ( .DIN(IR_opcode_field[2]), .CLK(clk), 
        .CLRB(n940), .SETB(1'b1), .Q(\IDinst/opcode_of_MEM[2]), .QN(n209) );
  dffascs1 \IDinst/IR_opcode_field_reg[2]  ( .DIN(\IDinst/n5648 ), .CLK(clk), 
        .CLRB(n941), .SETB(1'b1), .Q(IR_opcode_field[2]), .QN(n39) );
  dffascs1 \IDinst/opcode_of_WB_reg[3]  ( .DIN(\IDinst/opcode_of_MEM[3]), 
        .CLK(clk), .CLRB(n941), .SETB(1'b1), .QN(n9400) );
  dffascs1 \IDinst/opcode_of_MEM_reg[3]  ( .DIN(IR_opcode_field[3]), .CLK(clk), 
        .CLRB(n941), .SETB(1'b1), .Q(\IDinst/opcode_of_MEM[3]), .QN(n375) );
  dffascs1 \IDinst/IR_opcode_field_reg[3]  ( .DIN(\IDinst/n5647 ), .CLK(clk), 
        .CLRB(n941), .SETB(1'b1), .Q(IR_opcode_field[3]), .QN(n760) );
  dffascs1 \IDinst/opcode_of_WB_reg[4]  ( .DIN(\IDinst/opcode_of_MEM[4]), 
        .CLK(clk), .CLRB(n926), .SETB(1'b1), .QN(n9401) );
  dffascs1 \IDinst/opcode_of_MEM_reg[4]  ( .DIN(IR_opcode_field[4]), .CLK(clk), 
        .CLRB(n950), .SETB(1'b1), .Q(\IDinst/opcode_of_MEM[4]), .QN(n59) );
  dffascs1 \IDinst/IR_opcode_field_reg[4]  ( .DIN(\IDinst/n5646 ), .CLK(clk), 
        .CLRB(n950), .SETB(1'b1), .Q(IR_opcode_field[4]), .QN(n101) );
  dffascs1 \IDinst/opcode_of_WB_reg[5]  ( .DIN(\IDinst/opcode_of_MEM[5]), 
        .CLK(clk), .CLRB(n925), .SETB(1'b1), .Q(n9402) );
  dffascs1 \IDinst/opcode_of_MEM_reg[5]  ( .DIN(IR_opcode_field[5]), .CLK(clk), 
        .CLRB(n958), .SETB(1'b1), .Q(\IDinst/opcode_of_MEM[5]), .QN(n57) );
  dffascs1 \IDinst/IR_opcode_field_reg[5]  ( .DIN(\IDinst/n5645 ), .CLK(clk), 
        .CLRB(n958), .SETB(1'b1), .Q(IR_opcode_field[5]), .QN(n117) );
  dffascs1 \IDinst/IR_function_field_reg[0]  ( .DIN(\IDinst/n4876 ), .CLK(clk), 
        .CLRB(n1019), .SETB(1'b1), .Q(n19), .QN(n9458) );
  dffascs1 \IDinst/IR_function_field_reg[1]  ( .DIN(\IDinst/n4875 ), .CLK(clk), 
        .CLRB(n941), .SETB(1'b1), .Q(n2) );
  dffascs1 \IDinst/IR_function_field_reg[2]  ( .DIN(\IDinst/n4874 ), .CLK(clk), 
        .CLRB(n941), .SETB(1'b1), .Q(n17), .QN(n9457) );
  dffascs1 \IDinst/IR_function_field_reg[3]  ( .DIN(\IDinst/n4873 ), .CLK(clk), 
        .CLRB(n941), .SETB(1'b1), .Q(n137), .QN(n9456) );
  dffascs1 \IDinst/IR_function_field_reg[4]  ( .DIN(\IDinst/n4872 ), .CLK(clk), 
        .CLRB(n941), .SETB(1'b1), .QN(n9416) );
  dffascs1 \IDinst/mem_to_reg_reg  ( .DIN(\IDinst/n4866 ), .CLK(clk), 
        .CLRB(n941), .SETB(1'b1), .QN(n9413) );
  dffascs1 \IDinst/rt_addr_reg[0]  ( .DIN(\IDinst/n4865 ), .CLK(clk), 
        .CLRB(n942), .SETB(1'b1), .Q(n229), .QN(n9407) );
  dffascs1 \IDinst/RegFile_reg[25][7]  ( .DIN(\IDinst/n5851 ), .CLK(clk), 
        .CLRB(n850), .SETB(1'b1), .Q(\IDinst/RegFile[25][7] ) );
  dffascs1 \IDinst/RegFile_reg[25][6]  ( .DIN(\IDinst/n5852 ), .CLK(clk), 
        .CLRB(n846), .SETB(1'b1), .Q(\IDinst/RegFile[25][6] ) );
  dffascs1 \IDinst/RegFile_reg[25][5]  ( .DIN(\IDinst/n5853 ), .CLK(clk), 
        .CLRB(n853), .SETB(1'b1), .Q(\IDinst/RegFile[25][5] ) );
  dffascs1 \IDinst/RegFile_reg[25][4]  ( .DIN(\IDinst/n5854 ), .CLK(clk), 
        .CLRB(n869), .SETB(1'b1), .Q(\IDinst/RegFile[25][4] ) );
  dffascs1 \IDinst/RegFile_reg[25][3]  ( .DIN(\IDinst/n5855 ), .CLK(clk), 
        .CLRB(n841), .SETB(1'b1), .Q(\IDinst/RegFile[25][3] ) );
  dffascs1 \IDinst/RegFile_reg[25][2]  ( .DIN(\IDinst/n5856 ), .CLK(clk), 
        .CLRB(n838), .SETB(1'b1), .Q(\IDinst/RegFile[25][2] ) );
  dffascs1 \IDinst/RegFile_reg[25][1]  ( .DIN(\IDinst/n5857 ), .CLK(clk), 
        .CLRB(n834), .SETB(1'b1), .Q(\IDinst/RegFile[25][1] ) );
  dffascs1 \IDinst/RegFile_reg[25][0]  ( .DIN(\IDinst/n5858 ), .CLK(clk), 
        .CLRB(n927), .SETB(1'b1), .Q(\IDinst/RegFile[25][0] ) );
  dffascs1 \IDinst/RegFile_reg[17][7]  ( .DIN(\IDinst/n5787 ), .CLK(clk), 
        .CLRB(n850), .SETB(1'b1), .Q(\IDinst/RegFile[17][7] ) );
  dffascs1 \IDinst/RegFile_reg[17][6]  ( .DIN(\IDinst/n5788 ), .CLK(clk), 
        .CLRB(n847), .SETB(1'b1), .Q(\IDinst/RegFile[17][6] ) );
  dffascs1 \IDinst/RegFile_reg[17][5]  ( .DIN(\IDinst/n5789 ), .CLK(clk), 
        .CLRB(n854), .SETB(1'b1), .Q(\IDinst/RegFile[17][5] ) );
  dffascs1 \IDinst/RegFile_reg[17][4]  ( .DIN(\IDinst/n5790 ), .CLK(clk), 
        .CLRB(n869), .SETB(1'b1), .Q(\IDinst/RegFile[17][4] ) );
  dffascs1 \IDinst/RegFile_reg[17][3]  ( .DIN(\IDinst/n5791 ), .CLK(clk), 
        .CLRB(n842), .SETB(1'b1), .Q(\IDinst/RegFile[17][3] ) );
  dffascs1 \IDinst/RegFile_reg[17][2]  ( .DIN(\IDinst/n5792 ), .CLK(clk), 
        .CLRB(n839), .SETB(1'b1), .Q(\IDinst/RegFile[17][2] ) );
  dffascs1 \IDinst/RegFile_reg[17][1]  ( .DIN(\IDinst/n5793 ), .CLK(clk), 
        .CLRB(n835), .SETB(1'b1), .Q(\IDinst/RegFile[17][1] ) );
  dffascs1 \IDinst/RegFile_reg[17][0]  ( .DIN(\IDinst/n5794 ), .CLK(clk), 
        .CLRB(n930), .SETB(1'b1), .Q(\IDinst/RegFile[17][0] ) );
  dffascs1 \IDinst/RegFile_reg[9][7]  ( .DIN(\IDinst/n5723 ), .CLK(clk), 
        .CLRB(n851), .SETB(1'b1), .Q(\IDinst/RegFile[9][7] ) );
  dffascs1 \IDinst/RegFile_reg[9][6]  ( .DIN(\IDinst/n5724 ), .CLK(clk), 
        .CLRB(n847), .SETB(1'b1), .Q(\IDinst/RegFile[9][6] ) );
  dffascs1 \IDinst/RegFile_reg[9][5]  ( .DIN(\IDinst/n5725 ), .CLK(clk), 
        .CLRB(n855), .SETB(1'b1), .Q(\IDinst/RegFile[9][5] ) );
  dffascs1 \IDinst/RegFile_reg[9][4]  ( .DIN(\IDinst/n5726 ), .CLK(clk), 
        .CLRB(n870), .SETB(1'b1), .Q(\IDinst/RegFile[9][4] ) );
  dffascs1 \IDinst/RegFile_reg[9][3]  ( .DIN(\IDinst/n5727 ), .CLK(clk), 
        .CLRB(n843), .SETB(1'b1), .Q(\IDinst/RegFile[9][3] ) );
  dffascs1 \IDinst/RegFile_reg[9][2]  ( .DIN(\IDinst/n5728 ), .CLK(clk), 
        .CLRB(n839), .SETB(1'b1), .Q(\IDinst/RegFile[9][2] ) );
  dffascs1 \IDinst/RegFile_reg[9][1]  ( .DIN(\IDinst/n5729 ), .CLK(clk), 
        .CLRB(n836), .SETB(1'b1), .Q(\IDinst/RegFile[9][1] ) );
  dffascs1 \IDinst/RegFile_reg[9][0]  ( .DIN(\IDinst/n5730 ), .CLK(clk), 
        .CLRB(n933), .SETB(1'b1), .Q(\IDinst/RegFile[9][0] ) );
  dffascs1 \IDinst/RegFile_reg[1][7]  ( .DIN(\IDinst/n5659 ), .CLK(clk), 
        .CLRB(n852), .SETB(1'b1), .Q(\IDinst/RegFile[1][7] ) );
  dffascs1 \IDinst/RegFile_reg[1][6]  ( .DIN(\IDinst/n5660 ), .CLK(clk), 
        .CLRB(n848), .SETB(1'b1), .Q(\IDinst/RegFile[1][6] ) );
  dffascs1 \IDinst/RegFile_reg[1][5]  ( .DIN(\IDinst/n5661 ), .CLK(clk), 
        .CLRB(n856), .SETB(1'b1), .Q(\IDinst/RegFile[1][5] ) );
  dffascs1 \IDinst/RegFile_reg[1][4]  ( .DIN(\IDinst/n5662 ), .CLK(clk), 
        .CLRB(n871), .SETB(1'b1), .Q(\IDinst/RegFile[1][4] ) );
  dffascs1 \IDinst/RegFile_reg[1][3]  ( .DIN(\IDinst/n5663 ), .CLK(clk), 
        .CLRB(n844), .SETB(1'b1), .Q(\IDinst/RegFile[1][3] ) );
  dffascs1 \IDinst/RegFile_reg[1][2]  ( .DIN(\IDinst/n5664 ), .CLK(clk), 
        .CLRB(n840), .SETB(1'b1), .Q(\IDinst/RegFile[1][2] ) );
  dffascs1 \IDinst/RegFile_reg[1][1]  ( .DIN(\IDinst/n5665 ), .CLK(clk), 
        .CLRB(n837), .SETB(1'b1), .Q(\IDinst/RegFile[1][1] ) );
  dffascs1 \IDinst/RegFile_reg[1][0]  ( .DIN(\IDinst/n5666 ), .CLK(clk), 
        .CLRB(n936), .SETB(1'b1), .Q(\IDinst/RegFile[1][0] ) );
  dffascs1 \IDinst/RegFile_reg[28][7]  ( .DIN(\IDinst/n5875 ), .CLK(clk), 
        .CLRB(n849), .SETB(1'b1), .Q(\IDinst/RegFile[28][7] ) );
  dffascs1 \IDinst/RegFile_reg[28][6]  ( .DIN(\IDinst/n5876 ), .CLK(clk), 
        .CLRB(n846), .SETB(1'b1), .Q(\IDinst/RegFile[28][6] ) );
  dffascs1 \IDinst/RegFile_reg[28][5]  ( .DIN(\IDinst/n5877 ), .CLK(clk), 
        .CLRB(n853), .SETB(1'b1), .Q(\IDinst/RegFile[28][5] ) );
  dffascs1 \IDinst/RegFile_reg[28][4]  ( .DIN(\IDinst/n5878 ), .CLK(clk), 
        .CLRB(n868), .SETB(1'b1), .Q(\IDinst/RegFile[28][4] ) );
  dffascs1 \IDinst/RegFile_reg[28][3]  ( .DIN(\IDinst/n5879 ), .CLK(clk), 
        .CLRB(n841), .SETB(1'b1), .Q(\IDinst/RegFile[28][3] ) );
  dffascs1 \IDinst/RegFile_reg[28][2]  ( .DIN(\IDinst/n5880 ), .CLK(clk), 
        .CLRB(n838), .SETB(1'b1), .Q(\IDinst/RegFile[28][2] ) );
  dffascs1 \IDinst/RegFile_reg[28][1]  ( .DIN(\IDinst/n5881 ), .CLK(clk), 
        .CLRB(n834), .SETB(1'b1), .Q(\IDinst/RegFile[28][1] ) );
  dffascs1 \IDinst/RegFile_reg[28][0]  ( .DIN(\IDinst/n5882 ), .CLK(clk), 
        .CLRB(n928), .SETB(1'b1), .Q(\IDinst/RegFile[28][0] ) );
  dffascs1 \IDinst/RegFile_reg[20][7]  ( .DIN(\IDinst/n5811 ), .CLK(clk), 
        .CLRB(n850), .SETB(1'b1), .Q(\IDinst/RegFile[20][7] ) );
  dffascs1 \IDinst/RegFile_reg[20][6]  ( .DIN(\IDinst/n5812 ), .CLK(clk), 
        .CLRB(n846), .SETB(1'b1), .Q(\IDinst/RegFile[20][6] ) );
  dffascs1 \IDinst/RegFile_reg[20][5]  ( .DIN(\IDinst/n5813 ), .CLK(clk), 
        .CLRB(n854), .SETB(1'b1), .Q(\IDinst/RegFile[20][5] ) );
  dffascs1 \IDinst/RegFile_reg[20][4]  ( .DIN(\IDinst/n5814 ), .CLK(clk), 
        .CLRB(n869), .SETB(1'b1), .Q(\IDinst/RegFile[20][4] ) );
  dffascs1 \IDinst/RegFile_reg[20][3]  ( .DIN(\IDinst/n5815 ), .CLK(clk), 
        .CLRB(n842), .SETB(1'b1), .Q(\IDinst/RegFile[20][3] ) );
  dffascs1 \IDinst/RegFile_reg[20][2]  ( .DIN(\IDinst/n5816 ), .CLK(clk), 
        .CLRB(n838), .SETB(1'b1), .Q(\IDinst/RegFile[20][2] ) );
  dffascs1 \IDinst/RegFile_reg[20][1]  ( .DIN(\IDinst/n5817 ), .CLK(clk), 
        .CLRB(n835), .SETB(1'b1), .Q(\IDinst/RegFile[20][1] ) );
  dffascs1 \IDinst/RegFile_reg[20][0]  ( .DIN(\IDinst/n5818 ), .CLK(clk), 
        .CLRB(n931), .SETB(1'b1), .Q(\IDinst/RegFile[20][0] ) );
  dffascs1 \IDinst/RegFile_reg[12][7]  ( .DIN(\IDinst/n5747 ), .CLK(clk), 
        .CLRB(n851), .SETB(1'b1), .Q(\IDinst/RegFile[12][7] ) );
  dffascs1 \IDinst/RegFile_reg[12][6]  ( .DIN(\IDinst/n5748 ), .CLK(clk), 
        .CLRB(n847), .SETB(1'b1), .Q(\IDinst/RegFile[12][6] ) );
  dffascs1 \IDinst/RegFile_reg[12][5]  ( .DIN(\IDinst/n5749 ), .CLK(clk), 
        .CLRB(n855), .SETB(1'b1), .Q(\IDinst/RegFile[12][5] ) );
  dffascs1 \IDinst/RegFile_reg[12][4]  ( .DIN(\IDinst/n5750 ), .CLK(clk), 
        .CLRB(n870), .SETB(1'b1), .Q(\IDinst/RegFile[12][4] ) );
  dffascs1 \IDinst/RegFile_reg[12][3]  ( .DIN(\IDinst/n5751 ), .CLK(clk), 
        .CLRB(n843), .SETB(1'b1), .Q(\IDinst/RegFile[12][3] ) );
  dffascs1 \IDinst/RegFile_reg[12][2]  ( .DIN(\IDinst/n5752 ), .CLK(clk), 
        .CLRB(n839), .SETB(1'b1), .Q(\IDinst/RegFile[12][2] ) );
  dffascs1 \IDinst/RegFile_reg[12][1]  ( .DIN(\IDinst/n5753 ), .CLK(clk), 
        .CLRB(n836), .SETB(1'b1), .Q(\IDinst/RegFile[12][1] ) );
  dffascs1 \IDinst/RegFile_reg[12][0]  ( .DIN(\IDinst/n5754 ), .CLK(clk), 
        .CLRB(n934), .SETB(1'b1), .Q(\IDinst/RegFile[12][0] ) );
  dffascs1 \IDinst/RegFile_reg[4][7]  ( .DIN(\IDinst/n5683 ), .CLK(clk), 
        .CLRB(n852), .SETB(1'b1), .Q(\IDinst/RegFile[4][7] ) );
  dffascs1 \IDinst/RegFile_reg[4][6]  ( .DIN(\IDinst/n5684 ), .CLK(clk), 
        .CLRB(n848), .SETB(1'b1), .Q(\IDinst/RegFile[4][6] ) );
  dffascs1 \IDinst/RegFile_reg[4][5]  ( .DIN(\IDinst/n5685 ), .CLK(clk), 
        .CLRB(n855), .SETB(1'b1), .Q(\IDinst/RegFile[4][5] ) );
  dffascs1 \IDinst/RegFile_reg[4][4]  ( .DIN(\IDinst/n5686 ), .CLK(clk), 
        .CLRB(n871), .SETB(1'b1), .Q(\IDinst/RegFile[4][4] ) );
  dffascs1 \IDinst/RegFile_reg[4][3]  ( .DIN(\IDinst/n5687 ), .CLK(clk), 
        .CLRB(n844), .SETB(1'b1), .Q(\IDinst/RegFile[4][3] ) );
  dffascs1 \IDinst/RegFile_reg[4][2]  ( .DIN(\IDinst/n5688 ), .CLK(clk), 
        .CLRB(n840), .SETB(1'b1), .Q(\IDinst/RegFile[4][2] ) );
  dffascs1 \IDinst/RegFile_reg[4][1]  ( .DIN(\IDinst/n5689 ), .CLK(clk), 
        .CLRB(n836), .SETB(1'b1), .Q(\IDinst/RegFile[4][1] ) );
  dffascs1 \IDinst/RegFile_reg[4][0]  ( .DIN(\IDinst/n5690 ), .CLK(clk), 
        .CLRB(n937), .SETB(1'b1), .Q(\IDinst/RegFile[4][0] ) );
  dffascs1 \IDinst/RegFile_reg[29][7]  ( .DIN(\IDinst/n5883 ), .CLK(clk), 
        .CLRB(n849), .SETB(1'b1), .Q(\IDinst/RegFile[29][7] ) );
  dffascs1 \IDinst/RegFile_reg[29][6]  ( .DIN(\IDinst/n5884 ), .CLK(clk), 
        .CLRB(n845), .SETB(1'b1), .Q(\IDinst/RegFile[29][6] ) );
  dffascs1 \IDinst/RegFile_reg[29][5]  ( .DIN(\IDinst/n5885 ), .CLK(clk), 
        .CLRB(n853), .SETB(1'b1), .Q(\IDinst/RegFile[29][5] ) );
  dffascs1 \IDinst/RegFile_reg[29][4]  ( .DIN(\IDinst/n5886 ), .CLK(clk), 
        .CLRB(n868), .SETB(1'b1), .Q(\IDinst/RegFile[29][4] ) );
  dffascs1 \IDinst/RegFile_reg[29][3]  ( .DIN(\IDinst/n5887 ), .CLK(clk), 
        .CLRB(n841), .SETB(1'b1), .Q(\IDinst/RegFile[29][3] ) );
  dffascs1 \IDinst/RegFile_reg[29][2]  ( .DIN(\IDinst/n5888 ), .CLK(clk), 
        .CLRB(n837), .SETB(1'b1), .Q(\IDinst/RegFile[29][2] ) );
  dffascs1 \IDinst/RegFile_reg[29][1]  ( .DIN(\IDinst/n5889 ), .CLK(clk), 
        .CLRB(n834), .SETB(1'b1), .Q(\IDinst/RegFile[29][1] ) );
  dffascs1 \IDinst/RegFile_reg[29][0]  ( .DIN(\IDinst/n5890 ), .CLK(clk), 
        .CLRB(n929), .SETB(1'b1), .Q(\IDinst/RegFile[29][0] ) );
  dffascs1 \IDinst/RegFile_reg[21][7]  ( .DIN(\IDinst/n5819 ), .CLK(clk), 
        .CLRB(n850), .SETB(1'b1), .Q(\IDinst/RegFile[21][7] ) );
  dffascs1 \IDinst/RegFile_reg[21][6]  ( .DIN(\IDinst/n5820 ), .CLK(clk), 
        .CLRB(n846), .SETB(1'b1), .Q(\IDinst/RegFile[21][6] ) );
  dffascs1 \IDinst/RegFile_reg[21][5]  ( .DIN(\IDinst/n5821 ), .CLK(clk), 
        .CLRB(n854), .SETB(1'b1), .Q(\IDinst/RegFile[21][5] ) );
  dffascs1 \IDinst/RegFile_reg[21][4]  ( .DIN(\IDinst/n5822 ), .CLK(clk), 
        .CLRB(n869), .SETB(1'b1), .Q(\IDinst/RegFile[21][4] ) );
  dffascs1 \IDinst/RegFile_reg[21][3]  ( .DIN(\IDinst/n5823 ), .CLK(clk), 
        .CLRB(n842), .SETB(1'b1), .Q(\IDinst/RegFile[21][3] ) );
  dffascs1 \IDinst/RegFile_reg[21][2]  ( .DIN(\IDinst/n5824 ), .CLK(clk), 
        .CLRB(n838), .SETB(1'b1), .Q(\IDinst/RegFile[21][2] ) );
  dffascs1 \IDinst/RegFile_reg[21][1]  ( .DIN(\IDinst/n5825 ), .CLK(clk), 
        .CLRB(n835), .SETB(1'b1), .Q(\IDinst/RegFile[21][1] ) );
  dffascs1 \IDinst/RegFile_reg[21][0]  ( .DIN(\IDinst/n5826 ), .CLK(clk), 
        .CLRB(n932), .SETB(1'b1), .Q(\IDinst/RegFile[21][0] ) );
  dffascs1 \IDinst/RegFile_reg[13][7]  ( .DIN(\IDinst/n5755 ), .CLK(clk), 
        .CLRB(n851), .SETB(1'b1), .Q(\IDinst/RegFile[13][7] ) );
  dffascs1 \IDinst/RegFile_reg[13][6]  ( .DIN(\IDinst/n5756 ), .CLK(clk), 
        .CLRB(n847), .SETB(1'b1), .Q(\IDinst/RegFile[13][6] ) );
  dffascs1 \IDinst/RegFile_reg[13][5]  ( .DIN(\IDinst/n5757 ), .CLK(clk), 
        .CLRB(n854), .SETB(1'b1), .Q(\IDinst/RegFile[13][5] ) );
  dffascs1 \IDinst/RegFile_reg[13][4]  ( .DIN(\IDinst/n5758 ), .CLK(clk), 
        .CLRB(n870), .SETB(1'b1), .Q(\IDinst/RegFile[13][4] ) );
  dffascs1 \IDinst/RegFile_reg[13][3]  ( .DIN(\IDinst/n5759 ), .CLK(clk), 
        .CLRB(n843), .SETB(1'b1), .Q(\IDinst/RegFile[13][3] ) );
  dffascs1 \IDinst/RegFile_reg[13][2]  ( .DIN(\IDinst/n5760 ), .CLK(clk), 
        .CLRB(n839), .SETB(1'b1), .Q(\IDinst/RegFile[13][2] ) );
  dffascs1 \IDinst/RegFile_reg[13][1]  ( .DIN(\IDinst/n5761 ), .CLK(clk), 
        .CLRB(n835), .SETB(1'b1), .Q(\IDinst/RegFile[13][1] ) );
  dffascs1 \IDinst/RegFile_reg[13][0]  ( .DIN(\IDinst/n5762 ), .CLK(clk), 
        .CLRB(n935), .SETB(1'b1), .Q(\IDinst/RegFile[13][0] ) );
  dffascs1 \IDinst/RegFile_reg[5][7]  ( .DIN(\IDinst/n5691 ), .CLK(clk), 
        .CLRB(n852), .SETB(1'b1), .Q(\IDinst/RegFile[5][7] ) );
  dffascs1 \IDinst/RegFile_reg[5][6]  ( .DIN(\IDinst/n5692 ), .CLK(clk), 
        .CLRB(n848), .SETB(1'b1), .Q(\IDinst/RegFile[5][6] ) );
  dffascs1 \IDinst/RegFile_reg[5][5]  ( .DIN(\IDinst/n5693 ), .CLK(clk), 
        .CLRB(n855), .SETB(1'b1), .Q(\IDinst/RegFile[5][5] ) );
  dffascs1 \IDinst/RegFile_reg[5][4]  ( .DIN(\IDinst/n5694 ), .CLK(clk), 
        .CLRB(n871), .SETB(1'b1), .Q(\IDinst/RegFile[5][4] ) );
  dffascs1 \IDinst/RegFile_reg[5][3]  ( .DIN(\IDinst/n5695 ), .CLK(clk), 
        .CLRB(n843), .SETB(1'b1), .Q(\IDinst/RegFile[5][3] ) );
  dffascs1 \IDinst/RegFile_reg[5][2]  ( .DIN(\IDinst/n5696 ), .CLK(clk), 
        .CLRB(n840), .SETB(1'b1), .Q(\IDinst/RegFile[5][2] ) );
  dffascs1 \IDinst/RegFile_reg[5][1]  ( .DIN(\IDinst/n5697 ), .CLK(clk), 
        .CLRB(n836), .SETB(1'b1), .Q(\IDinst/RegFile[5][1] ) );
  dffascs1 \IDinst/RegFile_reg[5][0]  ( .DIN(\IDinst/n5698 ), .CLK(clk), 
        .CLRB(n938), .SETB(1'b1), .Q(\IDinst/RegFile[5][0] ) );
  dffascs1 \IDinst/RegFile_reg[24][7]  ( .DIN(\IDinst/n5843 ), .CLK(clk), 
        .CLRB(n850), .SETB(1'b1), .Q(\IDinst/RegFile[24][7] ) );
  dffascs1 \IDinst/RegFile_reg[24][6]  ( .DIN(\IDinst/n5844 ), .CLK(clk), 
        .CLRB(n846), .SETB(1'b1), .Q(\IDinst/RegFile[24][6] ) );
  dffascs1 \IDinst/RegFile_reg[24][5]  ( .DIN(\IDinst/n5845 ), .CLK(clk), 
        .CLRB(n853), .SETB(1'b1), .Q(\IDinst/RegFile[24][5] ) );
  dffascs1 \IDinst/RegFile_reg[24][4]  ( .DIN(\IDinst/n5846 ), .CLK(clk), 
        .CLRB(n869), .SETB(1'b1), .Q(\IDinst/RegFile[24][4] ) );
  dffascs1 \IDinst/RegFile_reg[24][3]  ( .DIN(\IDinst/n5847 ), .CLK(clk), 
        .CLRB(n842), .SETB(1'b1), .Q(\IDinst/RegFile[24][3] ) );
  dffascs1 \IDinst/RegFile_reg[24][2]  ( .DIN(\IDinst/n5848 ), .CLK(clk), 
        .CLRB(n838), .SETB(1'b1), .Q(\IDinst/RegFile[24][2] ) );
  dffascs1 \IDinst/RegFile_reg[24][1]  ( .DIN(\IDinst/n5849 ), .CLK(clk), 
        .CLRB(n834), .SETB(1'b1), .Q(\IDinst/RegFile[24][1] ) );
  dffascs1 \IDinst/RegFile_reg[24][0]  ( .DIN(\IDinst/n5850 ), .CLK(clk), 
        .CLRB(n927), .SETB(1'b1), .Q(\IDinst/RegFile[24][0] ) );
  dffascs1 \IDinst/RegFile_reg[16][7]  ( .DIN(\IDinst/n5779 ), .CLK(clk), 
        .CLRB(n851), .SETB(1'b1), .Q(\IDinst/RegFile[16][7] ) );
  dffascs1 \IDinst/RegFile_reg[16][6]  ( .DIN(\IDinst/n5780 ), .CLK(clk), 
        .CLRB(n847), .SETB(1'b1), .Q(\IDinst/RegFile[16][6] ) );
  dffascs1 \IDinst/RegFile_reg[16][5]  ( .DIN(\IDinst/n5781 ), .CLK(clk), 
        .CLRB(n854), .SETB(1'b1), .Q(\IDinst/RegFile[16][5] ) );
  dffascs1 \IDinst/RegFile_reg[16][4]  ( .DIN(\IDinst/n5782 ), .CLK(clk), 
        .CLRB(n869), .SETB(1'b1), .Q(\IDinst/RegFile[16][4] ) );
  dffascs1 \IDinst/RegFile_reg[16][3]  ( .DIN(\IDinst/n5783 ), .CLK(clk), 
        .CLRB(n842), .SETB(1'b1), .Q(\IDinst/RegFile[16][3] ) );
  dffascs1 \IDinst/RegFile_reg[16][2]  ( .DIN(\IDinst/n5784 ), .CLK(clk), 
        .CLRB(n839), .SETB(1'b1), .Q(\IDinst/RegFile[16][2] ) );
  dffascs1 \IDinst/RegFile_reg[16][1]  ( .DIN(\IDinst/n5785 ), .CLK(clk), 
        .CLRB(n835), .SETB(1'b1), .Q(\IDinst/RegFile[16][1] ) );
  dffascs1 \IDinst/RegFile_reg[16][0]  ( .DIN(\IDinst/n5786 ), .CLK(clk), 
        .CLRB(n930), .SETB(1'b1), .Q(\IDinst/RegFile[16][0] ) );
  dffascs1 \IDinst/RegFile_reg[8][7]  ( .DIN(\IDinst/n5715 ), .CLK(clk), 
        .CLRB(n851), .SETB(1'b1), .Q(\IDinst/RegFile[8][7] ) );
  dffascs1 \IDinst/RegFile_reg[8][6]  ( .DIN(\IDinst/n5716 ), .CLK(clk), 
        .CLRB(n848), .SETB(1'b1), .Q(\IDinst/RegFile[8][6] ) );
  dffascs1 \IDinst/RegFile_reg[8][5]  ( .DIN(\IDinst/n5717 ), .CLK(clk), 
        .CLRB(n855), .SETB(1'b1), .Q(\IDinst/RegFile[8][5] ) );
  dffascs1 \IDinst/RegFile_reg[8][4]  ( .DIN(\IDinst/n5718 ), .CLK(clk), 
        .CLRB(n870), .SETB(1'b1), .Q(\IDinst/RegFile[8][4] ) );
  dffascs1 \IDinst/RegFile_reg[8][3]  ( .DIN(\IDinst/n5719 ), .CLK(clk), 
        .CLRB(n843), .SETB(1'b1), .Q(\IDinst/RegFile[8][3] ) );
  dffascs1 \IDinst/RegFile_reg[8][2]  ( .DIN(\IDinst/n5720 ), .CLK(clk), 
        .CLRB(n840), .SETB(1'b1), .Q(\IDinst/RegFile[8][2] ) );
  dffascs1 \IDinst/RegFile_reg[8][1]  ( .DIN(\IDinst/n5721 ), .CLK(clk), 
        .CLRB(n836), .SETB(1'b1), .Q(\IDinst/RegFile[8][1] ) );
  dffascs1 \IDinst/RegFile_reg[8][0]  ( .DIN(\IDinst/n5722 ), .CLK(clk), 
        .CLRB(n933), .SETB(1'b1), .Q(\IDinst/RegFile[8][0] ) );
  dffascs1 \IDinst/RegFile_reg[0][7]  ( .DIN(\IDinst/n5651 ), .CLK(clk), 
        .CLRB(n852), .SETB(1'b1), .Q(\IDinst/RegFile[0][7] ) );
  dffascs1 \IDinst/RegFile_reg[0][6]  ( .DIN(\IDinst/n5652 ), .CLK(clk), 
        .CLRB(n848), .SETB(1'b1), .Q(\IDinst/RegFile[0][6] ) );
  dffascs1 \IDinst/RegFile_reg[0][5]  ( .DIN(\IDinst/n5653 ), .CLK(clk), 
        .CLRB(n856), .SETB(1'b1), .Q(\IDinst/RegFile[0][5] ) );
  dffascs1 \IDinst/RegFile_reg[0][4]  ( .DIN(\IDinst/n5654 ), .CLK(clk), 
        .CLRB(n871), .SETB(1'b1), .Q(\IDinst/RegFile[0][4] ) );
  dffascs1 \IDinst/RegFile_reg[0][3]  ( .DIN(\IDinst/n5655 ), .CLK(clk), 
        .CLRB(n844), .SETB(1'b1), .Q(\IDinst/RegFile[0][3] ) );
  dffascs1 \IDinst/RegFile_reg[0][2]  ( .DIN(\IDinst/n5656 ), .CLK(clk), 
        .CLRB(n840), .SETB(1'b1), .Q(\IDinst/RegFile[0][2] ) );
  dffascs1 \IDinst/RegFile_reg[0][1]  ( .DIN(\IDinst/n5657 ), .CLK(clk), 
        .CLRB(n837), .SETB(1'b1), .Q(\IDinst/RegFile[0][1] ) );
  dffascs1 \IDinst/RegFile_reg[0][0]  ( .DIN(\IDinst/n5658 ), .CLK(clk), 
        .CLRB(n936), .SETB(1'b1), .Q(\IDinst/RegFile[0][0] ) );
  dffascs1 \IDinst/RegFile_reg[26][7]  ( .DIN(\IDinst/n5859 ), .CLK(clk), 
        .CLRB(n850), .SETB(1'b1), .Q(\IDinst/RegFile[26][7] ) );
  dffascs1 \IDinst/RegFile_reg[26][6]  ( .DIN(\IDinst/n5860 ), .CLK(clk), 
        .CLRB(n846), .SETB(1'b1), .Q(\IDinst/RegFile[26][6] ) );
  dffascs1 \IDinst/RegFile_reg[26][5]  ( .DIN(\IDinst/n5861 ), .CLK(clk), 
        .CLRB(n853), .SETB(1'b1), .Q(\IDinst/RegFile[26][5] ) );
  dffascs1 \IDinst/RegFile_reg[26][4]  ( .DIN(\IDinst/n5862 ), .CLK(clk), 
        .CLRB(n868), .SETB(1'b1), .Q(\IDinst/RegFile[26][4] ) );
  dffascs1 \IDinst/RegFile_reg[26][3]  ( .DIN(\IDinst/n5863 ), .CLK(clk), 
        .CLRB(n841), .SETB(1'b1), .Q(\IDinst/RegFile[26][3] ) );
  dffascs1 \IDinst/RegFile_reg[26][2]  ( .DIN(\IDinst/n5864 ), .CLK(clk), 
        .CLRB(n838), .SETB(1'b1), .Q(\IDinst/RegFile[26][2] ) );
  dffascs1 \IDinst/RegFile_reg[26][1]  ( .DIN(\IDinst/n5865 ), .CLK(clk), 
        .CLRB(n834), .SETB(1'b1), .Q(\IDinst/RegFile[26][1] ) );
  dffascs1 \IDinst/RegFile_reg[26][0]  ( .DIN(\IDinst/n5866 ), .CLK(clk), 
        .CLRB(n927), .SETB(1'b1), .Q(\IDinst/RegFile[26][0] ) );
  dffascs1 \IDinst/RegFile_reg[18][7]  ( .DIN(\IDinst/n5795 ), .CLK(clk), 
        .CLRB(n850), .SETB(1'b1), .Q(\IDinst/RegFile[18][7] ) );
  dffascs1 \IDinst/RegFile_reg[18][6]  ( .DIN(\IDinst/n5796 ), .CLK(clk), 
        .CLRB(n847), .SETB(1'b1), .Q(\IDinst/RegFile[18][6] ) );
  dffascs1 \IDinst/RegFile_reg[18][5]  ( .DIN(\IDinst/n5797 ), .CLK(clk), 
        .CLRB(n854), .SETB(1'b1), .Q(\IDinst/RegFile[18][5] ) );
  dffascs1 \IDinst/RegFile_reg[18][4]  ( .DIN(\IDinst/n5798 ), .CLK(clk), 
        .CLRB(n869), .SETB(1'b1), .Q(\IDinst/RegFile[18][4] ) );
  dffascs1 \IDinst/RegFile_reg[18][3]  ( .DIN(\IDinst/n5799 ), .CLK(clk), 
        .CLRB(n842), .SETB(1'b1), .Q(\IDinst/RegFile[18][3] ) );
  dffascs1 \IDinst/RegFile_reg[18][2]  ( .DIN(\IDinst/n5800 ), .CLK(clk), 
        .CLRB(n839), .SETB(1'b1), .Q(\IDinst/RegFile[18][2] ) );
  dffascs1 \IDinst/RegFile_reg[18][1]  ( .DIN(\IDinst/n5801 ), .CLK(clk), 
        .CLRB(n835), .SETB(1'b1), .Q(\IDinst/RegFile[18][1] ) );
  dffascs1 \IDinst/RegFile_reg[18][0]  ( .DIN(\IDinst/n5802 ), .CLK(clk), 
        .CLRB(n930), .SETB(1'b1), .Q(\IDinst/RegFile[18][0] ) );
  dffascs1 \IDinst/RegFile_reg[10][7]  ( .DIN(\IDinst/n5731 ), .CLK(clk), 
        .CLRB(n851), .SETB(1'b1), .Q(\IDinst/RegFile[10][7] ) );
  dffascs1 \IDinst/RegFile_reg[10][6]  ( .DIN(\IDinst/n5732 ), .CLK(clk), 
        .CLRB(n847), .SETB(1'b1), .Q(\IDinst/RegFile[10][6] ) );
  dffascs1 \IDinst/RegFile_reg[10][5]  ( .DIN(\IDinst/n5733 ), .CLK(clk), 
        .CLRB(n855), .SETB(1'b1), .Q(\IDinst/RegFile[10][5] ) );
  dffascs1 \IDinst/RegFile_reg[10][4]  ( .DIN(\IDinst/n5734 ), .CLK(clk), 
        .CLRB(n870), .SETB(1'b1), .Q(\IDinst/RegFile[10][4] ) );
  dffascs1 \IDinst/RegFile_reg[10][3]  ( .DIN(\IDinst/n5735 ), .CLK(clk), 
        .CLRB(n843), .SETB(1'b1), .Q(\IDinst/RegFile[10][3] ) );
  dffascs1 \IDinst/RegFile_reg[10][2]  ( .DIN(\IDinst/n5736 ), .CLK(clk), 
        .CLRB(n839), .SETB(1'b1), .Q(\IDinst/RegFile[10][2] ) );
  dffascs1 \IDinst/RegFile_reg[10][1]  ( .DIN(\IDinst/n5737 ), .CLK(clk), 
        .CLRB(n836), .SETB(1'b1), .Q(\IDinst/RegFile[10][1] ) );
  dffascs1 \IDinst/RegFile_reg[10][0]  ( .DIN(\IDinst/n5738 ), .CLK(clk), 
        .CLRB(n934), .SETB(1'b1), .Q(\IDinst/RegFile[10][0] ) );
  dffascs1 \IDinst/RegFile_reg[2][7]  ( .DIN(\IDinst/n5667 ), .CLK(clk), 
        .CLRB(n852), .SETB(1'b1), .Q(\IDinst/RegFile[2][7] ) );
  dffascs1 \IDinst/RegFile_reg[2][6]  ( .DIN(\IDinst/n5668 ), .CLK(clk), 
        .CLRB(n848), .SETB(1'b1), .Q(\IDinst/RegFile[2][6] ) );
  dffascs1 \IDinst/RegFile_reg[2][5]  ( .DIN(\IDinst/n5669 ), .CLK(clk), 
        .CLRB(n856), .SETB(1'b1), .Q(\IDinst/RegFile[2][5] ) );
  dffascs1 \IDinst/RegFile_reg[2][4]  ( .DIN(\IDinst/n5670 ), .CLK(clk), 
        .CLRB(n871), .SETB(1'b1), .Q(\IDinst/RegFile[2][4] ) );
  dffascs1 \IDinst/RegFile_reg[2][3]  ( .DIN(\IDinst/n5671 ), .CLK(clk), 
        .CLRB(n844), .SETB(1'b1), .Q(\IDinst/RegFile[2][3] ) );
  dffascs1 \IDinst/RegFile_reg[2][2]  ( .DIN(\IDinst/n5672 ), .CLK(clk), 
        .CLRB(n840), .SETB(1'b1), .Q(\IDinst/RegFile[2][2] ) );
  dffascs1 \IDinst/RegFile_reg[2][1]  ( .DIN(\IDinst/n5673 ), .CLK(clk), 
        .CLRB(n837), .SETB(1'b1), .Q(\IDinst/RegFile[2][1] ) );
  dffascs1 \IDinst/RegFile_reg[2][0]  ( .DIN(\IDinst/n5674 ), .CLK(clk), 
        .CLRB(n937), .SETB(1'b1), .Q(\IDinst/RegFile[2][0] ) );
  dffascs1 \IDinst/RegFile_reg[27][7]  ( .DIN(\IDinst/n5867 ), .CLK(clk), 
        .CLRB(n849), .SETB(1'b1), .Q(\IDinst/RegFile[27][7] ) );
  dffascs1 \IDinst/RegFile_reg[27][6]  ( .DIN(\IDinst/n5868 ), .CLK(clk), 
        .CLRB(n846), .SETB(1'b1), .Q(\IDinst/RegFile[27][6] ) );
  dffascs1 \IDinst/RegFile_reg[27][5]  ( .DIN(\IDinst/n5869 ), .CLK(clk), 
        .CLRB(n853), .SETB(1'b1), .Q(\IDinst/RegFile[27][5] ) );
  dffascs1 \IDinst/RegFile_reg[27][4]  ( .DIN(\IDinst/n5870 ), .CLK(clk), 
        .CLRB(n868), .SETB(1'b1), .Q(\IDinst/RegFile[27][4] ) );
  dffascs1 \IDinst/RegFile_reg[27][3]  ( .DIN(\IDinst/n5871 ), .CLK(clk), 
        .CLRB(n841), .SETB(1'b1), .Q(\IDinst/RegFile[27][3] ) );
  dffascs1 \IDinst/RegFile_reg[27][2]  ( .DIN(\IDinst/n5872 ), .CLK(clk), 
        .CLRB(n838), .SETB(1'b1), .Q(\IDinst/RegFile[27][2] ) );
  dffascs1 \IDinst/RegFile_reg[27][1]  ( .DIN(\IDinst/n5873 ), .CLK(clk), 
        .CLRB(n834), .SETB(1'b1), .Q(\IDinst/RegFile[27][1] ) );
  dffascs1 \IDinst/RegFile_reg[27][0]  ( .DIN(\IDinst/n5874 ), .CLK(clk), 
        .CLRB(n928), .SETB(1'b1), .Q(\IDinst/RegFile[27][0] ) );
  dffascs1 \IDinst/RegFile_reg[19][7]  ( .DIN(\IDinst/n5803 ), .CLK(clk), 
        .CLRB(n850), .SETB(1'b1), .Q(\IDinst/RegFile[19][7] ) );
  dffascs1 \IDinst/RegFile_reg[19][6]  ( .DIN(\IDinst/n5804 ), .CLK(clk), 
        .CLRB(n846), .SETB(1'b1), .Q(\IDinst/RegFile[19][6] ) );
  dffascs1 \IDinst/RegFile_reg[19][5]  ( .DIN(\IDinst/n5805 ), .CLK(clk), 
        .CLRB(n854), .SETB(1'b1), .Q(\IDinst/RegFile[19][5] ) );
  dffascs1 \IDinst/RegFile_reg[19][4]  ( .DIN(\IDinst/n5806 ), .CLK(clk), 
        .CLRB(n869), .SETB(1'b1), .Q(\IDinst/RegFile[19][4] ) );
  dffascs1 \IDinst/RegFile_reg[19][3]  ( .DIN(\IDinst/n5807 ), .CLK(clk), 
        .CLRB(n842), .SETB(1'b1), .Q(\IDinst/RegFile[19][3] ) );
  dffascs1 \IDinst/RegFile_reg[19][2]  ( .DIN(\IDinst/n5808 ), .CLK(clk), 
        .CLRB(n838), .SETB(1'b1), .Q(\IDinst/RegFile[19][2] ) );
  dffascs1 \IDinst/RegFile_reg[19][1]  ( .DIN(\IDinst/n5809 ), .CLK(clk), 
        .CLRB(n835), .SETB(1'b1), .Q(\IDinst/RegFile[19][1] ) );
  dffascs1 \IDinst/RegFile_reg[19][0]  ( .DIN(\IDinst/n5810 ), .CLK(clk), 
        .CLRB(n931), .SETB(1'b1), .Q(\IDinst/RegFile[19][0] ) );
  dffascs1 \IDinst/RegFile_reg[11][7]  ( .DIN(\IDinst/n5739 ), .CLK(clk), 
        .CLRB(n851), .SETB(1'b1), .Q(\IDinst/RegFile[11][7] ) );
  dffascs1 \IDinst/RegFile_reg[11][6]  ( .DIN(\IDinst/n5740 ), .CLK(clk), 
        .CLRB(n847), .SETB(1'b1), .Q(\IDinst/RegFile[11][6] ) );
  dffascs1 \IDinst/RegFile_reg[11][5]  ( .DIN(\IDinst/n5741 ), .CLK(clk), 
        .CLRB(n855), .SETB(1'b1), .Q(\IDinst/RegFile[11][5] ) );
  dffascs1 \IDinst/RegFile_reg[11][4]  ( .DIN(\IDinst/n5742 ), .CLK(clk), 
        .CLRB(n870), .SETB(1'b1), .Q(\IDinst/RegFile[11][4] ) );
  dffascs1 \IDinst/RegFile_reg[11][3]  ( .DIN(\IDinst/n5743 ), .CLK(clk), 
        .CLRB(n843), .SETB(1'b1), .Q(\IDinst/RegFile[11][3] ) );
  dffascs1 \IDinst/RegFile_reg[11][2]  ( .DIN(\IDinst/n5744 ), .CLK(clk), 
        .CLRB(n839), .SETB(1'b1), .Q(\IDinst/RegFile[11][2] ) );
  dffascs1 \IDinst/RegFile_reg[11][1]  ( .DIN(\IDinst/n5745 ), .CLK(clk), 
        .CLRB(n836), .SETB(1'b1), .Q(\IDinst/RegFile[11][1] ) );
  dffascs1 \IDinst/RegFile_reg[11][0]  ( .DIN(\IDinst/n5746 ), .CLK(clk), 
        .CLRB(n934), .SETB(1'b1), .Q(\IDinst/RegFile[11][0] ) );
  dffascs1 \IDinst/RegFile_reg[3][7]  ( .DIN(\IDinst/n5675 ), .CLK(clk), 
        .CLRB(n852), .SETB(1'b1), .Q(\IDinst/RegFile[3][7] ) );
  dffascs1 \IDinst/RegFile_reg[3][6]  ( .DIN(\IDinst/n5676 ), .CLK(clk), 
        .CLRB(n848), .SETB(1'b1), .Q(\IDinst/RegFile[3][6] ) );
  dffascs1 \IDinst/RegFile_reg[3][5]  ( .DIN(\IDinst/n5677 ), .CLK(clk), 
        .CLRB(n855), .SETB(1'b1), .Q(\IDinst/RegFile[3][5] ) );
  dffascs1 \IDinst/RegFile_reg[3][4]  ( .DIN(\IDinst/n5678 ), .CLK(clk), 
        .CLRB(n871), .SETB(1'b1), .Q(\IDinst/RegFile[3][4] ) );
  dffascs1 \IDinst/RegFile_reg[3][3]  ( .DIN(\IDinst/n5679 ), .CLK(clk), 
        .CLRB(n844), .SETB(1'b1), .Q(\IDinst/RegFile[3][3] ) );
  dffascs1 \IDinst/RegFile_reg[3][2]  ( .DIN(\IDinst/n5680 ), .CLK(clk), 
        .CLRB(n840), .SETB(1'b1), .Q(\IDinst/RegFile[3][2] ) );
  dffascs1 \IDinst/RegFile_reg[3][1]  ( .DIN(\IDinst/n5681 ), .CLK(clk), 
        .CLRB(n836), .SETB(1'b1), .Q(\IDinst/RegFile[3][1] ) );
  dffascs1 \IDinst/RegFile_reg[3][0]  ( .DIN(\IDinst/n5682 ), .CLK(clk), 
        .CLRB(n937), .SETB(1'b1), .Q(\IDinst/RegFile[3][0] ) );
  dffascs1 \IDinst/RegFile_reg[30][7]  ( .DIN(\IDinst/n5891 ), .CLK(clk), 
        .CLRB(n849), .SETB(1'b1), .Q(\IDinst/RegFile[30][7] ) );
  dffascs1 \IDinst/RegFile_reg[30][6]  ( .DIN(\IDinst/n5892 ), .CLK(clk), 
        .CLRB(n845), .SETB(1'b1), .Q(\IDinst/RegFile[30][6] ) );
  dffascs1 \IDinst/RegFile_reg[30][5]  ( .DIN(\IDinst/n5893 ), .CLK(clk), 
        .CLRB(n853), .SETB(1'b1), .Q(\IDinst/RegFile[30][5] ) );
  dffascs1 \IDinst/RegFile_reg[30][4]  ( .DIN(\IDinst/n5894 ), .CLK(clk), 
        .CLRB(n868), .SETB(1'b1), .Q(\IDinst/RegFile[30][4] ) );
  dffascs1 \IDinst/RegFile_reg[30][3]  ( .DIN(\IDinst/n5895 ), .CLK(clk), 
        .CLRB(n841), .SETB(1'b1), .Q(\IDinst/RegFile[30][3] ) );
  dffascs1 \IDinst/RegFile_reg[30][2]  ( .DIN(\IDinst/n5896 ), .CLK(clk), 
        .CLRB(n837), .SETB(1'b1), .Q(\IDinst/RegFile[30][2] ) );
  dffascs1 \IDinst/RegFile_reg[30][1]  ( .DIN(\IDinst/n5897 ), .CLK(clk), 
        .CLRB(n834), .SETB(1'b1), .Q(\IDinst/RegFile[30][1] ) );
  dffascs1 \IDinst/RegFile_reg[30][0]  ( .DIN(\IDinst/n5898 ), .CLK(clk), 
        .CLRB(n929), .SETB(1'b1), .Q(\IDinst/RegFile[30][0] ) );
  dffascs1 \IDinst/RegFile_reg[22][7]  ( .DIN(\IDinst/n5827 ), .CLK(clk), 
        .CLRB(n850), .SETB(1'b1), .Q(\IDinst/RegFile[22][7] ) );
  dffascs1 \IDinst/RegFile_reg[22][6]  ( .DIN(\IDinst/n5828 ), .CLK(clk), 
        .CLRB(n846), .SETB(1'b1), .Q(\IDinst/RegFile[22][6] ) );
  dffascs1 \IDinst/RegFile_reg[22][5]  ( .DIN(\IDinst/n5829 ), .CLK(clk), 
        .CLRB(n854), .SETB(1'b1), .Q(\IDinst/RegFile[22][5] ) );
  dffascs1 \IDinst/RegFile_reg[22][4]  ( .DIN(\IDinst/n5830 ), .CLK(clk), 
        .CLRB(n869), .SETB(1'b1), .Q(\IDinst/RegFile[22][4] ) );
  dffascs1 \IDinst/RegFile_reg[22][3]  ( .DIN(\IDinst/n5831 ), .CLK(clk), 
        .CLRB(n842), .SETB(1'b1), .Q(\IDinst/RegFile[22][3] ) );
  dffascs1 \IDinst/RegFile_reg[22][2]  ( .DIN(\IDinst/n5832 ), .CLK(clk), 
        .CLRB(n838), .SETB(1'b1), .Q(\IDinst/RegFile[22][2] ) );
  dffascs1 \IDinst/RegFile_reg[22][1]  ( .DIN(\IDinst/n5833 ), .CLK(clk), 
        .CLRB(n835), .SETB(1'b1), .Q(\IDinst/RegFile[22][1] ) );
  dffascs1 \IDinst/RegFile_reg[22][0]  ( .DIN(\IDinst/n5834 ), .CLK(clk), 
        .CLRB(n932), .SETB(1'b1), .Q(\IDinst/RegFile[22][0] ) );
  dffascs1 \IDinst/RegFile_reg[14][7]  ( .DIN(\IDinst/n5763 ), .CLK(clk), 
        .CLRB(n851), .SETB(1'b1), .Q(\IDinst/RegFile[14][7] ) );
  dffascs1 \IDinst/RegFile_reg[14][6]  ( .DIN(\IDinst/n5764 ), .CLK(clk), 
        .CLRB(n847), .SETB(1'b1), .Q(\IDinst/RegFile[14][6] ) );
  dffascs1 \IDinst/RegFile_reg[14][5]  ( .DIN(\IDinst/n5765 ), .CLK(clk), 
        .CLRB(n854), .SETB(1'b1), .Q(\IDinst/RegFile[14][5] ) );
  dffascs1 \IDinst/RegFile_reg[14][4]  ( .DIN(\IDinst/n5766 ), .CLK(clk), 
        .CLRB(n870), .SETB(1'b1), .Q(\IDinst/RegFile[14][4] ) );
  dffascs1 \IDinst/RegFile_reg[14][3]  ( .DIN(\IDinst/n5767 ), .CLK(clk), 
        .CLRB(n843), .SETB(1'b1), .Q(\IDinst/RegFile[14][3] ) );
  dffascs1 \IDinst/RegFile_reg[14][2]  ( .DIN(\IDinst/n5768 ), .CLK(clk), 
        .CLRB(n839), .SETB(1'b1), .Q(\IDinst/RegFile[14][2] ) );
  dffascs1 \IDinst/RegFile_reg[14][1]  ( .DIN(\IDinst/n5769 ), .CLK(clk), 
        .CLRB(n835), .SETB(1'b1), .Q(\IDinst/RegFile[14][1] ) );
  dffascs1 \IDinst/RegFile_reg[14][0]  ( .DIN(\IDinst/n5770 ), .CLK(clk), 
        .CLRB(n935), .SETB(1'b1), .Q(\IDinst/RegFile[14][0] ) );
  dffascs1 \IDinst/RegFile_reg[6][7]  ( .DIN(\IDinst/n5699 ), .CLK(clk), 
        .CLRB(n852), .SETB(1'b1), .Q(\IDinst/RegFile[6][7] ) );
  dffascs1 \IDinst/RegFile_reg[6][6]  ( .DIN(\IDinst/n5700 ), .CLK(clk), 
        .CLRB(n848), .SETB(1'b1), .Q(\IDinst/RegFile[6][6] ) );
  dffascs1 \IDinst/RegFile_reg[6][5]  ( .DIN(\IDinst/n5701 ), .CLK(clk), 
        .CLRB(n855), .SETB(1'b1), .Q(\IDinst/RegFile[6][5] ) );
  dffascs1 \IDinst/RegFile_reg[6][4]  ( .DIN(\IDinst/n5702 ), .CLK(clk), 
        .CLRB(n870), .SETB(1'b1), .Q(\IDinst/RegFile[6][4] ) );
  dffascs1 \IDinst/RegFile_reg[6][3]  ( .DIN(\IDinst/n5703 ), .CLK(clk), 
        .CLRB(n843), .SETB(1'b1), .Q(\IDinst/RegFile[6][3] ) );
  dffascs1 \IDinst/RegFile_reg[6][2]  ( .DIN(\IDinst/n5704 ), .CLK(clk), 
        .CLRB(n840), .SETB(1'b1), .Q(\IDinst/RegFile[6][2] ) );
  dffascs1 \IDinst/RegFile_reg[6][1]  ( .DIN(\IDinst/n5705 ), .CLK(clk), 
        .CLRB(n836), .SETB(1'b1), .Q(\IDinst/RegFile[6][1] ) );
  dffascs1 \IDinst/RegFile_reg[6][0]  ( .DIN(\IDinst/n5706 ), .CLK(clk), 
        .CLRB(n938), .SETB(1'b1), .Q(\IDinst/RegFile[6][0] ) );
  dffascs1 \IDinst/RegFile_reg[31][7]  ( .DIN(\IDinst/n5899 ), .CLK(clk), 
        .CLRB(n849), .SETB(1'b1), .Q(\IDinst/RegFile[31][7] ) );
  dffascs1 \IDinst/RegFile_reg[31][6]  ( .DIN(\IDinst/n5900 ), .CLK(clk), 
        .CLRB(n845), .SETB(1'b1), .Q(\IDinst/RegFile[31][6] ) );
  dffascs1 \IDinst/RegFile_reg[31][5]  ( .DIN(\IDinst/n5901 ), .CLK(clk), 
        .CLRB(n853), .SETB(1'b1), .Q(\IDinst/RegFile[31][5] ) );
  dffascs1 \IDinst/RegFile_reg[31][4]  ( .DIN(\IDinst/n5902 ), .CLK(clk), 
        .CLRB(n868), .SETB(1'b1), .Q(\IDinst/RegFile[31][4] ) );
  dffascs1 \IDinst/RegFile_reg[31][3]  ( .DIN(\IDinst/n5903 ), .CLK(clk), 
        .CLRB(n841), .SETB(1'b1), .Q(\IDinst/RegFile[31][3] ) );
  dffascs1 \IDinst/RegFile_reg[31][2]  ( .DIN(\IDinst/n5904 ), .CLK(clk), 
        .CLRB(n837), .SETB(1'b1), .Q(\IDinst/RegFile[31][2] ) );
  dffascs1 \IDinst/RegFile_reg[31][1]  ( .DIN(\IDinst/n5905 ), .CLK(clk), 
        .CLRB(n834), .SETB(1'b1), .Q(\IDinst/RegFile[31][1] ) );
  dffascs1 \IDinst/RegFile_reg[31][0]  ( .DIN(\IDinst/n5906 ), .CLK(clk), 
        .CLRB(n963), .SETB(1'b1), .Q(\IDinst/RegFile[31][0] ) );
  dffascs1 \IDinst/RegFile_reg[23][7]  ( .DIN(\IDinst/n5835 ), .CLK(clk), 
        .CLRB(n850), .SETB(1'b1), .Q(\IDinst/RegFile[23][7] ) );
  dffascs1 \IDinst/RegFile_reg[23][6]  ( .DIN(\IDinst/n5836 ), .CLK(clk), 
        .CLRB(n846), .SETB(1'b1), .Q(\IDinst/RegFile[23][6] ) );
  dffascs1 \IDinst/RegFile_reg[23][5]  ( .DIN(\IDinst/n5837 ), .CLK(clk), 
        .CLRB(n853), .SETB(1'b1), .Q(\IDinst/RegFile[23][5] ) );
  dffascs1 \IDinst/RegFile_reg[23][4]  ( .DIN(\IDinst/n5838 ), .CLK(clk), 
        .CLRB(n869), .SETB(1'b1), .Q(\IDinst/RegFile[23][4] ) );
  dffascs1 \IDinst/RegFile_reg[23][3]  ( .DIN(\IDinst/n5839 ), .CLK(clk), 
        .CLRB(n842), .SETB(1'b1), .Q(\IDinst/RegFile[23][3] ) );
  dffascs1 \IDinst/RegFile_reg[23][2]  ( .DIN(\IDinst/n5840 ), .CLK(clk), 
        .CLRB(n838), .SETB(1'b1), .Q(\IDinst/RegFile[23][2] ) );
  dffascs1 \IDinst/RegFile_reg[23][1]  ( .DIN(\IDinst/n5841 ), .CLK(clk), 
        .CLRB(n834), .SETB(1'b1), .Q(\IDinst/RegFile[23][1] ) );
  dffascs1 \IDinst/RegFile_reg[23][0]  ( .DIN(\IDinst/n5842 ), .CLK(clk), 
        .CLRB(n932), .SETB(1'b1), .Q(\IDinst/RegFile[23][0] ) );
  dffascs1 \IDinst/RegFile_reg[15][7]  ( .DIN(\IDinst/n5771 ), .CLK(clk), 
        .CLRB(n851), .SETB(1'b1), .Q(\IDinst/RegFile[15][7] ) );
  dffascs1 \IDinst/RegFile_reg[15][6]  ( .DIN(\IDinst/n5772 ), .CLK(clk), 
        .CLRB(n847), .SETB(1'b1), .Q(\IDinst/RegFile[15][6] ) );
  dffascs1 \IDinst/RegFile_reg[15][5]  ( .DIN(\IDinst/n5773 ), .CLK(clk), 
        .CLRB(n854), .SETB(1'b1), .Q(\IDinst/RegFile[15][5] ) );
  dffascs1 \IDinst/RegFile_reg[15][4]  ( .DIN(\IDinst/n5774 ), .CLK(clk), 
        .CLRB(n870), .SETB(1'b1), .Q(\IDinst/RegFile[15][4] ) );
  dffascs1 \IDinst/RegFile_reg[15][3]  ( .DIN(\IDinst/n5775 ), .CLK(clk), 
        .CLRB(n842), .SETB(1'b1), .Q(\IDinst/RegFile[15][3] ) );
  dffascs1 \IDinst/RegFile_reg[15][2]  ( .DIN(\IDinst/n5776 ), .CLK(clk), 
        .CLRB(n839), .SETB(1'b1), .Q(\IDinst/RegFile[15][2] ) );
  dffascs1 \IDinst/RegFile_reg[15][1]  ( .DIN(\IDinst/n5777 ), .CLK(clk), 
        .CLRB(n835), .SETB(1'b1), .Q(\IDinst/RegFile[15][1] ) );
  dffascs1 \IDinst/RegFile_reg[15][0]  ( .DIN(\IDinst/n5778 ), .CLK(clk), 
        .CLRB(n936), .SETB(1'b1), .Q(\IDinst/RegFile[15][0] ) );
  dffascs1 \IDinst/RegFile_reg[7][7]  ( .DIN(\IDinst/n5707 ), .CLK(clk), 
        .CLRB(n851), .SETB(1'b1), .Q(\IDinst/RegFile[7][7] ) );
  dffascs1 \IDinst/RegFile_reg[7][6]  ( .DIN(\IDinst/n5708 ), .CLK(clk), 
        .CLRB(n848), .SETB(1'b1), .Q(\IDinst/RegFile[7][6] ) );
  dffascs1 \IDinst/RegFile_reg[7][5]  ( .DIN(\IDinst/n5709 ), .CLK(clk), 
        .CLRB(n855), .SETB(1'b1), .Q(\IDinst/RegFile[7][5] ) );
  dffascs1 \IDinst/RegFile_reg[7][4]  ( .DIN(\IDinst/n5710 ), .CLK(clk), 
        .CLRB(n870), .SETB(1'b1), .Q(\IDinst/RegFile[7][4] ) );
  dffascs1 \IDinst/RegFile_reg[7][3]  ( .DIN(\IDinst/n5711 ), .CLK(clk), 
        .CLRB(n843), .SETB(1'b1), .Q(\IDinst/RegFile[7][3] ) );
  dffascs1 \IDinst/RegFile_reg[7][2]  ( .DIN(\IDinst/n5712 ), .CLK(clk), 
        .CLRB(n840), .SETB(1'b1), .Q(\IDinst/RegFile[7][2] ) );
  dffascs1 \IDinst/RegFile_reg[7][1]  ( .DIN(\IDinst/n5713 ), .CLK(clk), 
        .CLRB(n836), .SETB(1'b1), .Q(\IDinst/RegFile[7][1] ) );
  dffascs1 \IDinst/RegFile_reg[7][0]  ( .DIN(\IDinst/n5714 ), .CLK(clk), 
        .CLRB(n939), .SETB(1'b1), .Q(\IDinst/RegFile[7][0] ) );
  dffascs1 \IDinst/WB_index_reg[1]  ( .DIN(\IDinst/reg_dst_of_MEM[1]), 
        .CLK(clk), .CLRB(n942), .SETB(1'b1), .Q(n58), .QN(\IDinst/n1432 ) );
  dffascs1 \IDinst/reg_dst_of_MEM_reg[1]  ( .DIN(\IDinst/reg_dst_of_EX[1]), 
        .CLK(clk), .CLRB(n942), .SETB(1'b1), .Q(\IDinst/reg_dst_of_MEM[1]), 
        .QN(n9455) );
  dffascs1 \IDinst/rt_addr_reg[1]  ( .DIN(\IDinst/n4864 ), .CLK(clk), 
        .CLRB(n942), .SETB(1'b1), .Q(n228), .QN(n9409) );
  dffascs1 \IDinst/WB_index_reg[2]  ( .DIN(\IDinst/reg_dst_of_MEM[2]), 
        .CLK(clk), .CLRB(n942), .SETB(1'b1), .Q(n203), .QN(\IDinst/n1431 ) );
  dffascs1 \IDinst/reg_dst_of_MEM_reg[2]  ( .DIN(\IDinst/reg_dst_of_EX[2]), 
        .CLK(clk), .CLRB(n942), .SETB(1'b1), .Q(\IDinst/reg_dst_of_MEM[2]), 
        .QN(n9421) );
  dffascs1 \IDinst/rt_addr_reg[2]  ( .DIN(\IDinst/n4863 ), .CLK(clk), 
        .CLRB(n942), .SETB(1'b1), .Q(n227), .QN(n9411) );
  dffascs1 \IDinst/WB_index_reg[3]  ( .DIN(\IDinst/reg_dst_of_MEM[3]), 
        .CLK(clk), .CLRB(n942), .SETB(1'b1), .Q(n47), .QN(\IDinst/n1430 ) );
  dffascs1 \IDinst/reg_dst_of_MEM_reg[3]  ( .DIN(\IDinst/reg_dst_of_EX[3]), 
        .CLK(clk), .CLRB(n943), .SETB(1'b1), .Q(\IDinst/reg_dst_of_MEM[3]), 
        .QN(n9420) );
  dffascs1 \IDinst/rt_addr_reg[3]  ( .DIN(\IDinst/n4862 ), .CLK(clk), 
        .CLRB(n943), .SETB(1'b1), .Q(n49) );
  dffascs1 \IDinst/WB_index_reg[4]  ( .DIN(\IDinst/reg_dst_of_MEM[4]), 
        .CLK(clk), .CLRB(n943), .SETB(1'b1), .Q(n376), .QN(\IDinst/n1403 ) );
  dffascs1 \IDinst/reg_dst_of_MEM_reg[4]  ( .DIN(\IDinst/reg_dst_of_EX[4]), 
        .CLK(clk), .CLRB(n943), .SETB(1'b1), .Q(\IDinst/reg_dst_of_MEM[4]), 
        .QN(n9419) );
  dffascs1 \IDinst/rt_addr_reg[4]  ( .DIN(\IDinst/n4861 ), .CLK(clk), 
        .CLRB(n943), .SETB(1'b1), .Q(n141) );
  dffascs1 \IDinst/reg_dst_reg  ( .DIN(\IDinst/n4867 ), .CLK(clk), .CLRB(n944), 
        .SETB(1'b1), .Q(reg_dst), .QN(n11) );
  dffascs1 \IDinst/reg_write_reg  ( .DIN(\IDinst/n4868 ), .CLK(clk), 
        .CLRB(n939), .SETB(1'b1), .Q(reg_write) );
  dffascs1 \IDinst/delay_slot_reg  ( .DIN(\IDinst/n4859 ), .CLK(clk), 
        .CLRB(n962), .SETB(1'b1), .Q(n119), .QN(\IDinst/n1440 ) );
  dffascs1 \IDinst/rd_addr_reg[1]  ( .DIN(\IDinst/n5910 ), .CLK(clk), 
        .CLRB(n943), .SETB(1'b1), .Q(n231), .QN(n9410) );
  dffascs1 \IDinst/rd_addr_reg[2]  ( .DIN(\IDinst/n5909 ), .CLK(clk), 
        .CLRB(n943), .SETB(1'b1), .Q(n230), .QN(n9412) );
  dffascs1 \IDinst/rd_addr_reg[3]  ( .DIN(\IDinst/n5908 ), .CLK(clk), 
        .CLRB(n943), .SETB(1'b1), .Q(n50) );
  dffascs1 \IDinst/rd_addr_reg[4]  ( .DIN(\IDinst/n5907 ), .CLK(clk), 
        .CLRB(n943), .SETB(1'b1), .Q(n142) );
  dffascs1 \IDinst/IR_function_field_reg[5]  ( .DIN(\IDinst/n4871 ), .CLK(clk), 
        .CLRB(n944), .SETB(1'b1), .Q(n377), .QN(n9454) );
  dffascs1 \IDinst/mem_write_reg  ( .DIN(\IDinst/n4869 ), .CLK(clk), 
        .CLRB(n926), .SETB(1'b1), .QN(n9415) );
  dffascs1 \IDinst/current_IR_reg[31]  ( .DIN(\IDinst/n5943 ), .CLK(clk), 
        .CLRB(n809), .SETB(1'b1), .Q(n323) );
  dffascs1 \IDinst/mem_read_reg  ( .DIN(\IDinst/n4870 ), .CLK(clk), 
        .CLRB(n926), .SETB(1'b1), .QN(n9414) );
  dffascs1 \IDinst/current_IR_reg[28]  ( .DIN(\IDinst/n5914 ), .CLK(clk), 
        .CLRB(n951), .SETB(1'b1), .Q(n325) );
  dffascs1 \IDinst/current_IR_reg[29]  ( .DIN(\IDinst/n5913 ), .CLK(clk), 
        .CLRB(n951), .SETB(1'b1), .Q(n327) );
  dffascs1 \IDinst/current_IR_reg[26]  ( .DIN(\IDinst/n5916 ), .CLK(clk), 
        .CLRB(n952), .SETB(1'b1), .Q(n319) );
  dffascs1 \IDinst/current_IR_reg[30]  ( .DIN(\IDinst/n5912 ), .CLK(clk), 
        .CLRB(n926), .SETB(1'b1), .Q(n317) );
  dffascs1 \IDinst/current_IR_reg[27]  ( .DIN(\IDinst/n5915 ), .CLK(clk), 
        .CLRB(n951), .SETB(1'b1), .Q(n321) );
  dffascs1 \IDinst/current_IR_reg[25]  ( .DIN(\IDinst/n5917 ), .CLK(clk), 
        .CLRB(n952), .SETB(1'b1), .Q(n311) );
  dffascs1 \IDinst/current_IR_reg[24]  ( .DIN(\IDinst/n5918 ), .CLK(clk), 
        .CLRB(n952), .SETB(1'b1), .Q(n315) );
  dffascs1 \IDinst/current_IR_reg[23]  ( .DIN(\IDinst/n5919 ), .CLK(clk), 
        .CLRB(n953), .SETB(1'b1), .Q(n313) );
  dffascs1 \IDinst/current_IR_reg[22]  ( .DIN(\IDinst/n5920 ), .CLK(clk), 
        .CLRB(n953), .SETB(1'b1), .Q(n307) );
  dffascs1 \IDinst/current_IR_reg[21]  ( .DIN(\IDinst/n5921 ), .CLK(clk), 
        .CLRB(n953), .SETB(1'b1), .Q(n309) );
  dffascs1 \IDinst/current_IR_reg[20]  ( .DIN(\IDinst/n5922 ), .CLK(clk), 
        .CLRB(n954), .SETB(1'b1), .Q(n277) );
  dffascs1 \IDinst/current_IR_reg[19]  ( .DIN(\IDinst/n5923 ), .CLK(clk), 
        .CLRB(n954), .SETB(1'b1), .Q(n281) );
  dffascs1 \IDinst/current_IR_reg[18]  ( .DIN(\IDinst/n5924 ), .CLK(clk), 
        .CLRB(n954), .SETB(1'b1), .Q(n279) );
  dffascs1 \IDinst/current_IR_reg[17]  ( .DIN(\IDinst/n5925 ), .CLK(clk), 
        .CLRB(n954), .SETB(1'b1), .Q(n275) );
  dffascs1 \IDinst/current_IR_reg[16]  ( .DIN(\IDinst/n5926 ), .CLK(clk), 
        .CLRB(n955), .SETB(1'b1), .Q(n273) );
  dffascs1 \IDinst/counter_reg[0]  ( .DIN(\IDinst/n5944 ), .CLK(clk), 
        .CLRB(n962), .SETB(1'b1), .Q(n48), .QN(n9453) );
  dffascs1 \IDinst/intr_slot_reg  ( .DIN(\IDinst/n5946 ), .CLK(clk), 
        .CLRB(n962), .SETB(1'b1), .Q(n215), .QN(\IDinst/n1445 ) );
  dffascs1 \IDinst/slot_num_reg[1]  ( .DIN(\IDinst/n4858 ), .CLK(clk), 
        .CLRB(n950), .SETB(1'b1), .Q(\IDinst/slot_num[1]), .QN(n60) );
  dffascs1 \IDinst/slot_num_reg[0]  ( .DIN(\IDinst/n4857 ), .CLK(clk), 
        .CLRB(n950), .SETB(1'b1), .Q(\IDinst/slot_num[0]), .QN(n378) );
  dffascs1 \IDinst/stall_reg  ( .DIN(\IDinst/n5945 ), .CLK(clk), .CLRB(n962), 
        .SETB(1'b1), .Q(stall) );
  dffascs1 \IDinst/rd_addr_reg[0]  ( .DIN(\IDinst/n5911 ), .CLK(clk), 
        .CLRB(n943), .SETB(1'b1), .Q(n232), .QN(n9408) );
  dffascs1 \IDinst/WB_index_reg[0]  ( .DIN(\IDinst/reg_dst_of_MEM[0]), 
        .CLK(clk), .CLRB(n942), .SETB(1'b1), .Q(n27), .QN(\IDinst/n1433 ) );
  dffascs1 \IDinst/reg_dst_of_MEM_reg[0]  ( .DIN(\IDinst/reg_dst_of_EX[0]), 
        .CLK(clk), .CLRB(n942), .SETB(1'b1), .Q(\IDinst/reg_dst_of_MEM[0]), 
        .QN(n9452) );
  dffascs1 \EXinst/mem_to_reg_EX_reg  ( .DIN(\EXinst/N1338 ), .CLK(clk), 
        .CLRB(n941), .SETB(1'b1), .Q(n374), .QN(n28) );
  dffascs1 \EXinst/reg_out_B_EX_reg[0]  ( .DIN(\EXinst/N1305 ), .CLK(clk), 
        .CLRB(n962), .SETB(1'b1), .Q(\DM_write_data[0] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[1]  ( .DIN(\EXinst/N1306 ), .CLK(clk), 
        .CLRB(n829), .SETB(1'b1), .Q(\DM_write_data[1] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[2]  ( .DIN(\EXinst/N1307 ), .CLK(clk), 
        .CLRB(n837), .SETB(1'b1), .Q(\DM_write_data[2] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[3]  ( .DIN(\EXinst/N1308 ), .CLK(clk), 
        .CLRB(n841), .SETB(1'b1), .Q(\DM_write_data[3] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[4]  ( .DIN(\EXinst/N1309 ), .CLK(clk), 
        .CLRB(n868), .SETB(1'b1), .Q(\DM_write_data[4] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[5]  ( .DIN(\EXinst/N1310 ), .CLK(clk), 
        .CLRB(n852), .SETB(1'b1), .Q(\DM_write_data[5] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[6]  ( .DIN(\EXinst/N1311 ), .CLK(clk), 
        .CLRB(n829), .SETB(1'b1), .Q(\DM_write_data[6] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[7]  ( .DIN(\EXinst/N1312 ), .CLK(clk), 
        .CLRB(n828), .SETB(1'b1), .Q(\DM_write_data[7] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[8]  ( .DIN(\EXinst/N1313 ), .CLK(clk), 
        .CLRB(n895), .SETB(1'b1), .Q(\DM_write_data[8] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[9]  ( .DIN(\EXinst/N1314 ), .CLK(clk), 
        .CLRB(n828), .SETB(1'b1), .Q(\DM_write_data[9] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[10]  ( .DIN(\EXinst/N1315 ), .CLK(clk), 
        .CLRB(n828), .SETB(1'b1), .Q(\DM_write_data[10] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[11]  ( .DIN(\EXinst/N1316 ), .CLK(clk), 
        .CLRB(n811), .SETB(1'b1), .Q(\DM_write_data[11] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[12]  ( .DIN(\EXinst/N1317 ), .CLK(clk), 
        .CLRB(n914), .SETB(1'b1), .Q(\DM_write_data[12] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[13]  ( .DIN(\EXinst/N1318 ), .CLK(clk), 
        .CLRB(n812), .SETB(1'b1), .Q(\DM_write_data[13] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[14]  ( .DIN(\EXinst/N1319 ), .CLK(clk), 
        .CLRB(n820), .SETB(1'b1), .Q(\DM_write_data[14] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[15]  ( .DIN(\EXinst/N1320 ), .CLK(clk), 
        .CLRB(n821), .SETB(1'b1), .Q(\DM_write_data[15] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[16]  ( .DIN(\EXinst/N1321 ), .CLK(clk), 
        .CLRB(n922), .SETB(1'b1), .Q(\DM_write_data[16] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[17]  ( .DIN(\EXinst/N1322 ), .CLK(clk), 
        .CLRB(n816), .SETB(1'b1), .Q(\DM_write_data[17] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[18]  ( .DIN(\EXinst/N1323 ), .CLK(clk), 
        .CLRB(n812), .SETB(1'b1), .Q(\DM_write_data[18] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[19]  ( .DIN(\EXinst/N1324 ), .CLK(clk), 
        .CLRB(n813), .SETB(1'b1), .Q(\DM_write_data[19] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[20]  ( .DIN(\EXinst/N1325 ), .CLK(clk), 
        .CLRB(n811), .SETB(1'b1), .Q(\DM_write_data[20] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[21]  ( .DIN(\EXinst/N1326 ), .CLK(clk), 
        .CLRB(n824), .SETB(1'b1), .Q(\DM_write_data[21] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[22]  ( .DIN(\EXinst/N1327 ), .CLK(clk), 
        .CLRB(n811), .SETB(1'b1), .Q(\DM_write_data[22] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[23]  ( .DIN(\EXinst/N1328 ), .CLK(clk), 
        .CLRB(n811), .SETB(1'b1), .Q(\DM_write_data[23] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[24]  ( .DIN(\EXinst/N1329 ), .CLK(clk), 
        .CLRB(n810), .SETB(1'b1), .Q(\DM_write_data[24] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[25]  ( .DIN(\EXinst/N1330 ), .CLK(clk), 
        .CLRB(n810), .SETB(1'b1), .Q(\DM_write_data[25] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[26]  ( .DIN(\EXinst/N1331 ), .CLK(clk), 
        .CLRB(n810), .SETB(1'b1), .Q(\DM_write_data[26] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[27]  ( .DIN(\EXinst/N1332 ), .CLK(clk), 
        .CLRB(n810), .SETB(1'b1), .Q(\DM_write_data[27] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[28]  ( .DIN(\EXinst/N1333 ), .CLK(clk), 
        .CLRB(n809), .SETB(1'b1), .Q(\DM_write_data[28] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[29]  ( .DIN(\EXinst/N1334 ), .CLK(clk), 
        .CLRB(n809), .SETB(1'b1), .Q(\DM_write_data[29] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[30]  ( .DIN(\EXinst/N1335 ), .CLK(clk), 
        .CLRB(n940), .SETB(1'b1), .Q(\DM_write_data[30] ) );
  dffascs1 \EXinst/reg_out_B_EX_reg[31]  ( .DIN(\EXinst/N1336 ), .CLK(clk), 
        .CLRB(n940), .SETB(1'b1), .Q(\DM_write_data[31] ) );
  dffascs1 \EXinst/byte_reg  ( .DIN(\EXinst/n1387 ), .CLK(clk), .CLRB(n939), 
        .SETB(1'b1), .Q(byte), .QN(n9417) );
  dffascs1 \EXinst/ALU_result_reg[0]  ( .DIN(\EXinst/n1432 ), .CLK(clk), 
        .CLRB(n963), .SETB(1'b1), .Q(\DM_addr[0] ) );
  dffascs1 \EXinst/ALU_result_reg[1]  ( .DIN(\EXinst/n1433 ), .CLK(clk), 
        .CLRB(n837), .SETB(1'b1), .Q(\DM_addr[1] ) );
  dffascs1 \EXinst/ALU_result_reg[2]  ( .DIN(\EXinst/n1434 ), .CLK(clk), 
        .CLRB(n841), .SETB(1'b1), .Q(\DM_addr[2] ) );
  dffascs1 \EXinst/ALU_result_reg[3]  ( .DIN(\EXinst/n1435 ), .CLK(clk), 
        .CLRB(n844), .SETB(1'b1), .Q(\DM_addr[3] ) );
  dffascs1 \EXinst/ALU_result_reg[4]  ( .DIN(\EXinst/n1436 ), .CLK(clk), 
        .CLRB(n871), .SETB(1'b1), .Q(\DM_addr[4] ) );
  dffascs1 \EXinst/ALU_result_reg[5]  ( .DIN(\EXinst/n1437 ), .CLK(clk), 
        .CLRB(n856), .SETB(1'b1), .Q(\DM_addr[5] ) );
  dffascs1 \EXinst/ALU_result_reg[6]  ( .DIN(\EXinst/n1438 ), .CLK(clk), 
        .CLRB(n849), .SETB(1'b1), .Q(\DM_addr[6] ) );
  dffascs1 \EXinst/ALU_result_reg[7]  ( .DIN(\EXinst/n1439 ), .CLK(clk), 
        .CLRB(n852), .SETB(1'b1), .Q(\DM_addr[7] ) );
  dffascs1 \EXinst/ALU_result_reg[8]  ( .DIN(\EXinst/n1440 ), .CLK(clk), 
        .CLRB(n899), .SETB(1'b1), .Q(\DM_addr[8] ) );
  dffascs1 \EXinst/ALU_result_reg[9]  ( .DIN(\EXinst/n1441 ), .CLK(clk), 
        .CLRB(n864), .SETB(1'b1), .Q(\DM_addr[9] ) );
  dffascs1 \EXinst/ALU_result_reg[10]  ( .DIN(\EXinst/n1442 ), .CLK(clk), 
        .CLRB(n860), .SETB(1'b1), .Q(\DM_addr[10] ) );
  dffascs1 \EXinst/ALU_result_reg[11]  ( .DIN(\EXinst/n1443 ), .CLK(clk), 
        .CLRB(n895), .SETB(1'b1), .Q(\DM_addr[11] ) );
  dffascs1 \EXinst/ALU_result_reg[12]  ( .DIN(\EXinst/n1444 ), .CLK(clk), 
        .CLRB(n918), .SETB(1'b1), .Q(\DM_addr[12] ) );
  dffascs1 \EXinst/ALU_result_reg[13]  ( .DIN(\EXinst/n1445 ), .CLK(clk), 
        .CLRB(n879), .SETB(1'b1), .Q(\DM_addr[13] ) );
  dffascs1 \EXinst/ALU_result_reg[14]  ( .DIN(\EXinst/n1446 ), .CLK(clk), 
        .CLRB(n868), .SETB(1'b1), .Q(\DM_addr[14] ) );
  dffascs1 \EXinst/ALU_result_reg[15]  ( .DIN(\EXinst/n1447 ), .CLK(clk), 
        .CLRB(n828), .SETB(1'b1), .Q(\DM_addr[15] ) );
  dffascs1 \EXinst/ALU_result_reg[16]  ( .DIN(\EXinst/n1448 ), .CLK(clk), 
        .CLRB(n914), .SETB(1'b1), .Q(\DM_addr[16] ) );
  dffascs1 \EXinst/ALU_result_reg[17]  ( .DIN(\EXinst/n1449 ), .CLK(clk), 
        .CLRB(n820), .SETB(1'b1), .Q(\DM_addr[17] ) );
  dffascs1 \EXinst/ALU_result_reg[18]  ( .DIN(\EXinst/n1450 ), .CLK(clk), 
        .CLRB(n875), .SETB(1'b1), .Q(\DM_addr[18] ) );
  dffascs1 \EXinst/ALU_result_reg[19]  ( .DIN(\EXinst/n1451 ), .CLK(clk), 
        .CLRB(n816), .SETB(1'b1), .Q(\DM_addr[19] ) );
  dffascs1 \EXinst/ALU_result_reg[20]  ( .DIN(\EXinst/n1452 ), .CLK(clk), 
        .CLRB(n888), .SETB(1'b1), .Q(\DM_addr[20] ) );
  dffascs1 \EXinst/ALU_result_reg[21]  ( .DIN(\EXinst/n1453 ), .CLK(clk), 
        .CLRB(n824), .SETB(1'b1), .Q(\DM_addr[21] ) );
  dffascs1 \EXinst/ALU_result_reg[22]  ( .DIN(\EXinst/n1454 ), .CLK(clk), 
        .CLRB(n884), .SETB(1'b1), .Q(\DM_addr[22] ) );
  dffascs1 \EXinst/ALU_result_reg[23]  ( .DIN(\EXinst/n1455 ), .CLK(clk), 
        .CLRB(n891), .SETB(1'b1), .Q(\DM_addr[23] ) );
  dffascs1 \EXinst/ALU_result_reg[24]  ( .DIN(\EXinst/n1456 ), .CLK(clk), 
        .CLRB(n906), .SETB(1'b1), .Q(\DM_addr[24] ) );
  dffascs1 \EXinst/ALU_result_reg[25]  ( .DIN(\EXinst/n1457 ), .CLK(clk), 
        .CLRB(n902), .SETB(1'b1), .Q(\DM_addr[25] ) );
  dffascs1 \EXinst/ALU_result_reg[26]  ( .DIN(\EXinst/n1458 ), .CLK(clk), 
        .CLRB(n913), .SETB(1'b1), .Q(\DM_addr[26] ) );
  dffascs1 \EXinst/ALU_result_reg[27]  ( .DIN(\EXinst/n1459 ), .CLK(clk), 
        .CLRB(n910), .SETB(1'b1), .Q(\DM_addr[27] ) );
  dffascs1 \EXinst/ALU_result_reg[28]  ( .DIN(\EXinst/n1460 ), .CLK(clk), 
        .CLRB(n922), .SETB(1'b1), .Q(\DM_addr[28] ) );
  dffascs1 \EXinst/ALU_result_reg[29]  ( .DIN(\EXinst/n1461 ), .CLK(clk), 
        .CLRB(n962), .SETB(1'b1), .Q(\DM_addr[29] ) );
  dffascs1 \EXinst/ALU_result_reg[30]  ( .DIN(\EXinst/n1462 ), .CLK(clk), 
        .CLRB(n963), .SETB(1'b1), .Q(\DM_addr[30] ) );
  dffascs1 \EXinst/ALU_result_reg[31]  ( .DIN(\EXinst/n1463 ), .CLK(clk), 
        .CLRB(n1018), .SETB(1'b1), .Q(\DM_addr[31] ) );
  dffascs1 \EXinst/mem_sign_ext_reg  ( .DIN(\EXinst/N1339 ), .CLK(clk), 
        .CLRB(n940), .SETB(1'b1), .Q(n380), .QN(n9418) );
  dffascs1 \EXinst/mem_write_EX_reg  ( .DIN(\EXinst/N1341 ), .CLK(clk), 
        .CLRB(n926), .SETB(1'b1), .Q(DM_write) );
  dffascs1 \EXinst/word_reg  ( .DIN(\EXinst/n1423 ), .CLK(clk), .CLRB(n940), 
        .SETB(1'b1), .Q(word) );
  dffascs1 \EXinst/reg_write_EX_reg  ( .DIN(\EXinst/N1337 ), .CLK(clk), 
        .CLRB(n939), .SETB(1'b1), .Q(reg_write_EX) );
  dffascs1 \EXinst/mem_read_EX_reg  ( .DIN(\EXinst/N1340 ), .CLK(clk), 
        .CLRB(n926), .SETB(1'b1), .Q(DM_read) );
  dffascs1 \MEMinst/reg_write_MEM_reg  ( .DIN(reg_write_EX), .CLK(clk), 
        .CLRB(n939), .SETB(1'b1), .Q(reg_write_MEM) );
  dffascs1 \MEMinst/RF_data_in_reg[0]  ( .DIN(\MEMinst/N57 ), .CLK(clk), 
        .CLRB(n963), .SETB(1'b1), .QN(n9393) );
  dffascs1 \MEMinst/RF_data_in_reg[1]  ( .DIN(\MEMinst/N58 ), .CLK(clk), 
        .CLRB(n837), .SETB(1'b1), .QN(n9394) );
  dffascs1 \MEMinst/RF_data_in_reg[2]  ( .DIN(\MEMinst/N59 ), .CLK(clk), 
        .CLRB(n840), .SETB(1'b1), .QN(n9395) );
  dffascs1 \MEMinst/RF_data_in_reg[3]  ( .DIN(\MEMinst/N60 ), .CLK(clk), 
        .CLRB(n844), .SETB(1'b1), .QN(n9396) );
  dffascs1 \MEMinst/RF_data_in_reg[4]  ( .DIN(\MEMinst/N61 ), .CLK(clk), 
        .CLRB(n871), .SETB(1'b1), .QN(n9397) );
  dffascs1 \MEMinst/RF_data_in_reg[5]  ( .DIN(\MEMinst/N62 ), .CLK(clk), 
        .CLRB(n856), .SETB(1'b1), .QN(n9398) );
  dffascs1 \MEMinst/RF_data_in_reg[6]  ( .DIN(\MEMinst/N63 ), .CLK(clk), 
        .CLRB(n848), .SETB(1'b1), .QN(n9399) );
  dffascs1 \MEMinst/RF_data_in_reg[7]  ( .DIN(\MEMinst/N64 ), .CLK(clk), 
        .CLRB(n852), .SETB(1'b1), .QN(n9404) );
  dffascs1 \MEMinst/RF_data_in_reg[8]  ( .DIN(\MEMinst/N65 ), .CLK(clk), 
        .CLRB(n898), .SETB(1'b1), .Q(n200) );
  dffascs1 \MEMinst/RF_data_in_reg[9]  ( .DIN(\MEMinst/N66 ), .CLK(clk), 
        .CLRB(n863), .SETB(1'b1), .Q(n198) );
  dffascs1 \MEMinst/RF_data_in_reg[10]  ( .DIN(\MEMinst/N67 ), .CLK(clk), 
        .CLRB(n860), .SETB(1'b1), .Q(n196) );
  dffascs1 \MEMinst/RF_data_in_reg[11]  ( .DIN(\MEMinst/N68 ), .CLK(clk), 
        .CLRB(n895), .SETB(1'b1), .Q(n194) );
  dffascs1 \MEMinst/RF_data_in_reg[12]  ( .DIN(\MEMinst/N69 ), .CLK(clk), 
        .CLRB(n918), .SETB(1'b1), .Q(n192) );
  dffascs1 \MEMinst/RF_data_in_reg[13]  ( .DIN(\MEMinst/N70 ), .CLK(clk), 
        .CLRB(n879), .SETB(1'b1), .Q(n190) );
  dffascs1 \MEMinst/RF_data_in_reg[14]  ( .DIN(\MEMinst/N71 ), .CLK(clk), 
        .CLRB(n868), .SETB(1'b1), .Q(n188) );
  dffascs1 \MEMinst/RF_data_in_reg[15]  ( .DIN(\MEMinst/N72 ), .CLK(clk), 
        .CLRB(n828), .SETB(1'b1), .Q(n129) );
  dffascs1 \MEMinst/RF_data_in_reg[16]  ( .DIN(\MEMinst/N73 ), .CLK(clk), 
        .CLRB(n914), .SETB(1'b1), .Q(n185) );
  dffascs1 \MEMinst/RF_data_in_reg[17]  ( .DIN(\MEMinst/N74 ), .CLK(clk), 
        .CLRB(n820), .SETB(1'b1), .Q(n183) );
  dffascs1 \MEMinst/RF_data_in_reg[18]  ( .DIN(\MEMinst/N75 ), .CLK(clk), 
        .CLRB(n875), .SETB(1'b1), .Q(n181) );
  dffascs1 \MEMinst/RF_data_in_reg[19]  ( .DIN(\MEMinst/N76 ), .CLK(clk), 
        .CLRB(n816), .SETB(1'b1), .Q(n179) );
  dffascs1 \MEMinst/RF_data_in_reg[20]  ( .DIN(\MEMinst/N77 ), .CLK(clk), 
        .CLRB(n888), .SETB(1'b1), .Q(n177) );
  dffascs1 \MEMinst/RF_data_in_reg[21]  ( .DIN(\MEMinst/N78 ), .CLK(clk), 
        .CLRB(n824), .SETB(1'b1), .Q(n175) );
  dffascs1 \MEMinst/RF_data_in_reg[22]  ( .DIN(\MEMinst/N79 ), .CLK(clk), 
        .CLRB(n883), .SETB(1'b1), .Q(n173) );
  dffascs1 \MEMinst/RF_data_in_reg[23]  ( .DIN(\MEMinst/N80 ), .CLK(clk), 
        .CLRB(n891), .SETB(1'b1), .Q(n171) );
  dffascs1 \MEMinst/RF_data_in_reg[24]  ( .DIN(\MEMinst/N81 ), .CLK(clk), 
        .CLRB(n906), .SETB(1'b1), .Q(n169) );
  dffascs1 \MEMinst/RF_data_in_reg[25]  ( .DIN(\MEMinst/N82 ), .CLK(clk), 
        .CLRB(n902), .SETB(1'b1), .Q(n167) );
  dffascs1 \MEMinst/RF_data_in_reg[26]  ( .DIN(\MEMinst/N83 ), .CLK(clk), 
        .CLRB(n913), .SETB(1'b1), .Q(n165) );
  dffascs1 \MEMinst/RF_data_in_reg[27]  ( .DIN(\MEMinst/N84 ), .CLK(clk), 
        .CLRB(n910), .SETB(1'b1), .Q(n163) );
  dffascs1 \MEMinst/RF_data_in_reg[28]  ( .DIN(\MEMinst/N85 ), .CLK(clk), 
        .CLRB(n922), .SETB(1'b1), .Q(n161) );
  dffascs1 \MEMinst/RF_data_in_reg[29]  ( .DIN(\MEMinst/N86 ), .CLK(clk), 
        .CLRB(n962), .SETB(1'b1), .Q(n159) );
  dffascs1 \MEMinst/RF_data_in_reg[30]  ( .DIN(\MEMinst/N87 ), .CLK(clk), 
        .CLRB(n963), .SETB(1'b1), .Q(n157) );
  dffascs1 \MEMinst/RF_data_in_reg[31]  ( .DIN(\MEMinst/N88 ), .CLK(clk), 
        .CLRB(n963), .SETB(1'b1), .Q(n155) );
  and2s1 U1 ( .DIN1(n676), .DIN2(n4121), .Q(n5) );
  nnd2s1 U2 ( .DIN1(n7004), .DIN2(n8950), .Q(n72) );
  nnd2s1 U3 ( .DIN1(n7107), .DIN2(n7108), .Q(n73) );
  nnd2s1 U4 ( .DIN1(n9361), .DIN2(n7108), .Q(n74) );
  xnr2s1 U5 ( .DIN1(n632), .DIN2(n9477), .Q(n87) );
  xnr2s1 U6 ( .DIN1(n632), .DIN2(n9479), .Q(n88) );
  xnr2s1 U7 ( .DIN1(n632), .DIN2(n9481), .Q(n89) );
  xnr2s1 U8 ( .DIN1(n632), .DIN2(n9483), .Q(n90) );
  xnr2s1 U9 ( .DIN1(n632), .DIN2(n9485), .Q(n91) );
  or2s1 U10 ( .DIN1(n1662), .DIN2(n662), .Q(n118) );
  or2s1 U11 ( .DIN1(n7059), .DIN2(n528), .Q(n127) );
  or2s1 U12 ( .DIN1(n528), .DIN2(stall), .Q(n128) );
  or2s1 U13 ( .DIN1(n1918), .DIN2(n441), .Q(n130) );
  or2s1 U14 ( .DIN1(n4535), .DIN2(n382), .Q(n131) );
  and2s1 U15 ( .DIN1(n5258), .DIN2(n5259), .Q(n138) );
  and2s1 U16 ( .DIN1(n5091), .DIN2(n5092), .Q(n139) );
  or2s1 U17 ( .DIN1(n5490), .DIN2(n438), .Q(n140) );
  or2s1 U18 ( .DIN1(n32), .DIN2(n438), .Q(n202) );
  or2s1 U19 ( .DIN1(n801), .DIN2(n742), .Q(n208) );
  or2s1 U20 ( .DIN1(n803), .DIN2(n4845), .Q(n210) );
  or2s1 U21 ( .DIN1(n1), .DIN2(n714), .Q(n211) );
  or2s1 U22 ( .DIN1(n4840), .DIN2(n747), .Q(n212) );
  or2s1 U23 ( .DIN1(n711), .DIN2(n439), .Q(n213) );
  or2s1 U24 ( .DIN1(n382), .DIN2(n4164), .Q(n214) );
  xnr2s1 U25 ( .DIN1(n430), .DIN2(n440), .Q(n216) );
  and2s1 U26 ( .DIN1(n3035), .DIN2(n3036), .Q(n217) );
  and2s1 U27 ( .DIN1(n3035), .DIN2(n3102), .Q(n218) );
  and2s1 U28 ( .DIN1(n3035), .DIN2(n3168), .Q(n219) );
  and2s1 U29 ( .DIN1(n3035), .DIN2(n3233), .Q(n220) );
  and2s1 U30 ( .DIN1(n3035), .DIN2(n3298), .Q(n221) );
  and2s1 U31 ( .DIN1(n3035), .DIN2(n3363), .Q(n222) );
  and2s1 U32 ( .DIN1(n3035), .DIN2(n3428), .Q(n223) );
  and2s1 U33 ( .DIN1(n3035), .DIN2(n3493), .Q(n224) );
  and4s1 U34 ( .DIN1(n5237), .DIN2(n5238), .DIN3(reg_write_MEM), .DIN4(n5239), 
        .Q(n226) );
  and2s1 U35 ( .DIN1(n9459), .DIN2(n1888), .Q(n328) );
  and2s1 U36 ( .DIN1(n4148), .DIN2(n5274), .Q(n329) );
  and2s1 U37 ( .DIN1(n4049), .DIN2(n1383), .Q(n338) );
  and2s1 U38 ( .DIN1(n4049), .DIN2(n4028), .Q(n339) );
  and2s1 U39 ( .DIN1(n4049), .DIN2(n4031), .Q(n340) );
  and2s1 U40 ( .DIN1(n4049), .DIN2(n4034), .Q(n341) );
  and2s1 U41 ( .DIN1(n4049), .DIN2(n4037), .Q(n342) );
  and2s1 U42 ( .DIN1(n4049), .DIN2(n4040), .Q(n343) );
  and2s1 U43 ( .DIN1(n4049), .DIN2(n4043), .Q(n344) );
  and2s1 U44 ( .DIN1(n4049), .DIN2(n4046), .Q(n345) );
  and2s1 U45 ( .DIN1(n4025), .DIN2(n1383), .Q(n346) );
  and2s1 U46 ( .DIN1(n4025), .DIN2(n4028), .Q(n347) );
  and2s1 U47 ( .DIN1(n4025), .DIN2(n4031), .Q(n348) );
  and2s1 U48 ( .DIN1(n4025), .DIN2(n4034), .Q(n349) );
  and2s1 U49 ( .DIN1(n4025), .DIN2(n4037), .Q(n350) );
  and2s1 U50 ( .DIN1(n4025), .DIN2(n4040), .Q(n351) );
  and2s1 U51 ( .DIN1(n4025), .DIN2(n4043), .Q(n352) );
  and2s1 U52 ( .DIN1(n4025), .DIN2(n4046), .Q(n353) );
  and2s1 U53 ( .DIN1(n4066), .DIN2(n1383), .Q(n354) );
  and2s1 U54 ( .DIN1(n4066), .DIN2(n4028), .Q(n355) );
  and2s1 U55 ( .DIN1(n4066), .DIN2(n4031), .Q(n356) );
  and2s1 U56 ( .DIN1(n4066), .DIN2(n4034), .Q(n357) );
  and2s1 U57 ( .DIN1(n4066), .DIN2(n4037), .Q(n358) );
  and2s1 U58 ( .DIN1(n4066), .DIN2(n4040), .Q(n359) );
  and2s1 U59 ( .DIN1(n4066), .DIN2(n4043), .Q(n360) );
  and2s1 U60 ( .DIN1(n4066), .DIN2(n4046), .Q(n361) );
  and2s1 U61 ( .DIN1(n4083), .DIN2(n1383), .Q(n362) );
  and2s1 U62 ( .DIN1(n4028), .DIN2(n4083), .Q(n363) );
  and2s1 U63 ( .DIN1(n4031), .DIN2(n4083), .Q(n364) );
  and2s1 U64 ( .DIN1(n4034), .DIN2(n4083), .Q(n365) );
  and2s1 U65 ( .DIN1(n4037), .DIN2(n4083), .Q(n366) );
  and2s1 U66 ( .DIN1(n4040), .DIN2(n4083), .Q(n367) );
  and2s1 U67 ( .DIN1(n4043), .DIN2(n4083), .Q(n368) );
  and2s1 U68 ( .DIN1(n4046), .DIN2(n4083), .Q(n369) );
  nnd4s1 U69 ( .DIN1(n5244), .DIN2(n5243), .DIN3(n1132), .DIN4(n1178), 
        .Q(n370) );
  nnd4s1 U70 ( .DIN1(n5244), .DIN2(n5243), .DIN3(n1180), .DIN4(n1122), 
        .Q(n371) );
  nnd3s1 U71 ( .DIN1(n4128), .DIN2(n130), .DIN3(n4148), .Q(n372) );
  nnd2s1 U72 ( .DIN1(n5073), .DIN2(n5074), .Q(n373) );
  hi1s1 U73 ( .DIN(n9211), .Q(n381) );
  hi1s1 U74 ( .DIN(n329), .Q(n382) );
  hi1s1 U75 ( .DIN(n329), .Q(n383) );
  hi1s1 U76 ( .DIN(n5404), .Q(n384) );
  hi1s1 U77 ( .DIN(n384), .Q(n385) );
  hi1s1 U78 ( .DIN(n74), .Q(n386) );
  hi1s1 U79 ( .DIN(n73), .Q(n387) );
  hi1s1 U80 ( .DIN(n87), .Q(n388) );
  hi1s1 U81 ( .DIN(n88), .Q(n389) );
  hi1s1 U82 ( .DIN(n89), .Q(n390) );
  hi1s1 U83 ( .DIN(n90), .Q(n391) );
  hi1s1 U84 ( .DIN(n91), .Q(n392) );
  xnr2s1 U85 ( .DIN1(n632), .DIN2(n739), .Q(n8466) );
  hi1s1 U86 ( .DIN(n8466), .Q(n393) );
  hi1s1 U87 ( .DIN(n8687), .Q(n394) );
  hi1s1 U88 ( .DIN(n394), .Q(n395) );
  hi1s1 U89 ( .DIN(n5), .Q(n396) );
  hi1s1 U90 ( .DIN(n5303), .Q(n397) );
  hi1s1 U91 ( .DIN(n5303), .Q(n398) );
  hi1s1 U92 ( .DIN(n1), .Q(n399) );
  hi1s1 U93 ( .DIN(n72), .Q(n400) );
  hi1s1 U94 ( .DIN(reg_out_A[31]), .Q(n401) );
  hi1s1 U95 ( .DIN(n127), .Q(n402) );
  hi1s1 U96 ( .DIN(n127), .Q(n403) );
  hi1s1 U97 ( .DIN(n127), .Q(n404) );
  hi1s1 U98 ( .DIN(n127), .Q(n405) );
  hi1s1 U99 ( .DIN(n79), .Q(n406) );
  hi1s1 U100 ( .DIN(n38), .Q(n407) );
  hi1s1 U101 ( .DIN(n83), .Q(n408) );
  hi1s1 U102 ( .DIN(n30), .Q(n409) );
  hi1s1 U103 ( .DIN(n68), .Q(n410) );
  hi1s1 U104 ( .DIN(n67), .Q(n411) );
  hi1s1 U105 ( .DIN(n78), .Q(n412) );
  hi1s1 U106 ( .DIN(n69), .Q(n413) );
  hi1s1 U107 ( .DIN(n37), .Q(n414) );
  hi1s1 U108 ( .DIN(n70), .Q(n415) );
  hi1s1 U109 ( .DIN(n82), .Q(n416) );
  hi1s1 U110 ( .DIN(n71), .Q(n417) );
  hi1s1 U111 ( .DIN(n85), .Q(n418) );
  hi1s1 U112 ( .DIN(n31), .Q(n419) );
  hi1s1 U113 ( .DIN(n86), .Q(n420) );
  hi1s1 U114 ( .DIN(n64), .Q(n421) );
  hi1s1 U115 ( .DIN(n84), .Q(n422) );
  hi1s1 U116 ( .DIN(n65), .Q(n423) );
  hi1s1 U117 ( .DIN(n66), .Q(n424) );
  hi1s1 U118 ( .DIN(n332), .Q(n425) );
  hi1s1 U119 ( .DIN(n80), .Q(n426) );
  hi1s1 U120 ( .DIN(n333), .Q(n427) );
  hi1s1 U121 ( .DIN(n81), .Q(n428) );
  hi1s1 U122 ( .DIN(n63), .Q(n429) );
  hi1s1 U123 ( .DIN(n331), .Q(n430) );
  hi1s1 U124 ( .DIN(n77), .Q(n431) );
  hi1s1 U125 ( .DIN(n330), .Q(n432) );
  hi1s1 U126 ( .DIN(n334), .Q(n433) );
  hi1s1 U127 ( .DIN(n335), .Q(n434) );
  hi1s1 U128 ( .DIN(n336), .Q(n435) );
  hi1s1 U129 ( .DIN(n372), .Q(n436) );
  hi1s1 U130 ( .DIN(n372), .Q(n437) );
  hi1s1 U131 ( .DIN(n337), .Q(n438) );
  hi1s1 U132 ( .DIN(n9489), .Q(n439) );
  hi1s1 U133 ( .DIN(n9489), .Q(n440) );
  hi1s1 U134 ( .DIN(n382), .Q(n441) );
  hi1s1 U135 ( .DIN(n328), .Q(n442) );
  hi1s1 U136 ( .DIN(n328), .Q(n443) );
  hi1s1 U137 ( .DIN(n217), .Q(n444) );
  hi1s1 U138 ( .DIN(n217), .Q(n445) );
  hi1s1 U139 ( .DIN(n218), .Q(n446) );
  hi1s1 U140 ( .DIN(n218), .Q(n447) );
  hi1s1 U141 ( .DIN(n219), .Q(n448) );
  hi1s1 U142 ( .DIN(n219), .Q(n449) );
  hi1s1 U143 ( .DIN(n220), .Q(n450) );
  hi1s1 U144 ( .DIN(n220), .Q(n451) );
  hi1s1 U145 ( .DIN(n221), .Q(n452) );
  hi1s1 U146 ( .DIN(n221), .Q(n453) );
  hi1s1 U147 ( .DIN(n222), .Q(n454) );
  hi1s1 U148 ( .DIN(n222), .Q(n455) );
  hi1s1 U149 ( .DIN(n223), .Q(n456) );
  hi1s1 U150 ( .DIN(n223), .Q(n457) );
  hi1s1 U151 ( .DIN(n224), .Q(n458) );
  hi1s1 U152 ( .DIN(n224), .Q(n459) );
  hi1s1 U153 ( .DIN(n368), .Q(n460) );
  hi1s1 U154 ( .DIN(n368), .Q(n461) );
  hi1s1 U155 ( .DIN(n369), .Q(n462) );
  hi1s1 U156 ( .DIN(n369), .Q(n463) );
  hi1s1 U157 ( .DIN(n366), .Q(n464) );
  hi1s1 U158 ( .DIN(n366), .Q(n465) );
  hi1s1 U159 ( .DIN(n367), .Q(n466) );
  hi1s1 U160 ( .DIN(n367), .Q(n467) );
  hi1s1 U161 ( .DIN(n364), .Q(n468) );
  hi1s1 U162 ( .DIN(n364), .Q(n469) );
  hi1s1 U163 ( .DIN(n365), .Q(n470) );
  hi1s1 U164 ( .DIN(n365), .Q(n471) );
  hi1s1 U165 ( .DIN(n362), .Q(n472) );
  hi1s1 U166 ( .DIN(n362), .Q(n473) );
  hi1s1 U167 ( .DIN(n363), .Q(n474) );
  hi1s1 U168 ( .DIN(n363), .Q(n475) );
  hi1s1 U169 ( .DIN(n338), .Q(n476) );
  hi1s1 U170 ( .DIN(n338), .Q(n477) );
  hi1s1 U171 ( .DIN(n354), .Q(n478) );
  hi1s1 U172 ( .DIN(n354), .Q(n479) );
  hi1s1 U173 ( .DIN(n361), .Q(n480) );
  hi1s1 U174 ( .DIN(n361), .Q(n481) );
  hi1s1 U175 ( .DIN(n346), .Q(n482) );
  hi1s1 U176 ( .DIN(n346), .Q(n483) );
  hi1s1 U177 ( .DIN(n353), .Q(n484) );
  hi1s1 U178 ( .DIN(n353), .Q(n485) );
  hi1s1 U179 ( .DIN(n345), .Q(n486) );
  hi1s1 U180 ( .DIN(n345), .Q(n487) );
  hi1s1 U181 ( .DIN(n357), .Q(n488) );
  hi1s1 U182 ( .DIN(n357), .Q(n489) );
  hi1s1 U183 ( .DIN(n359), .Q(n490) );
  hi1s1 U184 ( .DIN(n359), .Q(n491) );
  hi1s1 U185 ( .DIN(n343), .Q(n492) );
  hi1s1 U186 ( .DIN(n343), .Q(n493) );
  hi1s1 U187 ( .DIN(n355), .Q(n494) );
  hi1s1 U188 ( .DIN(n355), .Q(n495) );
  hi1s1 U189 ( .DIN(n339), .Q(n496) );
  hi1s1 U190 ( .DIN(n339), .Q(n497) );
  hi1s1 U191 ( .DIN(n341), .Q(n498) );
  hi1s1 U192 ( .DIN(n341), .Q(n499) );
  hi1s1 U193 ( .DIN(n349), .Q(n500) );
  hi1s1 U194 ( .DIN(n349), .Q(n501) );
  hi1s1 U195 ( .DIN(n351), .Q(n502) );
  hi1s1 U196 ( .DIN(n351), .Q(n503) );
  hi1s1 U197 ( .DIN(n360), .Q(n504) );
  hi1s1 U198 ( .DIN(n360), .Q(n505) );
  hi1s1 U199 ( .DIN(n347), .Q(n506) );
  hi1s1 U200 ( .DIN(n347), .Q(n507) );
  hi1s1 U201 ( .DIN(n356), .Q(n508) );
  hi1s1 U202 ( .DIN(n356), .Q(n509) );
  hi1s1 U203 ( .DIN(n358), .Q(n510) );
  hi1s1 U204 ( .DIN(n358), .Q(n511) );
  hi1s1 U205 ( .DIN(n342), .Q(n512) );
  hi1s1 U206 ( .DIN(n342), .Q(n513) );
  hi1s1 U207 ( .DIN(n344), .Q(n514) );
  hi1s1 U208 ( .DIN(n344), .Q(n515) );
  hi1s1 U209 ( .DIN(n352), .Q(n516) );
  hi1s1 U210 ( .DIN(n352), .Q(n517) );
  hi1s1 U211 ( .DIN(n340), .Q(n518) );
  hi1s1 U212 ( .DIN(n340), .Q(n519) );
  hi1s1 U213 ( .DIN(n348), .Q(n520) );
  hi1s1 U214 ( .DIN(n348), .Q(n521) );
  hi1s1 U215 ( .DIN(n350), .Q(n522) );
  hi1s1 U216 ( .DIN(n350), .Q(n523) );
  hi1s1 U217 ( .DIN(n226), .Q(n524) );
  hi1s1 U218 ( .DIN(n226), .Q(n525) );
  hi1s1 U219 ( .DIN(n374), .Q(n526) );
  hi1s1 U220 ( .DIN(n9453), .Q(n527) );
  hi1s1 U221 ( .DIN(n9453), .Q(n528) );
  hi1s1 U222 ( .DIN(n214), .Q(n529) );
  hi1s1 U223 ( .DIN(n214), .Q(n530) );
  hi1s1 U224 ( .DIN(n211), .Q(n531) );
  hi1s1 U225 ( .DIN(n211), .Q(n532) );
  hi1s1 U226 ( .DIN(\IDinst/N48 ), .Q(n533) );
  hi1s1 U227 ( .DIN(n533), .Q(n534) );
  hi1s1 U228 ( .DIN(n533), .Q(n535) );
  hi1s1 U229 ( .DIN(n373), .Q(n536) );
  hi1s1 U230 ( .DIN(n373), .Q(n537) );
  hi1s1 U231 ( .DIN(\IDinst/N43 ), .Q(n538) );
  hi1s1 U232 ( .DIN(n538), .Q(n539) );
  hi1s1 U233 ( .DIN(n370), .Q(n540) );
  hi1s1 U234 ( .DIN(n370), .Q(n541) );
  hi1s1 U235 ( .DIN(n371), .Q(n542) );
  hi1s1 U236 ( .DIN(n371), .Q(n543) );
  hi1s1 U237 ( .DIN(n212), .Q(n544) );
  hi1s1 U238 ( .DIN(n212), .Q(n545) );
  hi1s1 U239 ( .DIN(n208), .Q(n546) );
  hi1s1 U240 ( .DIN(n208), .Q(n547) );
  hi1s1 U241 ( .DIN(n7041), .Q(n548) );
  hi1s1 U242 ( .DIN(n7041), .Q(n549) );
  hi1s1 U243 ( .DIN(n48), .Q(n550) );
  hi1s1 U244 ( .DIN(n48), .Q(n551) );
  hi1s1 U245 ( .DIN(n213), .Q(n552) );
  hi1s1 U246 ( .DIN(n213), .Q(n553) );
  hi1s1 U247 ( .DIN(n210), .Q(n554) );
  hi1s1 U248 ( .DIN(n210), .Q(n555) );
  hi1s1 U249 ( .DIN(n465), .Q(n556) );
  hi1s1 U250 ( .DIN(n464), .Q(n557) );
  hi1s1 U251 ( .DIN(n467), .Q(n558) );
  hi1s1 U252 ( .DIN(n466), .Q(n559) );
  hi1s1 U253 ( .DIN(n461), .Q(n560) );
  hi1s1 U254 ( .DIN(n460), .Q(n561) );
  hi1s1 U255 ( .DIN(n463), .Q(n562) );
  hi1s1 U256 ( .DIN(n462), .Q(n563) );
  hi1s1 U257 ( .DIN(n473), .Q(n564) );
  hi1s1 U258 ( .DIN(n472), .Q(n565) );
  hi1s1 U259 ( .DIN(n475), .Q(n566) );
  hi1s1 U260 ( .DIN(n474), .Q(n567) );
  hi1s1 U261 ( .DIN(n469), .Q(n568) );
  hi1s1 U262 ( .DIN(n468), .Q(n569) );
  hi1s1 U263 ( .DIN(n471), .Q(n570) );
  hi1s1 U264 ( .DIN(n470), .Q(n571) );
  hi1s1 U265 ( .DIN(n511), .Q(n572) );
  hi1s1 U266 ( .DIN(n510), .Q(n573) );
  hi1s1 U267 ( .DIN(n491), .Q(n574) );
  hi1s1 U268 ( .DIN(n490), .Q(n575) );
  hi1s1 U269 ( .DIN(n505), .Q(n576) );
  hi1s1 U270 ( .DIN(n504), .Q(n577) );
  hi1s1 U271 ( .DIN(n481), .Q(n578) );
  hi1s1 U272 ( .DIN(n480), .Q(n579) );
  hi1s1 U273 ( .DIN(n479), .Q(n580) );
  hi1s1 U274 ( .DIN(n478), .Q(n581) );
  hi1s1 U275 ( .DIN(n495), .Q(n582) );
  hi1s1 U276 ( .DIN(n494), .Q(n583) );
  hi1s1 U277 ( .DIN(n509), .Q(n584) );
  hi1s1 U278 ( .DIN(n508), .Q(n585) );
  hi1s1 U279 ( .DIN(n489), .Q(n586) );
  hi1s1 U280 ( .DIN(n488), .Q(n587) );
  hi1s1 U281 ( .DIN(n523), .Q(n588) );
  hi1s1 U282 ( .DIN(n522), .Q(n589) );
  hi1s1 U283 ( .DIN(n503), .Q(n590) );
  hi1s1 U284 ( .DIN(n502), .Q(n591) );
  hi1s1 U285 ( .DIN(n517), .Q(n592) );
  hi1s1 U286 ( .DIN(n516), .Q(n593) );
  hi1s1 U287 ( .DIN(n485), .Q(n594) );
  hi1s1 U288 ( .DIN(n484), .Q(n595) );
  hi1s1 U289 ( .DIN(n483), .Q(n596) );
  hi1s1 U290 ( .DIN(n482), .Q(n597) );
  hi1s1 U291 ( .DIN(n507), .Q(n598) );
  hi1s1 U292 ( .DIN(n506), .Q(n599) );
  hi1s1 U293 ( .DIN(n521), .Q(n600) );
  hi1s1 U294 ( .DIN(n520), .Q(n601) );
  hi1s1 U295 ( .DIN(n501), .Q(n602) );
  hi1s1 U296 ( .DIN(n500), .Q(n603) );
  hi1s1 U297 ( .DIN(n513), .Q(n604) );
  hi1s1 U298 ( .DIN(n512), .Q(n605) );
  hi1s1 U299 ( .DIN(n493), .Q(n606) );
  hi1s1 U300 ( .DIN(n492), .Q(n607) );
  hi1s1 U301 ( .DIN(n515), .Q(n608) );
  hi1s1 U302 ( .DIN(n514), .Q(n609) );
  hi1s1 U303 ( .DIN(n487), .Q(n610) );
  hi1s1 U304 ( .DIN(n486), .Q(n611) );
  hi1s1 U305 ( .DIN(n477), .Q(n612) );
  hi1s1 U306 ( .DIN(n476), .Q(n613) );
  hi1s1 U307 ( .DIN(n497), .Q(n614) );
  hi1s1 U308 ( .DIN(n496), .Q(n615) );
  hi1s1 U309 ( .DIN(n519), .Q(n616) );
  hi1s1 U310 ( .DIN(n518), .Q(n617) );
  hi1s1 U311 ( .DIN(n499), .Q(n618) );
  hi1s1 U312 ( .DIN(n498), .Q(n619) );
  hi1s1 U313 ( .DIN(n5375), .Q(n620) );
  hi1s1 U314 ( .DIN(n140), .Q(n621) );
  hi1s1 U315 ( .DIN(n140), .Q(n622) );
  hi1s1 U316 ( .DIN(n140), .Q(n623) );
  hi1s1 U317 ( .DIN(n1466), .Q(n624) );
  hi1s1 U318 ( .DIN(n1466), .Q(n625) );
  hi1s1 U319 ( .DIN(n525), .Q(n626) );
  hi1s1 U320 ( .DIN(n524), .Q(n627) );
  hi1s1 U321 ( .DIN(n202), .Q(n628) );
  hi1s1 U322 ( .DIN(n202), .Q(n629) );
  hi1s1 U323 ( .DIN(n202), .Q(n630) );
  hi1s1 U324 ( .DIN(n5423), .Q(n631) );
  hi1s1 U325 ( .DIN(n631), .Q(n632) );
  hi1s1 U326 ( .DIN(n631), .Q(n633) );
  hi1s1 U327 ( .DIN(\IDinst/N48 ), .Q(n634) );
  hi1s1 U328 ( .DIN(\IDinst/N43 ), .Q(n635) );
  hi1s1 U329 ( .DIN(\IDinst/N43 ), .Q(n636) );
  hi1s1 U330 ( .DIN(n131), .Q(n637) );
  hi1s1 U331 ( .DIN(n131), .Q(n638) );
  hi1s1 U332 ( .DIN(n131), .Q(n639) );
  hi1s1 U333 ( .DIN(n131), .Q(n640) );
  hi1s1 U334 ( .DIN(n138), .Q(n641) );
  hi1s1 U335 ( .DIN(n138), .Q(n642) );
  hi1s1 U336 ( .DIN(n138), .Q(n643) );
  hi1s1 U337 ( .DIN(n138), .Q(n644) );
  hi1s1 U338 ( .DIN(n624), .Q(n645) );
  hi1s1 U339 ( .DIN(n625), .Q(n646) );
  hi1s1 U340 ( .DIN(n624), .Q(n647) );
  hi1s1 U341 ( .DIN(n625), .Q(n648) );
  hi1s1 U342 ( .DIN(n130), .Q(n649) );
  hi1s1 U343 ( .DIN(n130), .Q(n650) );
  hi1s1 U344 ( .DIN(n130), .Q(n651) );
  hi1s1 U345 ( .DIN(n130), .Q(n652) );
  hi1s1 U346 ( .DIN(n5381), .Q(n653) );
  hi1s1 U347 ( .DIN(n5381), .Q(n654) );
  hi1s1 U348 ( .DIN(n5381), .Q(n655) );
  hi1s1 U349 ( .DIN(n5381), .Q(n656) );
  hi1s1 U350 ( .DIN(n118), .Q(n657) );
  hi1s1 U351 ( .DIN(n118), .Q(n658) );
  hi1s1 U352 ( .DIN(n118), .Q(n659) );
  hi1s1 U353 ( .DIN(n118), .Q(n660) );
  hi1s1 U354 ( .DIN(n128), .Q(n661) );
  hi1s1 U355 ( .DIN(n128), .Q(n662) );
  hi1s1 U356 ( .DIN(n128), .Q(n663) );
  hi1s1 U357 ( .DIN(n128), .Q(n664) );
  hi1s1 U358 ( .DIN(n139), .Q(n665) );
  hi1s1 U359 ( .DIN(n139), .Q(n666) );
  hi1s1 U360 ( .DIN(n139), .Q(n667) );
  hi1s1 U361 ( .DIN(n139), .Q(n668) );
  hi1s1 U362 ( .DIN(n138), .Q(n669) );
  hi1s1 U363 ( .DIN(n669), .Q(n670) );
  hi1s1 U364 ( .DIN(n669), .Q(n671) );
  hi1s1 U365 ( .DIN(n669), .Q(n672) );
  hi1s1 U366 ( .DIN(n669), .Q(n673) );
  hi1s1 U367 ( .DIN(n131), .Q(n674) );
  hi1s1 U368 ( .DIN(n674), .Q(n675) );
  hi1s1 U369 ( .DIN(n674), .Q(n676) );
  hi1s1 U370 ( .DIN(n674), .Q(n677) );
  hi1s1 U371 ( .DIN(n674), .Q(n678) );
  hi1s1 U372 ( .DIN(n139), .Q(n679) );
  hi1s1 U373 ( .DIN(n679), .Q(n680) );
  hi1s1 U374 ( .DIN(n679), .Q(n681) );
  hi1s1 U375 ( .DIN(n679), .Q(n682) );
  hi1s1 U376 ( .DIN(n679), .Q(n683) );
  hi1s1 U377 ( .DIN(n662), .Q(n684) );
  hi1s1 U378 ( .DIN(n663), .Q(n685) );
  hi1s1 U379 ( .DIN(n661), .Q(n686) );
  hi1s1 U380 ( .DIN(n662), .Q(n687) );
  hi1s1 U381 ( .DIN(n3496), .Q(n688) );
  hi1s1 U382 ( .DIN(n688), .Q(n689) );
  hi1s1 U383 ( .DIN(n3562), .Q(n690) );
  hi1s1 U384 ( .DIN(n690), .Q(n691) );
  hi1s1 U385 ( .DIN(n2509), .Q(n692) );
  hi1s1 U386 ( .DIN(n692), .Q(n693) );
  hi1s1 U387 ( .DIN(n3628), .Q(n694) );
  hi1s1 U388 ( .DIN(n694), .Q(n695) );
  hi1s1 U389 ( .DIN(n2577), .Q(n696) );
  hi1s1 U390 ( .DIN(n696), .Q(n697) );
  hi1s1 U391 ( .DIN(n3694), .Q(n698) );
  hi1s1 U392 ( .DIN(n698), .Q(n699) );
  nb1s1 U393 ( .DIN(n5306), .Q(n700) );
  hi1s1 U394 ( .DIN(n2643), .Q(n701) );
  hi1s1 U395 ( .DIN(n701), .Q(n702) );
  hi1s1 U396 ( .DIN(n3760), .Q(n703) );
  hi1s1 U397 ( .DIN(n703), .Q(n704) );
  hi1s1 U398 ( .DIN(n5375), .Q(n705) );
  hi1s1 U399 ( .DIN(n705), .Q(n706) );
  hi1s1 U400 ( .DIN(n9488), .Q(n707) );
  nnd2s1 U401 ( .DIN1(n2572), .DIN2(n2772), .Q(n708) );
  hi1s1 U402 ( .DIN(n3826), .Q(n709) );
  hi1s1 U403 ( .DIN(n709), .Q(n710) );
  hi1s1 U404 ( .DIN(n711), .Q(n712) );
  xor2s1 U405 ( .DIN1(\IDinst/n1403 ), .DIN2(n634), .Q(n5079) );
  hi1s1 U406 ( .DIN(n5079), .Q(n713) );
  hi1s1 U407 ( .DIN(n714), .Q(n715) );
  nb1s1 U408 ( .DIN(reg_out_B[5]), .Q(n716) );
  hi1s1 U409 ( .DIN(n717), .Q(n718) );
  and2s1 U410 ( .DIN1(n5949), .DIN2(n792), .Q(n719) );
  hi1s1 U411 ( .DIN(n5359), .Q(n720) );
  nnd2s1 U412 ( .DIN1(n2572), .DIN2(n2838), .Q(n721) );
  nnd4s1 U413 ( .DIN1(n9032), .DIN2(n9033), .DIN3(n9034), .DIN4(n788), 
        .Q(n722) );
  hi1s1 U414 ( .DIN(n5368), .Q(n723) );
  nnd2s1 U415 ( .DIN1(n3035), .DIN2(n3955), .Q(n724) );
  hi1s1 U416 ( .DIN(n5826), .Q(n725) );
  hi1s1 U417 ( .DIN(n725), .Q(n726) );
  nor2s1 U418 ( .DIN1(n9213), .DIN2(n9214), .Q(n727) );
  xor2s1 U419 ( .DIN1(n9419), .DIN2(n635), .Q(n4933) );
  hi1s1 U420 ( .DIN(n4933), .Q(n728) );
  xor2s1 U421 ( .DIN1(\IDinst/n1430 ), .DIN2(n682), .Q(n5076) );
  hi1s1 U422 ( .DIN(n5076), .Q(n729) );
  nb1s1 U423 ( .DIN(n7339), .Q(n730) );
  nnd2s1 U424 ( .DIN1(n1428), .DIN2(n1429), .Q(n1394) );
  hi1s1 U425 ( .DIN(n1394), .Q(n731) );
  hi1s1 U426 ( .DIN(n4555), .Q(n732) );
  nb1s1 U427 ( .DIN(n9486), .Q(n733) );
  hi1s1 U428 ( .DIN(n62), .Q(n734) );
  hi1s1 U429 ( .DIN(n735), .Q(n736) );
  nnd2s1 U430 ( .DIN1(n2572), .DIN2(n2904), .Q(n737) );
  nnd2s1 U431 ( .DIN1(n3035), .DIN2(n4021), .Q(n738) );
  hi1s1 U432 ( .DIN(n206), .Q(n739) );
  hi1s1 U433 ( .DIN(n206), .Q(n740) );
  hi1s1 U434 ( .DIN(n205), .Q(n741) );
  hi1s1 U435 ( .DIN(n205), .Q(n742) );
  nnd2s1 U436 ( .DIN1(n5426), .DIN2(n9212), .Q(n743) );
  nb1s1 U437 ( .DIN(n5413), .Q(n744) );
  nb1s1 U438 ( .DIN(n5413), .Q(n745) );
  hi1s1 U439 ( .DIN(n207), .Q(n746) );
  hi1s1 U440 ( .DIN(n207), .Q(n747) );
  nor2s1 U441 ( .DIN1(n5075), .DIN2(n5244), .Q(n748) );
  nnd3s1 U442 ( .DIN1(n9458), .DIN2(n2), .DIN3(n9234), .Q(n749) );
  or2s1 U443 ( .DIN1(n778), .DIN2(n4157), .Q(n4284) );
  hi1s1 U444 ( .DIN(n4284), .Q(n750) );
  hi1s1 U445 ( .DIN(n4284), .Q(n751) );
  hi1s1 U446 ( .DIN(n204), .Q(n752) );
  hi1s1 U447 ( .DIN(n204), .Q(n753) );
  or2s1 U448 ( .DIN1(n399), .DIN2(n715), .Q(n5353) );
  hi1s1 U449 ( .DIN(n5353), .Q(n754) );
  hi1s1 U450 ( .DIN(n5353), .Q(n755) );
  nnd2s1 U451 ( .DIN1(n4149), .DIN2(n4534), .Q(n4285) );
  hi1s1 U452 ( .DIN(n4285), .Q(n756) );
  hi1s1 U453 ( .DIN(n4285), .Q(n757) );
  or2s1 U454 ( .DIN1(n9489), .DIN2(n712), .Q(n5313) );
  hi1s1 U455 ( .DIN(n5313), .Q(n758) );
  hi1s1 U456 ( .DIN(n5313), .Q(n759) );
  xor2s1 U457 ( .DIN1(\IDinst/n1403 ), .DIN2(n636), .Q(n5240) );
  hi1s1 U458 ( .DIN(n5240), .Q(n761) );
  xor2s1 U459 ( .DIN1(n9419), .DIN2(n533), .Q(n4941) );
  hi1s1 U460 ( .DIN(n4941), .Q(n762) );
  hi1s1 U461 ( .DIN(n7202), .Q(n763) );
  nnd2s1 U462 ( .DIN1(n1425), .DIN2(n1426), .Q(n1393) );
  hi1s1 U463 ( .DIN(n1393), .Q(n764) );
  nnd2s1 U464 ( .DIN1(n2572), .DIN2(n2970), .Q(n765) );
  nnd2s1 U465 ( .DIN1(n3035), .DIN2(n4098), .Q(n766) );
  and2s1 U466 ( .DIN1(n9232), .DIN2(n723), .Q(n5469) );
  hi1s1 U467 ( .DIN(n5469), .Q(n767) );
  hi1s1 U468 ( .DIN(n5469), .Q(n768) );
  nor2s1 U469 ( .DIN1(n9218), .DIN2(n9244), .Q(n769) );
  nor2s1 U470 ( .DIN1(n5073), .DIN2(n5075), .Q(n770) );
  or2s1 U471 ( .DIN1(n714), .DIN2(n399), .Q(n5351) );
  hi1s1 U472 ( .DIN(n5351), .Q(n771) );
  hi1s1 U473 ( .DIN(n5351), .Q(n772) );
  or2s1 U474 ( .DIN1(n1), .DIN2(n715), .Q(n5352) );
  hi1s1 U475 ( .DIN(n5352), .Q(n773) );
  hi1s1 U476 ( .DIN(n5352), .Q(n774) );
  nnd2s1 U477 ( .DIN1(n9234), .DIN2(n9237), .Q(n5338) );
  hi1s1 U478 ( .DIN(n5338), .Q(n775) );
  hi1s1 U479 ( .DIN(n5338), .Q(n776) );
  and2s1 U480 ( .DIN1(n329), .DIN2(n4712), .Q(n4149) );
  hi1s1 U481 ( .DIN(n4149), .Q(n777) );
  hi1s1 U482 ( .DIN(n4149), .Q(n778) );
  or2s1 U483 ( .DIN1(n624), .DIN2(n9383), .Q(n1794) );
  hi1s1 U484 ( .DIN(n1794), .Q(n779) );
  hi1s1 U485 ( .DIN(n1794), .Q(n780) );
  hi1s1 U486 ( .DIN(n4298), .Q(n781) );
  hi1s1 U487 ( .DIN(n8728), .Q(n782) );
  or2s1 U488 ( .DIN1(n440), .DIN2(n712), .Q(n5312) );
  hi1s1 U489 ( .DIN(n5312), .Q(n783) );
  hi1s1 U490 ( .DIN(n5312), .Q(n784) );
  nnd2s1 U491 ( .DIN1(n9036), .DIN2(n4878), .Q(n785) );
  nnd2s1 U492 ( .DIN1(n9036), .DIN2(n4878), .Q(n786) );
  nnd2s1 U493 ( .DIN1(n9036), .DIN2(n4878), .Q(n787) );
  nnd2s1 U494 ( .DIN1(n9036), .DIN2(n4878), .Q(n788) );
  or2s1 U495 ( .DIN1(n707), .DIN2(n9489), .Q(n5314) );
  hi1s1 U496 ( .DIN(n5314), .Q(n789) );
  hi1s1 U497 ( .DIN(n5314), .Q(n790) );
  hi1s1 U498 ( .DIN(n7040), .Q(n791) );
  hi1s1 U499 ( .DIN(n29), .Q(n792) );
  hi1s1 U500 ( .DIN(n9404), .Q(n793) );
  hi1s1 U501 ( .DIN(n9399), .Q(n794) );
  hi1s1 U502 ( .DIN(n9398), .Q(n795) );
  hi1s1 U503 ( .DIN(n9397), .Q(n796) );
  hi1s1 U504 ( .DIN(n9396), .Q(n797) );
  hi1s1 U505 ( .DIN(n9394), .Q(n798) );
  hi1s1 U506 ( .DIN(n9393), .Q(n799) );
  hi1s1 U507 ( .DIN(n9395), .Q(n800) );
  hi1s1 U508 ( .DIN(n61), .Q(n801) );
  nb1s1 U509 ( .DIN(n4840), .Q(n802) );
  nb1s1 U510 ( .DIN(n4840), .Q(n803) );
  hi1s1 U511 ( .DIN(n9459), .Q(n804) );
  hi1s1 U512 ( .DIN(n56), .Q(n805) );
  hi1s1 U513 ( .DIN(n56), .Q(n806) );
  hi1s1 U514 ( .DIN(n55), .Q(n807) );
  hi1s1 U515 ( .DIN(n55), .Q(n808) );
  nb1s1 U516 ( .DIN(n1001), .Q(n809) );
  nb1s1 U517 ( .DIN(n1001), .Q(n810) );
  nb1s1 U518 ( .DIN(n1024), .Q(n811) );
  nb1s1 U519 ( .DIN(n1000), .Q(n812) );
  nb1s1 U520 ( .DIN(n1000), .Q(n813) );
  nb1s1 U521 ( .DIN(n1000), .Q(n814) );
  nb1s1 U522 ( .DIN(n999), .Q(n815) );
  nb1s1 U523 ( .DIN(n999), .Q(n816) );
  nb1s1 U524 ( .DIN(n999), .Q(n817) );
  nb1s1 U525 ( .DIN(n998), .Q(n818) );
  nb1s1 U526 ( .DIN(n998), .Q(n819) );
  nb1s1 U527 ( .DIN(n998), .Q(n820) );
  nb1s1 U528 ( .DIN(n997), .Q(n821) );
  nb1s1 U529 ( .DIN(n997), .Q(n822) );
  nb1s1 U530 ( .DIN(n997), .Q(n823) );
  nb1s1 U531 ( .DIN(n996), .Q(n824) );
  nb1s1 U532 ( .DIN(n996), .Q(n825) );
  nb1s1 U533 ( .DIN(n996), .Q(n826) );
  nb1s1 U534 ( .DIN(n995), .Q(n827) );
  nb1s1 U535 ( .DIN(n995), .Q(n828) );
  nb1s1 U536 ( .DIN(n995), .Q(n829) );
  nb1s1 U537 ( .DIN(n1003), .Q(n830) );
  nb1s1 U538 ( .DIN(n1003), .Q(n831) );
  nb1s1 U539 ( .DIN(n1004), .Q(n832) );
  nb1s1 U540 ( .DIN(n994), .Q(n833) );
  nb1s1 U541 ( .DIN(n994), .Q(n834) );
  nb1s1 U542 ( .DIN(n994), .Q(n835) );
  nb1s1 U543 ( .DIN(n993), .Q(n836) );
  nb1s1 U544 ( .DIN(n993), .Q(n837) );
  nb1s1 U545 ( .DIN(n993), .Q(n838) );
  nb1s1 U546 ( .DIN(n992), .Q(n839) );
  nb1s1 U547 ( .DIN(n992), .Q(n840) );
  nb1s1 U548 ( .DIN(n992), .Q(n841) );
  nb1s1 U549 ( .DIN(n991), .Q(n842) );
  nb1s1 U550 ( .DIN(n991), .Q(n843) );
  nb1s1 U551 ( .DIN(n991), .Q(n844) );
  nb1s1 U552 ( .DIN(n1005), .Q(n845) );
  nb1s1 U553 ( .DIN(n1005), .Q(n846) );
  nb1s1 U554 ( .DIN(n994), .Q(n847) );
  nb1s1 U555 ( .DIN(n990), .Q(n848) );
  nb1s1 U556 ( .DIN(n990), .Q(n849) );
  nb1s1 U557 ( .DIN(n990), .Q(n850) );
  nb1s1 U558 ( .DIN(n989), .Q(n851) );
  nb1s1 U559 ( .DIN(n989), .Q(n852) );
  nb1s1 U560 ( .DIN(n989), .Q(n853) );
  nb1s1 U561 ( .DIN(n1006), .Q(n854) );
  nb1s1 U562 ( .DIN(n1006), .Q(n855) );
  nb1s1 U563 ( .DIN(n1023), .Q(n856) );
  nb1s1 U564 ( .DIN(n988), .Q(n857) );
  nb1s1 U565 ( .DIN(n988), .Q(n858) );
  nb1s1 U566 ( .DIN(n988), .Q(n859) );
  nb1s1 U567 ( .DIN(n987), .Q(n860) );
  nb1s1 U568 ( .DIN(n987), .Q(n861) );
  nb1s1 U569 ( .DIN(n987), .Q(n862) );
  nb1s1 U570 ( .DIN(n1007), .Q(n863) );
  nb1s1 U571 ( .DIN(n1007), .Q(n864) );
  nb1s1 U572 ( .DIN(n998), .Q(n865) );
  nb1s1 U573 ( .DIN(n986), .Q(n866) );
  nb1s1 U574 ( .DIN(n986), .Q(n867) );
  nb1s1 U575 ( .DIN(n986), .Q(n868) );
  nb1s1 U576 ( .DIN(n985), .Q(n869) );
  nb1s1 U577 ( .DIN(n985), .Q(n870) );
  nb1s1 U578 ( .DIN(n985), .Q(n871) );
  nb1s1 U579 ( .DIN(n984), .Q(n872) );
  nb1s1 U580 ( .DIN(n984), .Q(n873) );
  nb1s1 U581 ( .DIN(n984), .Q(n874) );
  nb1s1 U582 ( .DIN(n983), .Q(n875) );
  nb1s1 U583 ( .DIN(n983), .Q(n876) );
  nb1s1 U584 ( .DIN(n983), .Q(n877) );
  nb1s1 U585 ( .DIN(n1008), .Q(n878) );
  nb1s1 U586 ( .DIN(n1008), .Q(n879) );
  nb1s1 U587 ( .DIN(n1022), .Q(n880) );
  nb1s1 U588 ( .DIN(n982), .Q(n881) );
  nb1s1 U589 ( .DIN(n982), .Q(n882) );
  nb1s1 U590 ( .DIN(n982), .Q(n883) );
  nb1s1 U591 ( .DIN(n981), .Q(n884) );
  nb1s1 U592 ( .DIN(n981), .Q(n885) );
  nb1s1 U593 ( .DIN(n981), .Q(n886) );
  nb1s1 U594 ( .DIN(n1009), .Q(n887) );
  nb1s1 U595 ( .DIN(n1009), .Q(n888) );
  nb1s1 U596 ( .DIN(n996), .Q(n889) );
  nb1s1 U597 ( .DIN(n1010), .Q(n890) );
  nb1s1 U598 ( .DIN(n1010), .Q(n891) );
  nb1s1 U599 ( .DIN(n995), .Q(n892) );
  nb1s1 U600 ( .DIN(n980), .Q(n893) );
  nb1s1 U601 ( .DIN(n980), .Q(n894) );
  nb1s1 U602 ( .DIN(n980), .Q(n895) );
  nb1s1 U603 ( .DIN(n979), .Q(n896) );
  nb1s1 U604 ( .DIN(n979), .Q(n897) );
  nb1s1 U605 ( .DIN(n979), .Q(n898) );
  nb1s1 U606 ( .DIN(n978), .Q(n899) );
  nb1s1 U607 ( .DIN(n978), .Q(n900) );
  nb1s1 U608 ( .DIN(n978), .Q(n901) );
  nb1s1 U609 ( .DIN(n977), .Q(n902) );
  nb1s1 U610 ( .DIN(n977), .Q(n903) );
  nb1s1 U611 ( .DIN(n977), .Q(n904) );
  nb1s1 U612 ( .DIN(n1011), .Q(n905) );
  nb1s1 U613 ( .DIN(n1011), .Q(n906) );
  nb1s1 U614 ( .DIN(n1021), .Q(n907) );
  nb1s1 U615 ( .DIN(n976), .Q(n908) );
  nb1s1 U616 ( .DIN(n976), .Q(n909) );
  nb1s1 U617 ( .DIN(n976), .Q(n910) );
  nb1s1 U618 ( .DIN(n1012), .Q(n911) );
  nb1s1 U619 ( .DIN(n1012), .Q(n912) );
  nb1s1 U620 ( .DIN(n997), .Q(n913) );
  nb1s1 U621 ( .DIN(n975), .Q(n914) );
  nb1s1 U622 ( .DIN(n975), .Q(n915) );
  nb1s1 U623 ( .DIN(n975), .Q(n916) );
  nb1s1 U624 ( .DIN(n974), .Q(n917) );
  nb1s1 U625 ( .DIN(n974), .Q(n918) );
  nb1s1 U626 ( .DIN(n974), .Q(n919) );
  nb1s1 U627 ( .DIN(n973), .Q(n920) );
  nb1s1 U628 ( .DIN(n973), .Q(n921) );
  nb1s1 U629 ( .DIN(n973), .Q(n922) );
  nb1s1 U630 ( .DIN(n1013), .Q(n923) );
  nb1s1 U631 ( .DIN(n1013), .Q(n924) );
  nb1s1 U632 ( .DIN(n1002), .Q(n925) );
  nb1s1 U633 ( .DIN(n1014), .Q(n926) );
  nb1s1 U634 ( .DIN(n1014), .Q(n927) );
  nb1s1 U635 ( .DIN(n1020), .Q(n928) );
  nb1s1 U636 ( .DIN(n972), .Q(n929) );
  nb1s1 U637 ( .DIN(n972), .Q(n930) );
  nb1s1 U638 ( .DIN(n972), .Q(n931) );
  nb1s1 U639 ( .DIN(n971), .Q(n932) );
  nb1s1 U640 ( .DIN(n971), .Q(n933) );
  nb1s1 U641 ( .DIN(n971), .Q(n934) );
  nb1s1 U642 ( .DIN(n970), .Q(n935) );
  nb1s1 U643 ( .DIN(n970), .Q(n936) );
  nb1s1 U644 ( .DIN(n970), .Q(n937) );
  nb1s1 U645 ( .DIN(n969), .Q(n938) );
  nb1s1 U646 ( .DIN(n969), .Q(n939) );
  nb1s1 U647 ( .DIN(n969), .Q(n940) );
  nb1s1 U648 ( .DIN(n968), .Q(n941) );
  nb1s1 U649 ( .DIN(n968), .Q(n942) );
  nb1s1 U650 ( .DIN(n968), .Q(n943) );
  nb1s1 U651 ( .DIN(n967), .Q(n944) );
  nb1s1 U652 ( .DIN(n967), .Q(n945) );
  nb1s1 U653 ( .DIN(n967), .Q(n946) );
  nb1s1 U654 ( .DIN(n966), .Q(n947) );
  nb1s1 U655 ( .DIN(n966), .Q(n948) );
  nb1s1 U656 ( .DIN(n966), .Q(n949) );
  nb1s1 U657 ( .DIN(n1016), .Q(n950) );
  nb1s1 U658 ( .DIN(n1016), .Q(n951) );
  nb1s1 U659 ( .DIN(n1000), .Q(n952) );
  nb1s1 U660 ( .DIN(n965), .Q(n953) );
  nb1s1 U661 ( .DIN(n965), .Q(n954) );
  nb1s1 U662 ( .DIN(n965), .Q(n955) );
  nb1s1 U663 ( .DIN(n1017), .Q(n956) );
  nb1s1 U664 ( .DIN(n1017), .Q(n957) );
  nb1s1 U665 ( .DIN(n999), .Q(n958) );
  nb1s1 U666 ( .DIN(n964), .Q(n959) );
  nb1s1 U667 ( .DIN(n964), .Q(n960) );
  nb1s1 U668 ( .DIN(n964), .Q(n961) );
  nb1s1 U669 ( .DIN(n1018), .Q(n962) );
  nb1s1 U670 ( .DIN(n1018), .Q(n963) );
  nb1s1 U671 ( .DIN(n1017), .Q(n964) );
  nb1s1 U672 ( .DIN(n1017), .Q(n965) );
  nb1s1 U673 ( .DIN(n1016), .Q(n966) );
  nb1s1 U674 ( .DIN(n1016), .Q(n967) );
  nb1s1 U675 ( .DIN(n1015), .Q(n968) );
  nb1s1 U676 ( .DIN(n1015), .Q(n969) );
  nb1s1 U677 ( .DIN(n1015), .Q(n970) );
  nb1s1 U678 ( .DIN(n1014), .Q(n971) );
  nb1s1 U679 ( .DIN(n1014), .Q(n972) );
  nb1s1 U680 ( .DIN(n1013), .Q(n973) );
  nb1s1 U681 ( .DIN(n1013), .Q(n974) );
  nb1s1 U682 ( .DIN(n1012), .Q(n975) );
  nb1s1 U683 ( .DIN(n1012), .Q(n976) );
  nb1s1 U684 ( .DIN(n1011), .Q(n977) );
  nb1s1 U685 ( .DIN(n1011), .Q(n978) );
  nb1s1 U686 ( .DIN(n1010), .Q(n979) );
  nb1s1 U687 ( .DIN(n1010), .Q(n980) );
  nb1s1 U688 ( .DIN(n1009), .Q(n981) );
  nb1s1 U689 ( .DIN(n1009), .Q(n982) );
  nb1s1 U690 ( .DIN(n1008), .Q(n983) );
  nb1s1 U691 ( .DIN(n1008), .Q(n984) );
  nb1s1 U692 ( .DIN(n1007), .Q(n985) );
  nb1s1 U693 ( .DIN(n1007), .Q(n986) );
  nb1s1 U694 ( .DIN(n1006), .Q(n987) );
  nb1s1 U695 ( .DIN(n1006), .Q(n988) );
  nb1s1 U696 ( .DIN(n1005), .Q(n989) );
  nb1s1 U697 ( .DIN(n1005), .Q(n990) );
  nb1s1 U698 ( .DIN(n1004), .Q(n991) );
  nb1s1 U699 ( .DIN(n1004), .Q(n992) );
  nb1s1 U700 ( .DIN(n1004), .Q(n993) );
  nb1s1 U701 ( .DIN(n1003), .Q(n994) );
  nb1s1 U702 ( .DIN(n1003), .Q(n995) );
  nb1s1 U703 ( .DIN(n1002), .Q(n996) );
  nb1s1 U704 ( .DIN(n1002), .Q(n997) );
  nb1s1 U705 ( .DIN(n1002), .Q(n998) );
  nb1s1 U706 ( .DIN(n1001), .Q(n999) );
  nb1s1 U707 ( .DIN(n1001), .Q(n1000) );
  nb1s1 U708 ( .DIN(n1024), .Q(n1001) );
  nb1s1 U709 ( .DIN(n1024), .Q(n1002) );
  nb1s1 U710 ( .DIN(n1024), .Q(n1003) );
  nb1s1 U711 ( .DIN(n1023), .Q(n1004) );
  nb1s1 U712 ( .DIN(n1023), .Q(n1005) );
  nb1s1 U713 ( .DIN(n1023), .Q(n1006) );
  nb1s1 U714 ( .DIN(n1022), .Q(n1007) );
  nb1s1 U715 ( .DIN(n1022), .Q(n1008) );
  nb1s1 U716 ( .DIN(n1022), .Q(n1009) );
  nb1s1 U717 ( .DIN(n1021), .Q(n1010) );
  nb1s1 U718 ( .DIN(n1021), .Q(n1011) );
  nb1s1 U719 ( .DIN(n1021), .Q(n1012) );
  nb1s1 U720 ( .DIN(n1020), .Q(n1013) );
  nb1s1 U721 ( .DIN(n1020), .Q(n1014) );
  nb1s1 U722 ( .DIN(n1020), .Q(n1015) );
  nb1s1 U723 ( .DIN(n1019), .Q(n1016) );
  nb1s1 U724 ( .DIN(n1019), .Q(n1017) );
  nb1s1 U725 ( .DIN(n1019), .Q(n1018) );
  nb1s1 U726 ( .DIN(n9588), .Q(n1019) );
  nb1s1 U727 ( .DIN(n9588), .Q(n1020) );
  nb1s1 U728 ( .DIN(n9588), .Q(n1021) );
  nb1s1 U729 ( .DIN(n9588), .Q(n1022) );
  nb1s1 U730 ( .DIN(n9588), .Q(n1023) );
  nb1s1 U731 ( .DIN(n9588), .Q(n1024) );
  hi1s1 U732 ( .DIN(n1065), .Q(n1025) );
  hi1s1 U733 ( .DIN(n1122), .Q(n1026) );
  hi1s1 U734 ( .DIN(n1122), .Q(n1027) );
  hi1s1 U735 ( .DIN(n1123), .Q(n1028) );
  hi1s1 U736 ( .DIN(n1123), .Q(n1029) );
  hi1s1 U737 ( .DIN(n1123), .Q(n1030) );
  hi1s1 U738 ( .DIN(n1123), .Q(n1031) );
  hi1s1 U739 ( .DIN(n1123), .Q(n1032) );
  hi1s1 U740 ( .DIN(n1123), .Q(n1033) );
  hi1s1 U741 ( .DIN(n1123), .Q(n1034) );
  hi1s1 U742 ( .DIN(n1123), .Q(n1035) );
  hi1s1 U743 ( .DIN(n1123), .Q(n1036) );
  hi1s1 U744 ( .DIN(n1123), .Q(n1037) );
  hi1s1 U745 ( .DIN(n1124), .Q(n1038) );
  hi1s1 U746 ( .DIN(n1124), .Q(n1039) );
  hi1s1 U747 ( .DIN(n1124), .Q(n1040) );
  hi1s1 U748 ( .DIN(n1124), .Q(n1041) );
  hi1s1 U749 ( .DIN(n1124), .Q(n1042) );
  hi1s1 U750 ( .DIN(n1124), .Q(n1043) );
  hi1s1 U751 ( .DIN(n1124), .Q(n1044) );
  hi1s1 U752 ( .DIN(n1124), .Q(n1045) );
  hi1s1 U753 ( .DIN(n1124), .Q(n1046) );
  hi1s1 U754 ( .DIN(n1124), .Q(n1047) );
  hi1s1 U755 ( .DIN(n1125), .Q(n1048) );
  hi1s1 U756 ( .DIN(n1125), .Q(n1049) );
  hi1s1 U757 ( .DIN(n1125), .Q(n1050) );
  hi1s1 U758 ( .DIN(n1125), .Q(n1051) );
  hi1s1 U759 ( .DIN(n1125), .Q(n1052) );
  hi1s1 U760 ( .DIN(n1125), .Q(n1053) );
  hi1s1 U761 ( .DIN(n1125), .Q(n1054) );
  hi1s1 U762 ( .DIN(n1125), .Q(n1055) );
  hi1s1 U763 ( .DIN(n1125), .Q(n1056) );
  hi1s1 U764 ( .DIN(n1125), .Q(n1057) );
  hi1s1 U765 ( .DIN(n1096), .Q(n1058) );
  hi1s1 U766 ( .DIN(n1125), .Q(n1059) );
  hi1s1 U767 ( .DIN(n1124), .Q(n1060) );
  hi1s1 U768 ( .DIN(n1123), .Q(n1061) );
  hi1s1 U769 ( .DIN(\IDinst/N39 ), .Q(n1062) );
  hi1s1 U770 ( .DIN(\IDinst/N39 ), .Q(n1063) );
  hi1s1 U771 ( .DIN(\IDinst/N39 ), .Q(n1064) );
  hi1s1 U772 ( .DIN(n1130), .Q(n1065) );
  hi1s1 U773 ( .DIN(n1129), .Q(n1066) );
  hi1s1 U774 ( .DIN(n1132), .Q(n1067) );
  hi1s1 U775 ( .DIN(n1132), .Q(n1068) );
  hi1s1 U776 ( .DIN(n1132), .Q(n1069) );
  hi1s1 U777 ( .DIN(n1131), .Q(n1070) );
  hi1s1 U778 ( .DIN(n1131), .Q(n1071) );
  hi1s1 U779 ( .DIN(n1131), .Q(n1072) );
  hi1s1 U780 ( .DIN(n1130), .Q(n1073) );
  hi1s1 U781 ( .DIN(n1130), .Q(n1074) );
  hi1s1 U782 ( .DIN(n1130), .Q(n1075) );
  hi1s1 U783 ( .DIN(n1129), .Q(n1076) );
  hi1s1 U784 ( .DIN(n1129), .Q(n1077) );
  hi1s1 U785 ( .DIN(n1129), .Q(n1078) );
  hi1s1 U786 ( .DIN(n1131), .Q(n1079) );
  hi1s1 U787 ( .DIN(n1130), .Q(n1080) );
  hi1s1 U788 ( .DIN(n1129), .Q(n1081) );
  hi1s1 U789 ( .DIN(n1128), .Q(n1082) );
  hi1s1 U790 ( .DIN(n1128), .Q(n1083) );
  hi1s1 U791 ( .DIN(n1127), .Q(n1084) );
  hi1s1 U792 ( .DIN(n1128), .Q(n1085) );
  hi1s1 U793 ( .DIN(n1127), .Q(n1086) );
  hi1s1 U794 ( .DIN(n1128), .Q(n1087) );
  hi1s1 U795 ( .DIN(n1129), .Q(n1088) );
  hi1s1 U796 ( .DIN(n1132), .Q(n1089) );
  hi1s1 U797 ( .DIN(n1129), .Q(n1090) );
  hi1s1 U798 ( .DIN(n1127), .Q(n1091) );
  hi1s1 U799 ( .DIN(n1128), .Q(n1092) );
  hi1s1 U800 ( .DIN(n1126), .Q(n1093) );
  hi1s1 U801 ( .DIN(n1126), .Q(n1094) );
  hi1s1 U802 ( .DIN(n1130), .Q(n1095) );
  hi1s1 U803 ( .DIN(n1132), .Q(n1096) );
  hi1s1 U804 ( .DIN(n1128), .Q(n1097) );
  hi1s1 U805 ( .DIN(n1128), .Q(n1098) );
  hi1s1 U806 ( .DIN(n1128), .Q(n1099) );
  hi1s1 U807 ( .DIN(n1127), .Q(n1100) );
  hi1s1 U808 ( .DIN(n1127), .Q(n1101) );
  hi1s1 U809 ( .DIN(n1127), .Q(n1102) );
  hi1s1 U810 ( .DIN(n1129), .Q(n1103) );
  hi1s1 U811 ( .DIN(n1132), .Q(n1104) );
  hi1s1 U812 ( .DIN(n1131), .Q(n1105) );
  hi1s1 U813 ( .DIN(n1126), .Q(n1106) );
  hi1s1 U814 ( .DIN(n1126), .Q(n1107) );
  hi1s1 U815 ( .DIN(n1126), .Q(n1108) );
  hi1s1 U816 ( .DIN(n1127), .Q(n1109) );
  hi1s1 U817 ( .DIN(n1126), .Q(n1110) );
  hi1s1 U818 ( .DIN(n1126), .Q(n1111) );
  hi1s1 U819 ( .DIN(n1127), .Q(n1112) );
  hi1s1 U820 ( .DIN(n1131), .Q(n1113) );
  hi1s1 U821 ( .DIN(n1131), .Q(n1114) );
  hi1s1 U822 ( .DIN(n1126), .Q(n1115) );
  hi1s1 U823 ( .DIN(n1128), .Q(n1116) );
  hi1s1 U824 ( .DIN(n1127), .Q(n1117) );
  hi1s1 U825 ( .DIN(n1132), .Q(n1118) );
  hi1s1 U826 ( .DIN(n1131), .Q(n1119) );
  hi1s1 U827 ( .DIN(n1130), .Q(n1120) );
  hi1s1 U828 ( .DIN(n1130), .Q(n1121) );
  hi1s1 U829 ( .DIN(n1129), .Q(n1122) );
  hi1s1 U830 ( .DIN(n1130), .Q(n1123) );
  hi1s1 U831 ( .DIN(n1126), .Q(n1124) );
  hi1s1 U832 ( .DIN(n1132), .Q(n1125) );
  hi1s1 U833 ( .DIN(\IDinst/N39 ), .Q(n1126) );
  hi1s1 U834 ( .DIN(\IDinst/N39 ), .Q(n1127) );
  hi1s1 U835 ( .DIN(\IDinst/N39 ), .Q(n1128) );
  hi1s1 U836 ( .DIN(\IDinst/N39 ), .Q(n1129) );
  hi1s1 U837 ( .DIN(\IDinst/N39 ), .Q(n1130) );
  hi1s1 U838 ( .DIN(\IDinst/N39 ), .Q(n1131) );
  hi1s1 U839 ( .DIN(\IDinst/N39 ), .Q(n1132) );
  hi1s1 U840 ( .DIN(n1153), .Q(n1133) );
  hi1s1 U841 ( .DIN(n1178), .Q(n1134) );
  hi1s1 U842 ( .DIN(n1178), .Q(n1135) );
  hi1s1 U843 ( .DIN(n1178), .Q(n1136) );
  hi1s1 U844 ( .DIN(n1178), .Q(n1137) );
  hi1s1 U845 ( .DIN(n1178), .Q(n1138) );
  hi1s1 U846 ( .DIN(n1178), .Q(n1139) );
  hi1s1 U847 ( .DIN(n1178), .Q(n1140) );
  hi1s1 U848 ( .DIN(n1179), .Q(n1141) );
  hi1s1 U849 ( .DIN(n1179), .Q(n1142) );
  hi1s1 U850 ( .DIN(n1179), .Q(n1143) );
  hi1s1 U851 ( .DIN(n1179), .Q(n1144) );
  hi1s1 U852 ( .DIN(n1179), .Q(n1145) );
  hi1s1 U853 ( .DIN(n1179), .Q(n1146) );
  hi1s1 U854 ( .DIN(n1179), .Q(n1147) );
  hi1s1 U855 ( .DIN(n1179), .Q(n1148) );
  hi1s1 U856 ( .DIN(n1179), .Q(n1149) );
  hi1s1 U857 ( .DIN(n1179), .Q(n1150) );
  hi1s1 U858 ( .DIN(n1154), .Q(n1151) );
  hi1s1 U859 ( .DIN(n1179), .Q(n1152) );
  hi1s1 U860 ( .DIN(n1180), .Q(n1153) );
  hi1s1 U861 ( .DIN(n1180), .Q(n1154) );
  hi1s1 U862 ( .DIN(n1180), .Q(n1155) );
  hi1s1 U863 ( .DIN(n1180), .Q(n1156) );
  hi1s1 U864 ( .DIN(n1180), .Q(n1157) );
  hi1s1 U865 ( .DIN(n1151), .Q(n1158) );
  hi1s1 U866 ( .DIN(n1180), .Q(n1159) );
  hi1s1 U867 ( .DIN(n1180), .Q(n1160) );
  hi1s1 U868 ( .DIN(n1151), .Q(n1161) );
  hi1s1 U869 ( .DIN(n1150), .Q(n1162) );
  hi1s1 U870 ( .DIN(n1180), .Q(n1163) );
  hi1s1 U871 ( .DIN(n1180), .Q(n1164) );
  hi1s1 U872 ( .DIN(n1180), .Q(n1165) );
  hi1s1 U873 ( .DIN(n1180), .Q(n1166) );
  hi1s1 U874 ( .DIN(n1149), .Q(n1167) );
  hi1s1 U875 ( .DIN(n1180), .Q(n1168) );
  hi1s1 U876 ( .DIN(n1180), .Q(n1169) );
  hi1s1 U877 ( .DIN(n1151), .Q(n1170) );
  hi1s1 U878 ( .DIN(n1133), .Q(n1171) );
  hi1s1 U879 ( .DIN(n1147), .Q(n1172) );
  hi1s1 U880 ( .DIN(n1180), .Q(n1173) );
  hi1s1 U881 ( .DIN(n1151), .Q(n1174) );
  hi1s1 U882 ( .DIN(n1180), .Q(n1175) );
  hi1s1 U883 ( .DIN(n1133), .Q(n1176) );
  hi1s1 U884 ( .DIN(n1180), .Q(n1177) );
  hi1s1 U885 ( .DIN(n1148), .Q(n1178) );
  hi1s1 U886 ( .DIN(n1133), .Q(n1179) );
  hi1s1 U887 ( .DIN(\IDinst/N40 ), .Q(n1180) );
  hi1s1 U888 ( .DIN(n1190), .Q(n1181) );
  hi1s1 U889 ( .DIN(\IDinst/N41 ), .Q(n1182) );
  hi1s1 U890 ( .DIN(\IDinst/N41 ), .Q(n1183) );
  hi1s1 U891 ( .DIN(\IDinst/N41 ), .Q(n1184) );
  hi1s1 U892 ( .DIN(\IDinst/N41 ), .Q(n1185) );
  hi1s1 U893 ( .DIN(\IDinst/N41 ), .Q(n1186) );
  hi1s1 U894 ( .DIN(\IDinst/N41 ), .Q(n1187) );
  hi1s1 U895 ( .DIN(\IDinst/N41 ), .Q(n1188) );
  hi1s1 U896 ( .DIN(\IDinst/N41 ), .Q(n1189) );
  hi1s1 U897 ( .DIN(n1182), .Q(n1190) );
  hi1s1 U898 ( .DIN(n1182), .Q(n1191) );
  hi1s1 U899 ( .DIN(n1185), .Q(n1192) );
  hi1s1 U900 ( .DIN(n1184), .Q(n1193) );
  hi1s1 U901 ( .DIN(n1187), .Q(n1194) );
  hi1s1 U902 ( .DIN(n1183), .Q(n1195) );
  hi1s1 U903 ( .DIN(n1189), .Q(n1196) );
  hi1s1 U904 ( .DIN(n1188), .Q(n1197) );
  hi1s1 U905 ( .DIN(n1295), .Q(n1198) );
  hi1s1 U906 ( .DIN(n1296), .Q(n1199) );
  hi1s1 U907 ( .DIN(n1296), .Q(n1200) );
  hi1s1 U908 ( .DIN(n1296), .Q(n1201) );
  hi1s1 U909 ( .DIN(n1296), .Q(n1202) );
  hi1s1 U910 ( .DIN(n1296), .Q(n1203) );
  hi1s1 U911 ( .DIN(n1296), .Q(n1204) );
  hi1s1 U912 ( .DIN(n1296), .Q(n1205) );
  hi1s1 U913 ( .DIN(n1296), .Q(n1206) );
  hi1s1 U914 ( .DIN(n1296), .Q(n1207) );
  hi1s1 U915 ( .DIN(n1296), .Q(n1208) );
  hi1s1 U916 ( .DIN(n1297), .Q(n1209) );
  hi1s1 U917 ( .DIN(n1297), .Q(n1210) );
  hi1s1 U918 ( .DIN(n1297), .Q(n1211) );
  hi1s1 U919 ( .DIN(n1297), .Q(n1212) );
  hi1s1 U920 ( .DIN(n1297), .Q(n1213) );
  hi1s1 U921 ( .DIN(n1297), .Q(n1214) );
  hi1s1 U922 ( .DIN(n1297), .Q(n1215) );
  hi1s1 U923 ( .DIN(n1297), .Q(n1216) );
  hi1s1 U924 ( .DIN(n1297), .Q(n1217) );
  hi1s1 U925 ( .DIN(n1297), .Q(n1218) );
  hi1s1 U926 ( .DIN(n1298), .Q(n1219) );
  hi1s1 U927 ( .DIN(n1298), .Q(n1220) );
  hi1s1 U928 ( .DIN(n1298), .Q(n1221) );
  hi1s1 U929 ( .DIN(n1298), .Q(n1222) );
  hi1s1 U930 ( .DIN(n1298), .Q(n1223) );
  hi1s1 U931 ( .DIN(n1298), .Q(n1224) );
  hi1s1 U932 ( .DIN(n1298), .Q(n1225) );
  hi1s1 U933 ( .DIN(n1298), .Q(n1226) );
  hi1s1 U934 ( .DIN(n1298), .Q(n1227) );
  hi1s1 U935 ( .DIN(n1298), .Q(n1228) );
  hi1s1 U936 ( .DIN(n1299), .Q(n1229) );
  hi1s1 U937 ( .DIN(n1299), .Q(n1230) );
  hi1s1 U938 ( .DIN(n1299), .Q(n1231) );
  hi1s1 U939 ( .DIN(n1299), .Q(n1232) );
  hi1s1 U940 ( .DIN(n1299), .Q(n1233) );
  hi1s1 U941 ( .DIN(n1299), .Q(n1234) );
  hi1s1 U942 ( .DIN(n1299), .Q(n1235) );
  hi1s1 U943 ( .DIN(n1299), .Q(n1236) );
  hi1s1 U944 ( .DIN(n1299), .Q(n1237) );
  hi1s1 U945 ( .DIN(n1300), .Q(n1238) );
  hi1s1 U946 ( .DIN(n1301), .Q(n1239) );
  hi1s1 U947 ( .DIN(n1310), .Q(n1240) );
  hi1s1 U948 ( .DIN(n1310), .Q(n1241) );
  hi1s1 U949 ( .DIN(n1310), .Q(n1242) );
  hi1s1 U950 ( .DIN(n1309), .Q(n1243) );
  hi1s1 U951 ( .DIN(n1309), .Q(n1244) );
  hi1s1 U952 ( .DIN(n1309), .Q(n1245) );
  hi1s1 U953 ( .DIN(n1308), .Q(n1246) );
  hi1s1 U954 ( .DIN(n1308), .Q(n1247) );
  hi1s1 U955 ( .DIN(n1308), .Q(n1248) );
  hi1s1 U956 ( .DIN(n1305), .Q(n1249) );
  hi1s1 U957 ( .DIN(n1302), .Q(n1250) );
  hi1s1 U958 ( .DIN(\IDinst/N44 ), .Q(n1251) );
  hi1s1 U959 ( .DIN(n1305), .Q(n1252) );
  hi1s1 U960 ( .DIN(n1306), .Q(n1253) );
  hi1s1 U961 ( .DIN(n1303), .Q(n1254) );
  hi1s1 U962 ( .DIN(n1307), .Q(n1255) );
  hi1s1 U963 ( .DIN(n1307), .Q(n1256) );
  hi1s1 U964 ( .DIN(n1307), .Q(n1257) );
  hi1s1 U965 ( .DIN(n1306), .Q(n1258) );
  hi1s1 U966 ( .DIN(n1306), .Q(n1259) );
  hi1s1 U967 ( .DIN(n1306), .Q(n1260) );
  hi1s1 U968 ( .DIN(n1305), .Q(n1261) );
  hi1s1 U969 ( .DIN(n1305), .Q(n1262) );
  hi1s1 U970 ( .DIN(n1305), .Q(n1263) );
  hi1s1 U971 ( .DIN(n1304), .Q(n1264) );
  hi1s1 U972 ( .DIN(n1304), .Q(n1265) );
  hi1s1 U973 ( .DIN(n1304), .Q(n1266) );
  hi1s1 U974 ( .DIN(n1309), .Q(n1267) );
  hi1s1 U975 ( .DIN(n1302), .Q(n1268) );
  hi1s1 U976 ( .DIN(n1310), .Q(n1269) );
  hi1s1 U977 ( .DIN(n1300), .Q(n1270) );
  hi1s1 U978 ( .DIN(\IDinst/N44 ), .Q(n1271) );
  hi1s1 U979 ( .DIN(n1310), .Q(n1272) );
  hi1s1 U980 ( .DIN(n1310), .Q(n1273) );
  hi1s1 U981 ( .DIN(n1308), .Q(n1274) );
  hi1s1 U982 ( .DIN(n1307), .Q(n1275) );
  hi1s1 U983 ( .DIN(n1309), .Q(n1276) );
  hi1s1 U984 ( .DIN(n1300), .Q(n1277) );
  hi1s1 U985 ( .DIN(n1301), .Q(n1278) );
  hi1s1 U986 ( .DIN(n1306), .Q(n1279) );
  hi1s1 U987 ( .DIN(n1303), .Q(n1280) );
  hi1s1 U988 ( .DIN(n1304), .Q(n1281) );
  hi1s1 U989 ( .DIN(\IDinst/N44 ), .Q(n1282) );
  hi1s1 U990 ( .DIN(n1304), .Q(n1283) );
  hi1s1 U991 ( .DIN(n1308), .Q(n1284) );
  hi1s1 U992 ( .DIN(n1307), .Q(n1285) );
  hi1s1 U993 ( .DIN(\IDinst/N44 ), .Q(n1286) );
  hi1s1 U994 ( .DIN(\IDinst/N44 ), .Q(n1287) );
  hi1s1 U995 ( .DIN(n1303), .Q(n1288) );
  hi1s1 U996 ( .DIN(n1303), .Q(n1289) );
  hi1s1 U997 ( .DIN(n1303), .Q(n1290) );
  hi1s1 U998 ( .DIN(n1302), .Q(n1291) );
  hi1s1 U999 ( .DIN(n1302), .Q(n1292) );
  hi1s1 U1000 ( .DIN(n1302), .Q(n1293) );
  hi1s1 U1001 ( .DIN(n1301), .Q(n1294) );
  hi1s1 U1002 ( .DIN(n1301), .Q(n1295) );
  hi1s1 U1003 ( .DIN(n1301), .Q(n1296) );
  hi1s1 U1004 ( .DIN(n1300), .Q(n1297) );
  hi1s1 U1005 ( .DIN(n1300), .Q(n1298) );
  hi1s1 U1006 ( .DIN(n1300), .Q(n1299) );
  hi1s1 U1007 ( .DIN(n1311), .Q(n1300) );
  hi1s1 U1008 ( .DIN(n1311), .Q(n1301) );
  hi1s1 U1009 ( .DIN(n1311), .Q(n1302) );
  hi1s1 U1010 ( .DIN(n1311), .Q(n1303) );
  hi1s1 U1011 ( .DIN(n1311), .Q(n1304) );
  hi1s1 U1012 ( .DIN(n1311), .Q(n1305) );
  hi1s1 U1013 ( .DIN(n1311), .Q(n1306) );
  hi1s1 U1014 ( .DIN(n1299), .Q(n1307) );
  hi1s1 U1015 ( .DIN(n1311), .Q(n1308) );
  hi1s1 U1016 ( .DIN(n1311), .Q(n1309) );
  hi1s1 U1017 ( .DIN(n1311), .Q(n1310) );
  hi1s1 U1018 ( .DIN(\IDinst/N44 ), .Q(n1311) );
  hi1s1 U1019 ( .DIN(n1360), .Q(n1312) );
  hi1s1 U1020 ( .DIN(n1360), .Q(n1313) );
  hi1s1 U1021 ( .DIN(n1360), .Q(n1314) );
  hi1s1 U1022 ( .DIN(n1360), .Q(n1315) );
  hi1s1 U1023 ( .DIN(n1360), .Q(n1316) );
  hi1s1 U1024 ( .DIN(n1361), .Q(n1317) );
  hi1s1 U1025 ( .DIN(n1361), .Q(n1318) );
  hi1s1 U1026 ( .DIN(n1361), .Q(n1319) );
  hi1s1 U1027 ( .DIN(n1361), .Q(n1320) );
  hi1s1 U1028 ( .DIN(n1361), .Q(n1321) );
  hi1s1 U1029 ( .DIN(n1361), .Q(n1322) );
  hi1s1 U1030 ( .DIN(n1361), .Q(n1323) );
  hi1s1 U1031 ( .DIN(n1361), .Q(n1324) );
  hi1s1 U1032 ( .DIN(n1361), .Q(n1325) );
  hi1s1 U1033 ( .DIN(n1361), .Q(n1326) );
  hi1s1 U1034 ( .DIN(n1347), .Q(n1327) );
  hi1s1 U1035 ( .DIN(n1349), .Q(n1328) );
  hi1s1 U1036 ( .DIN(n1340), .Q(n1329) );
  hi1s1 U1037 ( .DIN(n1344), .Q(n1330) );
  hi1s1 U1038 ( .DIN(n1361), .Q(n1331) );
  hi1s1 U1039 ( .DIN(\IDinst/N45 ), .Q(n1332) );
  hi1s1 U1040 ( .DIN(n1362), .Q(n1333) );
  hi1s1 U1041 ( .DIN(n1363), .Q(n1334) );
  hi1s1 U1042 ( .DIN(n1363), .Q(n1335) );
  hi1s1 U1043 ( .DIN(n1363), .Q(n1336) );
  hi1s1 U1044 ( .DIN(n1362), .Q(n1337) );
  hi1s1 U1045 ( .DIN(n1362), .Q(n1338) );
  hi1s1 U1046 ( .DIN(n1362), .Q(n1339) );
  hi1s1 U1047 ( .DIN(n1362), .Q(n1340) );
  hi1s1 U1048 ( .DIN(n1363), .Q(n1341) );
  hi1s1 U1049 ( .DIN(n1363), .Q(n1342) );
  hi1s1 U1050 ( .DIN(\IDinst/N45 ), .Q(n1343) );
  hi1s1 U1051 ( .DIN(\IDinst/N45 ), .Q(n1344) );
  hi1s1 U1052 ( .DIN(\IDinst/N45 ), .Q(n1345) );
  hi1s1 U1053 ( .DIN(\IDinst/N45 ), .Q(n1346) );
  hi1s1 U1054 ( .DIN(n1362), .Q(n1347) );
  hi1s1 U1055 ( .DIN(n1363), .Q(n1348) );
  hi1s1 U1056 ( .DIN(n1362), .Q(n1349) );
  hi1s1 U1057 ( .DIN(n1362), .Q(n1350) );
  hi1s1 U1058 ( .DIN(n1362), .Q(n1351) );
  hi1s1 U1059 ( .DIN(\IDinst/N45 ), .Q(n1352) );
  hi1s1 U1060 ( .DIN(n1363), .Q(n1353) );
  hi1s1 U1061 ( .DIN(\IDinst/N45 ), .Q(n1354) );
  hi1s1 U1062 ( .DIN(n1362), .Q(n1355) );
  hi1s1 U1063 ( .DIN(n1363), .Q(n1356) );
  hi1s1 U1064 ( .DIN(n1362), .Q(n1357) );
  hi1s1 U1065 ( .DIN(n1363), .Q(n1358) );
  hi1s1 U1066 ( .DIN(n1363), .Q(n1359) );
  hi1s1 U1067 ( .DIN(n1363), .Q(n1360) );
  hi1s1 U1068 ( .DIN(\IDinst/N45 ), .Q(n1361) );
  hi1s1 U1069 ( .DIN(n1352), .Q(n1362) );
  hi1s1 U1070 ( .DIN(n1332), .Q(n1363) );
  hi1s1 U1071 ( .DIN(n1372), .Q(n1364) );
  hi1s1 U1072 ( .DIN(\IDinst/N46 ), .Q(n1365) );
  hi1s1 U1073 ( .DIN(\IDinst/N46 ), .Q(n1366) );
  hi1s1 U1074 ( .DIN(\IDinst/N46 ), .Q(n1367) );
  hi1s1 U1075 ( .DIN(\IDinst/N46 ), .Q(n1368) );
  hi1s1 U1076 ( .DIN(\IDinst/N46 ), .Q(n1369) );
  hi1s1 U1077 ( .DIN(\IDinst/N46 ), .Q(n1370) );
  hi1s1 U1078 ( .DIN(\IDinst/N46 ), .Q(n1371) );
  hi1s1 U1079 ( .DIN(n1366), .Q(n1372) );
  hi1s1 U1080 ( .DIN(n1364), .Q(n1373) );
  hi1s1 U1081 ( .DIN(n1367), .Q(n1374) );
  hi1s1 U1082 ( .DIN(n1364), .Q(n1375) );
  hi1s1 U1083 ( .DIN(n1364), .Q(n1376) );
  hi1s1 U1084 ( .DIN(n1367), .Q(n1377) );
  hi1s1 U1085 ( .DIN(n1366), .Q(n1378) );
  hi1s1 U1086 ( .DIN(n1364), .Q(n1379) );
  hi1s1 U1087 ( .DIN(n1365), .Q(n1380) );
  hi1s1 U1088 ( .DIN(reset), .Q(n9588) );
  nor4s1 U1089 ( .DIN1(n1381), .DIN2(n1382), .DIN3(n47), 
        .DIN4(\IDinst/reg_dst_of_MEM[1]), .Q(PIPEEMPTY) );
  nnd3s1 U1090 ( .DIN1(FREEZE), .DIN2(n1383), .DIN3(\IDinst/n1403 ), .Q(n1382)
         );
  nnd4s1 U1091 ( .DIN1(n1384), .DIN2(n1385), .DIN3(n9419), .DIN4(n1386), 
        .Q(n1381) );
  and3s1 U1092 ( .DIN1(n9421), .DIN2(n9452), .DIN3(n9420), .Q(n1386) );
  nnd2s1 U1093 ( .DIN1(reg_dst), .DIN2(n1387), .Q(n1385) );
  nnd4s1 U1094 ( .DIN1(n9408), .DIN2(n9410), .DIN3(n1388), .DIN4(n9412), 
        .Q(n1387) );
  nor2s1 U1095 ( .DIN1(n142), .DIN2(n50), .Q(n1388) );
  nnd2s1 U1096 ( .DIN1(n1389), .DIN2(n11), .Q(n1384) );
  nnd4s1 U1097 ( .DIN1(n9407), .DIN2(n9409), .DIN3(n1390), .DIN4(n9411), 
        .Q(n1389) );
  nor2s1 U1098 ( .DIN1(n141), .DIN2(n49), .Q(n1390) );
  nnd3s1 U1099 ( .DIN1(n1391), .DIN2(n1392), .DIN3(n764), .Q(\MEMinst/N88 ) );
  nnd2s1 U1100 ( .DIN1(\DM_read_data[31] ), .DIN2(n731), .Q(n1392) );
  nnd2s1 U1101 ( .DIN1(n526), .DIN2(\DM_addr[31] ), .Q(n1391) );
  nnd3s1 U1102 ( .DIN1(n1395), .DIN2(n1396), .DIN3(n764), .Q(\MEMinst/N87 ) );
  nnd2s1 U1103 ( .DIN1(\DM_read_data[30] ), .DIN2(n731), .Q(n1396) );
  nnd2s1 U1104 ( .DIN1(n28), .DIN2(\DM_addr[30] ), .Q(n1395) );
  nnd3s1 U1105 ( .DIN1(n1397), .DIN2(n1398), .DIN3(n764), .Q(\MEMinst/N86 ) );
  nnd2s1 U1106 ( .DIN1(\DM_read_data[29] ), .DIN2(n731), .Q(n1398) );
  nnd2s1 U1107 ( .DIN1(n526), .DIN2(\DM_addr[29] ), .Q(n1397) );
  nnd3s1 U1108 ( .DIN1(n1399), .DIN2(n1400), .DIN3(n764), .Q(\MEMinst/N85 ) );
  nnd2s1 U1109 ( .DIN1(\DM_read_data[28] ), .DIN2(n731), .Q(n1400) );
  nnd2s1 U1110 ( .DIN1(n28), .DIN2(\DM_addr[28] ), .Q(n1399) );
  nnd3s1 U1111 ( .DIN1(n1401), .DIN2(n1402), .DIN3(n764), .Q(\MEMinst/N84 ) );
  nnd2s1 U1112 ( .DIN1(\DM_read_data[27] ), .DIN2(n731), .Q(n1402) );
  nnd2s1 U1113 ( .DIN1(n526), .DIN2(\DM_addr[27] ), .Q(n1401) );
  nnd3s1 U1114 ( .DIN1(n1403), .DIN2(n1404), .DIN3(n764), .Q(\MEMinst/N83 ) );
  nnd2s1 U1115 ( .DIN1(\DM_read_data[26] ), .DIN2(n731), .Q(n1404) );
  nnd2s1 U1116 ( .DIN1(n28), .DIN2(\DM_addr[26] ), .Q(n1403) );
  nnd3s1 U1117 ( .DIN1(n1405), .DIN2(n1406), .DIN3(n764), .Q(\MEMinst/N82 ) );
  nnd2s1 U1118 ( .DIN1(\DM_read_data[25] ), .DIN2(n731), .Q(n1406) );
  nnd2s1 U1119 ( .DIN1(n526), .DIN2(\DM_addr[25] ), .Q(n1405) );
  nnd3s1 U1120 ( .DIN1(n1407), .DIN2(n1408), .DIN3(n764), .Q(\MEMinst/N81 ) );
  nnd2s1 U1121 ( .DIN1(\DM_read_data[24] ), .DIN2(n731), .Q(n1408) );
  nnd2s1 U1122 ( .DIN1(n28), .DIN2(\DM_addr[24] ), .Q(n1407) );
  nnd3s1 U1123 ( .DIN1(n1409), .DIN2(n1410), .DIN3(n764), .Q(\MEMinst/N80 ) );
  nnd2s1 U1124 ( .DIN1(\DM_read_data[23] ), .DIN2(n731), .Q(n1410) );
  nnd2s1 U1125 ( .DIN1(n526), .DIN2(\DM_addr[23] ), .Q(n1409) );
  nnd3s1 U1126 ( .DIN1(n1411), .DIN2(n1412), .DIN3(n764), .Q(\MEMinst/N79 ) );
  nnd2s1 U1127 ( .DIN1(\DM_read_data[22] ), .DIN2(n731), .Q(n1412) );
  nnd2s1 U1128 ( .DIN1(n28), .DIN2(\DM_addr[22] ), .Q(n1411) );
  nnd3s1 U1129 ( .DIN1(n1413), .DIN2(n1414), .DIN3(n764), .Q(\MEMinst/N78 ) );
  nnd2s1 U1130 ( .DIN1(\DM_read_data[21] ), .DIN2(n731), .Q(n1414) );
  nnd2s1 U1131 ( .DIN1(n526), .DIN2(\DM_addr[21] ), .Q(n1413) );
  nnd3s1 U1132 ( .DIN1(n1415), .DIN2(n1416), .DIN3(n764), .Q(\MEMinst/N77 ) );
  nnd2s1 U1133 ( .DIN1(\DM_read_data[20] ), .DIN2(n731), .Q(n1416) );
  nnd2s1 U1134 ( .DIN1(n28), .DIN2(\DM_addr[20] ), .Q(n1415) );
  nnd3s1 U1135 ( .DIN1(n1417), .DIN2(n1418), .DIN3(n764), .Q(\MEMinst/N76 ) );
  nnd2s1 U1136 ( .DIN1(\DM_read_data[19] ), .DIN2(n731), .Q(n1418) );
  nnd2s1 U1137 ( .DIN1(n526), .DIN2(\DM_addr[19] ), .Q(n1417) );
  nnd3s1 U1138 ( .DIN1(n1419), .DIN2(n1420), .DIN3(n764), .Q(\MEMinst/N75 ) );
  nnd2s1 U1139 ( .DIN1(\DM_read_data[18] ), .DIN2(n731), .Q(n1420) );
  nnd2s1 U1140 ( .DIN1(n28), .DIN2(\DM_addr[18] ), .Q(n1419) );
  nnd3s1 U1141 ( .DIN1(n1421), .DIN2(n1422), .DIN3(n764), .Q(\MEMinst/N74 ) );
  nnd2s1 U1142 ( .DIN1(\DM_read_data[17] ), .DIN2(n731), .Q(n1422) );
  nnd2s1 U1143 ( .DIN1(n526), .DIN2(\DM_addr[17] ), .Q(n1421) );
  nnd3s1 U1144 ( .DIN1(n1423), .DIN2(n1424), .DIN3(n764), .Q(\MEMinst/N73 ) );
  nnd4s1 U1145 ( .DIN1(word), .DIN2(n9417), .DIN3(n1427), 
        .DIN4(\DM_read_data[15] ), .Q(n1425) );
  nor2s1 U1146 ( .DIN1(n9418), .DIN2(n526), .Q(n1427) );
  nnd2s1 U1147 ( .DIN1(\DM_read_data[16] ), .DIN2(n731), .Q(n1424) );
  nnd2s1 U1148 ( .DIN1(n380), .DIN2(n1430), .Q(n1428) );
  or2s1 U1149 ( .DIN1(byte), .DIN2(word), .Q(n1430) );
  nnd2s1 U1150 ( .DIN1(n28), .DIN2(\DM_addr[16] ), .Q(n1423) );
  nnd3s1 U1151 ( .DIN1(n1431), .DIN2(n1426), .DIN3(n1432), .Q(\MEMinst/N72 )
         );
  nnd2s1 U1152 ( .DIN1(n526), .DIN2(\DM_addr[15] ), .Q(n1432) );
  nnd2s1 U1153 ( .DIN1(n1433), .DIN2(\DM_read_data[15] ), .Q(n1431) );
  nnd3s1 U1154 ( .DIN1(n1434), .DIN2(n1426), .DIN3(n1435), .Q(\MEMinst/N71 )
         );
  nnd2s1 U1155 ( .DIN1(n28), .DIN2(\DM_addr[14] ), .Q(n1435) );
  nnd2s1 U1156 ( .DIN1(\DM_read_data[14] ), .DIN2(n1433), .Q(n1434) );
  nnd3s1 U1157 ( .DIN1(n1436), .DIN2(n1426), .DIN3(n1437), .Q(\MEMinst/N70 )
         );
  nnd2s1 U1158 ( .DIN1(n526), .DIN2(\DM_addr[13] ), .Q(n1437) );
  nnd2s1 U1159 ( .DIN1(\DM_read_data[13] ), .DIN2(n1433), .Q(n1436) );
  nnd3s1 U1160 ( .DIN1(n1438), .DIN2(n1426), .DIN3(n1439), .Q(\MEMinst/N69 )
         );
  nnd2s1 U1161 ( .DIN1(n28), .DIN2(\DM_addr[12] ), .Q(n1439) );
  nnd2s1 U1162 ( .DIN1(\DM_read_data[12] ), .DIN2(n1433), .Q(n1438) );
  nnd3s1 U1163 ( .DIN1(n1440), .DIN2(n1426), .DIN3(n1441), .Q(\MEMinst/N68 )
         );
  nnd2s1 U1164 ( .DIN1(n526), .DIN2(\DM_addr[11] ), .Q(n1441) );
  nnd2s1 U1165 ( .DIN1(\DM_read_data[11] ), .DIN2(n1433), .Q(n1440) );
  nnd3s1 U1166 ( .DIN1(n1442), .DIN2(n1426), .DIN3(n1443), .Q(\MEMinst/N67 )
         );
  nnd2s1 U1167 ( .DIN1(n28), .DIN2(\DM_addr[10] ), .Q(n1443) );
  nnd2s1 U1168 ( .DIN1(\DM_read_data[10] ), .DIN2(n1433), .Q(n1442) );
  nnd3s1 U1169 ( .DIN1(n1444), .DIN2(n1426), .DIN3(n1445), .Q(\MEMinst/N66 )
         );
  nnd2s1 U1170 ( .DIN1(n526), .DIN2(\DM_addr[9] ), .Q(n1445) );
  nnd2s1 U1171 ( .DIN1(\DM_read_data[9] ), .DIN2(n1433), .Q(n1444) );
  nnd3s1 U1172 ( .DIN1(n1446), .DIN2(n1426), .DIN3(n1447), .Q(\MEMinst/N65 )
         );
  nnd2s1 U1173 ( .DIN1(n28), .DIN2(\DM_addr[8] ), .Q(n1447) );
  nnd3s1 U1174 ( .DIN1(n1448), .DIN2(n1429), .DIN3(\DM_read_data[7] ), 
        .Q(n1426) );
  nnd2s1 U1175 ( .DIN1(\DM_read_data[8] ), .DIN2(n1433), .Q(n1446) );
  nor2s1 U1176 ( .DIN1(n1448), .DIN2(n28), .Q(n1433) );
  nor2s1 U1177 ( .DIN1(n9417), .DIN2(n9418), .Q(n1448) );
  nnd2s1 U1178 ( .DIN1(n1449), .DIN2(n1450), .Q(\MEMinst/N64 ) );
  nnd2s1 U1179 ( .DIN1(n526), .DIN2(\DM_addr[7] ), .Q(n1450) );
  nnd2s1 U1180 ( .DIN1(\DM_read_data[7] ), .DIN2(n1429), .Q(n1449) );
  nnd2s1 U1181 ( .DIN1(n1451), .DIN2(n1452), .Q(\MEMinst/N63 ) );
  nnd2s1 U1182 ( .DIN1(n28), .DIN2(\DM_addr[6] ), .Q(n1452) );
  nnd2s1 U1183 ( .DIN1(\DM_read_data[6] ), .DIN2(n1429), .Q(n1451) );
  nnd2s1 U1184 ( .DIN1(n1453), .DIN2(n1454), .Q(\MEMinst/N62 ) );
  nnd2s1 U1185 ( .DIN1(n526), .DIN2(\DM_addr[5] ), .Q(n1454) );
  nnd2s1 U1186 ( .DIN1(\DM_read_data[5] ), .DIN2(n1429), .Q(n1453) );
  nnd2s1 U1187 ( .DIN1(n1455), .DIN2(n1456), .Q(\MEMinst/N61 ) );
  nnd2s1 U1188 ( .DIN1(n28), .DIN2(\DM_addr[4] ), .Q(n1456) );
  nnd2s1 U1189 ( .DIN1(\DM_read_data[4] ), .DIN2(n1429), .Q(n1455) );
  nnd2s1 U1190 ( .DIN1(n1457), .DIN2(n1458), .Q(\MEMinst/N60 ) );
  nnd2s1 U1191 ( .DIN1(n526), .DIN2(\DM_addr[3] ), .Q(n1458) );
  nnd2s1 U1192 ( .DIN1(\DM_read_data[3] ), .DIN2(n1429), .Q(n1457) );
  nnd2s1 U1193 ( .DIN1(n1459), .DIN2(n1460), .Q(\MEMinst/N59 ) );
  nnd2s1 U1194 ( .DIN1(n28), .DIN2(\DM_addr[2] ), .Q(n1460) );
  nnd2s1 U1195 ( .DIN1(\DM_read_data[2] ), .DIN2(n1429), .Q(n1459) );
  nnd2s1 U1196 ( .DIN1(n1461), .DIN2(n1462), .Q(\MEMinst/N58 ) );
  nnd2s1 U1197 ( .DIN1(n526), .DIN2(\DM_addr[1] ), .Q(n1462) );
  nnd2s1 U1198 ( .DIN1(\DM_read_data[1] ), .DIN2(n1429), .Q(n1461) );
  nnd2s1 U1199 ( .DIN1(n1463), .DIN2(n1464), .Q(\MEMinst/N57 ) );
  nnd2s1 U1200 ( .DIN1(n28), .DIN2(\DM_addr[0] ), .Q(n1464) );
  nnd2s1 U1201 ( .DIN1(\DM_read_data[0] ), .DIN2(n1429), .Q(n1463) );
  hi1s1 U1202 ( .DIN(n526), .Q(n1429) );
  nnd2s1 U1203 ( .DIN1(n118), .DIN2(n1465), .Q(\IFinst/n848 ) );
  or2s1 U1204 ( .DIN1(n646), .DIN2(n9383), .Q(n1465) );
  nnd2s1 U1205 ( .DIN1(n1467), .DIN2(n1468), .Q(\IFinst/n847 ) );
  nnd2s1 U1206 ( .DIN1(n9523), .DIN2(n625), .Q(n1467) );
  nnd2s1 U1207 ( .DIN1(n1469), .DIN2(n1470), .Q(\IFinst/n846 ) );
  nnd2s1 U1208 ( .DIN1(n9490), .DIN2(n624), .Q(n1469) );
  nnd2s1 U1209 ( .DIN1(n1471), .DIN2(n1472), .Q(\IFinst/n845 ) );
  nnd2s1 U1210 ( .DIN1(n646), .DIN2(\NPC[2] ), .Q(n1472) );
  nnd2s1 U1211 ( .DIN1(n9492), .DIN2(n625), .Q(n1471) );
  nnd2s1 U1212 ( .DIN1(n1473), .DIN2(n1474), .Q(\IFinst/n844 ) );
  nnd2s1 U1213 ( .DIN1(n645), .DIN2(\NPC[3] ), .Q(n1474) );
  nnd2s1 U1214 ( .DIN1(n9493), .DIN2(n624), .Q(n1473) );
  nnd2s1 U1215 ( .DIN1(n1475), .DIN2(n1476), .Q(\IFinst/n843 ) );
  nnd2s1 U1216 ( .DIN1(n648), .DIN2(\NPC[4] ), .Q(n1476) );
  nnd2s1 U1217 ( .DIN1(n9494), .DIN2(n625), .Q(n1475) );
  nnd2s1 U1218 ( .DIN1(n1477), .DIN2(n1478), .Q(\IFinst/n842 ) );
  nnd2s1 U1219 ( .DIN1(n647), .DIN2(\NPC[5] ), .Q(n1478) );
  nnd2s1 U1220 ( .DIN1(n9495), .DIN2(n624), .Q(n1477) );
  nnd2s1 U1221 ( .DIN1(n1479), .DIN2(n1480), .Q(\IFinst/n841 ) );
  nnd2s1 U1222 ( .DIN1(n646), .DIN2(\NPC[6] ), .Q(n1480) );
  nnd2s1 U1223 ( .DIN1(n9496), .DIN2(n625), .Q(n1479) );
  nnd2s1 U1224 ( .DIN1(n1481), .DIN2(n1482), .Q(\IFinst/n840 ) );
  nnd2s1 U1225 ( .DIN1(n645), .DIN2(\NPC[7] ), .Q(n1482) );
  nnd2s1 U1226 ( .DIN1(n9497), .DIN2(n624), .Q(n1481) );
  nnd2s1 U1227 ( .DIN1(n1483), .DIN2(n1484), .Q(\IFinst/n839 ) );
  nnd2s1 U1228 ( .DIN1(n648), .DIN2(\NPC[8] ), .Q(n1484) );
  nnd2s1 U1229 ( .DIN1(n9498), .DIN2(n625), .Q(n1483) );
  nnd2s1 U1230 ( .DIN1(n1485), .DIN2(n1486), .Q(\IFinst/n838 ) );
  nnd2s1 U1231 ( .DIN1(n647), .DIN2(\NPC[9] ), .Q(n1486) );
  nnd2s1 U1232 ( .DIN1(n9499), .DIN2(n624), .Q(n1485) );
  nnd2s1 U1233 ( .DIN1(n1487), .DIN2(n1488), .Q(\IFinst/n837 ) );
  nnd2s1 U1234 ( .DIN1(n646), .DIN2(\NPC[10] ), .Q(n1488) );
  nnd2s1 U1235 ( .DIN1(n9500), .DIN2(n625), .Q(n1487) );
  nnd2s1 U1236 ( .DIN1(n1489), .DIN2(n1490), .Q(\IFinst/n836 ) );
  nnd2s1 U1237 ( .DIN1(n645), .DIN2(\NPC[11] ), .Q(n1490) );
  nnd2s1 U1238 ( .DIN1(n9501), .DIN2(n624), .Q(n1489) );
  nnd2s1 U1239 ( .DIN1(n1491), .DIN2(n1492), .Q(\IFinst/n835 ) );
  nnd2s1 U1240 ( .DIN1(n648), .DIN2(\NPC[12] ), .Q(n1492) );
  nnd2s1 U1241 ( .DIN1(n9502), .DIN2(n625), .Q(n1491) );
  nnd2s1 U1242 ( .DIN1(n1493), .DIN2(n1494), .Q(\IFinst/n834 ) );
  nnd2s1 U1243 ( .DIN1(n647), .DIN2(\NPC[13] ), .Q(n1494) );
  nnd2s1 U1244 ( .DIN1(n9503), .DIN2(n624), .Q(n1493) );
  nnd2s1 U1245 ( .DIN1(n1495), .DIN2(n1496), .Q(\IFinst/n833 ) );
  nnd2s1 U1246 ( .DIN1(n646), .DIN2(\NPC[14] ), .Q(n1496) );
  nnd2s1 U1247 ( .DIN1(n9504), .DIN2(n625), .Q(n1495) );
  nnd2s1 U1248 ( .DIN1(n1497), .DIN2(n1498), .Q(\IFinst/n832 ) );
  nnd2s1 U1249 ( .DIN1(n645), .DIN2(\NPC[15] ), .Q(n1498) );
  nnd2s1 U1250 ( .DIN1(n9505), .DIN2(n624), .Q(n1497) );
  nnd2s1 U1251 ( .DIN1(n1499), .DIN2(n1500), .Q(\IFinst/n831 ) );
  nnd2s1 U1252 ( .DIN1(n648), .DIN2(\NPC[16] ), .Q(n1500) );
  nnd2s1 U1253 ( .DIN1(n9506), .DIN2(n625), .Q(n1499) );
  nnd2s1 U1254 ( .DIN1(n1501), .DIN2(n1502), .Q(\IFinst/n830 ) );
  nnd2s1 U1255 ( .DIN1(n647), .DIN2(\NPC[17] ), .Q(n1502) );
  nnd2s1 U1256 ( .DIN1(n9507), .DIN2(n624), .Q(n1501) );
  nnd2s1 U1257 ( .DIN1(n1503), .DIN2(n1504), .Q(\IFinst/n829 ) );
  nnd2s1 U1258 ( .DIN1(n646), .DIN2(\NPC[18] ), .Q(n1504) );
  nnd2s1 U1259 ( .DIN1(n9508), .DIN2(n625), .Q(n1503) );
  nnd2s1 U1260 ( .DIN1(n1505), .DIN2(n1506), .Q(\IFinst/n828 ) );
  nnd2s1 U1261 ( .DIN1(n645), .DIN2(\NPC[19] ), .Q(n1506) );
  nnd2s1 U1262 ( .DIN1(n9509), .DIN2(n624), .Q(n1505) );
  nnd2s1 U1263 ( .DIN1(n1507), .DIN2(n1508), .Q(\IFinst/n827 ) );
  nnd2s1 U1264 ( .DIN1(n648), .DIN2(\NPC[20] ), .Q(n1508) );
  nnd2s1 U1265 ( .DIN1(n9510), .DIN2(n625), .Q(n1507) );
  nnd2s1 U1266 ( .DIN1(n1509), .DIN2(n1510), .Q(\IFinst/n826 ) );
  nnd2s1 U1267 ( .DIN1(n647), .DIN2(\NPC[21] ), .Q(n1510) );
  nnd2s1 U1268 ( .DIN1(n9511), .DIN2(n624), .Q(n1509) );
  nnd2s1 U1269 ( .DIN1(n1511), .DIN2(n1512), .Q(\IFinst/n825 ) );
  nnd2s1 U1270 ( .DIN1(n646), .DIN2(\NPC[22] ), .Q(n1512) );
  nnd2s1 U1271 ( .DIN1(n9512), .DIN2(n625), .Q(n1511) );
  nnd2s1 U1272 ( .DIN1(n1513), .DIN2(n1514), .Q(\IFinst/n824 ) );
  nnd2s1 U1273 ( .DIN1(n645), .DIN2(\NPC[23] ), .Q(n1514) );
  nnd2s1 U1274 ( .DIN1(n9513), .DIN2(n624), .Q(n1513) );
  nnd2s1 U1275 ( .DIN1(n1515), .DIN2(n1516), .Q(\IFinst/n823 ) );
  nnd2s1 U1276 ( .DIN1(n648), .DIN2(\NPC[24] ), .Q(n1516) );
  nnd2s1 U1277 ( .DIN1(n9514), .DIN2(n625), .Q(n1515) );
  nnd2s1 U1278 ( .DIN1(n1517), .DIN2(n1518), .Q(\IFinst/n822 ) );
  nnd2s1 U1279 ( .DIN1(n647), .DIN2(\NPC[25] ), .Q(n1518) );
  nnd2s1 U1280 ( .DIN1(n9515), .DIN2(n624), .Q(n1517) );
  nnd2s1 U1281 ( .DIN1(n1519), .DIN2(n1520), .Q(\IFinst/n821 ) );
  nnd2s1 U1282 ( .DIN1(n646), .DIN2(\NPC[26] ), .Q(n1520) );
  nnd2s1 U1283 ( .DIN1(n9516), .DIN2(n625), .Q(n1519) );
  nnd2s1 U1284 ( .DIN1(n1521), .DIN2(n1522), .Q(\IFinst/n820 ) );
  nnd2s1 U1285 ( .DIN1(n645), .DIN2(\NPC[27] ), .Q(n1522) );
  nnd2s1 U1286 ( .DIN1(n9517), .DIN2(n624), .Q(n1521) );
  nnd2s1 U1287 ( .DIN1(n1523), .DIN2(n1524), .Q(\IFinst/n819 ) );
  nnd2s1 U1288 ( .DIN1(n648), .DIN2(\NPC[28] ), .Q(n1524) );
  nnd2s1 U1289 ( .DIN1(n9518), .DIN2(n625), .Q(n1523) );
  nnd2s1 U1290 ( .DIN1(n1525), .DIN2(n1526), .Q(\IFinst/n818 ) );
  nnd2s1 U1291 ( .DIN1(n647), .DIN2(\NPC[29] ), .Q(n1526) );
  nnd2s1 U1292 ( .DIN1(n9519), .DIN2(n624), .Q(n1525) );
  nnd2s1 U1293 ( .DIN1(n1527), .DIN2(n1528), .Q(\IFinst/n817 ) );
  nnd2s1 U1294 ( .DIN1(n646), .DIN2(\NPC[30] ), .Q(n1528) );
  nnd2s1 U1295 ( .DIN1(n9521), .DIN2(n625), .Q(n1527) );
  nnd2s1 U1296 ( .DIN1(n1529), .DIN2(n1530), .Q(\IFinst/n816 ) );
  nnd2s1 U1297 ( .DIN1(n645), .DIN2(\NPC[31] ), .Q(n1530) );
  nnd2s1 U1298 ( .DIN1(n9522), .DIN2(n624), .Q(n1529) );
  nnd2s1 U1299 ( .DIN1(n1531), .DIN2(n1532), .Q(\IFinst/n749 ) );
  nnd2s1 U1300 ( .DIN1(n9524), .DIN2(n684), .Q(n1532) );
  nnd2s1 U1301 ( .DIN1(\IR[31] ), .DIN2(n664), .Q(n1531) );
  nnd2s1 U1302 ( .DIN1(n1533), .DIN2(n1534), .Q(\IFinst/n746 ) );
  nnd2s1 U1303 ( .DIN1(n663), .DIN2(n322), .Q(n1534) );
  nnd2s1 U1304 ( .DIN1(n9525), .DIN2(n685), .Q(n1533) );
  nnd2s1 U1305 ( .DIN1(n1535), .DIN2(n1536), .Q(\IFinst/n744 ) );
  nnd2s1 U1306 ( .DIN1(n9526), .DIN2(n687), .Q(n1536) );
  nnd2s1 U1307 ( .DIN1(\IR[30] ), .DIN2(n662), .Q(n1535) );
  nnd2s1 U1308 ( .DIN1(n1537), .DIN2(n1538), .Q(\IFinst/n741 ) );
  nnd2s1 U1309 ( .DIN1(n662), .DIN2(n316), .Q(n1538) );
  nnd2s1 U1310 ( .DIN1(n9527), .DIN2(n686), .Q(n1537) );
  nnd2s1 U1311 ( .DIN1(n1539), .DIN2(n1540), .Q(\IFinst/n739 ) );
  nnd2s1 U1312 ( .DIN1(n9528), .DIN2(n684), .Q(n1540) );
  nnd2s1 U1313 ( .DIN1(\IR[29] ), .DIN2(n663), .Q(n1539) );
  nnd2s1 U1314 ( .DIN1(n1541), .DIN2(n1542), .Q(\IFinst/n736 ) );
  nnd2s1 U1315 ( .DIN1(n661), .DIN2(n326), .Q(n1542) );
  nnd2s1 U1316 ( .DIN1(n9529), .DIN2(n685), .Q(n1541) );
  nnd2s1 U1317 ( .DIN1(n1543), .DIN2(n1544), .Q(\IFinst/n734 ) );
  nnd2s1 U1318 ( .DIN1(n9530), .DIN2(n687), .Q(n1544) );
  nnd2s1 U1319 ( .DIN1(\IR[28] ), .DIN2(n661), .Q(n1543) );
  nnd2s1 U1320 ( .DIN1(n1545), .DIN2(n1546), .Q(\IFinst/n731 ) );
  nnd2s1 U1321 ( .DIN1(n664), .DIN2(n324), .Q(n1546) );
  nnd2s1 U1322 ( .DIN1(n9531), .DIN2(n686), .Q(n1545) );
  nnd2s1 U1323 ( .DIN1(n1547), .DIN2(n1548), .Q(\IFinst/n729 ) );
  nnd2s1 U1324 ( .DIN1(n9532), .DIN2(n684), .Q(n1548) );
  nnd2s1 U1325 ( .DIN1(\IR[27] ), .DIN2(n664), .Q(n1547) );
  nnd2s1 U1326 ( .DIN1(n1549), .DIN2(n1550), .Q(\IFinst/n726 ) );
  nnd2s1 U1327 ( .DIN1(n663), .DIN2(n320), .Q(n1550) );
  nnd2s1 U1328 ( .DIN1(n9533), .DIN2(n685), .Q(n1549) );
  nnd2s1 U1329 ( .DIN1(n1551), .DIN2(n1552), .Q(\IFinst/n724 ) );
  nnd2s1 U1330 ( .DIN1(n9534), .DIN2(n687), .Q(n1552) );
  nnd2s1 U1331 ( .DIN1(\IR[26] ), .DIN2(n662), .Q(n1551) );
  nnd2s1 U1332 ( .DIN1(n1553), .DIN2(n1554), .Q(\IFinst/n721 ) );
  nnd2s1 U1333 ( .DIN1(n662), .DIN2(n318), .Q(n1554) );
  nnd2s1 U1334 ( .DIN1(n9535), .DIN2(n686), .Q(n1553) );
  nnd2s1 U1335 ( .DIN1(n1555), .DIN2(n1556), .Q(\IFinst/n719 ) );
  nnd2s1 U1336 ( .DIN1(n9536), .DIN2(n684), .Q(n1556) );
  nnd2s1 U1337 ( .DIN1(\IR[25] ), .DIN2(n663), .Q(n1555) );
  nnd2s1 U1338 ( .DIN1(n1557), .DIN2(n1558), .Q(\IFinst/n716 ) );
  nnd2s1 U1339 ( .DIN1(n661), .DIN2(n310), .Q(n1558) );
  nnd2s1 U1340 ( .DIN1(n9537), .DIN2(n685), .Q(n1557) );
  nnd2s1 U1341 ( .DIN1(n1559), .DIN2(n1560), .Q(\IFinst/n714 ) );
  nnd2s1 U1342 ( .DIN1(n9538), .DIN2(n687), .Q(n1560) );
  nnd2s1 U1343 ( .DIN1(\IR[24] ), .DIN2(n661), .Q(n1559) );
  nnd2s1 U1344 ( .DIN1(n1561), .DIN2(n1562), .Q(\IFinst/n711 ) );
  nnd2s1 U1345 ( .DIN1(n664), .DIN2(n314), .Q(n1562) );
  nnd2s1 U1346 ( .DIN1(n9539), .DIN2(n686), .Q(n1561) );
  nnd2s1 U1347 ( .DIN1(n1563), .DIN2(n1564), .Q(\IFinst/n709 ) );
  nnd2s1 U1348 ( .DIN1(n9540), .DIN2(n684), .Q(n1564) );
  nnd2s1 U1349 ( .DIN1(\IR[23] ), .DIN2(n664), .Q(n1563) );
  nnd2s1 U1350 ( .DIN1(n1565), .DIN2(n1566), .Q(\IFinst/n706 ) );
  nnd2s1 U1351 ( .DIN1(n663), .DIN2(n312), .Q(n1566) );
  nnd2s1 U1352 ( .DIN1(n9541), .DIN2(n685), .Q(n1565) );
  nnd2s1 U1353 ( .DIN1(n1567), .DIN2(n1568), .Q(\IFinst/n704 ) );
  nnd2s1 U1354 ( .DIN1(n9542), .DIN2(n687), .Q(n1568) );
  nnd2s1 U1355 ( .DIN1(\IR[22] ), .DIN2(n662), .Q(n1567) );
  nnd2s1 U1356 ( .DIN1(n1569), .DIN2(n1570), .Q(\IFinst/n701 ) );
  nnd2s1 U1357 ( .DIN1(n662), .DIN2(n306), .Q(n1570) );
  nnd2s1 U1358 ( .DIN1(n9543), .DIN2(n686), .Q(n1569) );
  nnd2s1 U1359 ( .DIN1(n1571), .DIN2(n1572), .Q(\IFinst/n699 ) );
  nnd2s1 U1360 ( .DIN1(n9544), .DIN2(n684), .Q(n1572) );
  nnd2s1 U1361 ( .DIN1(\IR[21] ), .DIN2(n663), .Q(n1571) );
  nnd2s1 U1362 ( .DIN1(n1573), .DIN2(n1574), .Q(\IFinst/n696 ) );
  nnd2s1 U1363 ( .DIN1(n661), .DIN2(n308), .Q(n1574) );
  nnd2s1 U1364 ( .DIN1(n9545), .DIN2(n685), .Q(n1573) );
  nnd2s1 U1365 ( .DIN1(n1575), .DIN2(n1576), .Q(\IFinst/n694 ) );
  nnd2s1 U1366 ( .DIN1(n9546), .DIN2(n687), .Q(n1576) );
  nnd2s1 U1367 ( .DIN1(\IR[20] ), .DIN2(n661), .Q(n1575) );
  nnd2s1 U1368 ( .DIN1(n1577), .DIN2(n1578), .Q(\IFinst/n691 ) );
  nnd2s1 U1369 ( .DIN1(n664), .DIN2(n276), .Q(n1578) );
  nnd2s1 U1370 ( .DIN1(n9547), .DIN2(n686), .Q(n1577) );
  nnd2s1 U1371 ( .DIN1(n1579), .DIN2(n1580), .Q(\IFinst/n689 ) );
  nnd2s1 U1372 ( .DIN1(n9548), .DIN2(n684), .Q(n1580) );
  nnd2s1 U1373 ( .DIN1(\IR[19] ), .DIN2(n664), .Q(n1579) );
  nnd2s1 U1374 ( .DIN1(n1581), .DIN2(n1582), .Q(\IFinst/n686 ) );
  nnd2s1 U1375 ( .DIN1(n663), .DIN2(n280), .Q(n1582) );
  nnd2s1 U1376 ( .DIN1(n9549), .DIN2(n685), .Q(n1581) );
  nnd2s1 U1377 ( .DIN1(n1583), .DIN2(n1584), .Q(\IFinst/n684 ) );
  nnd2s1 U1378 ( .DIN1(n9550), .DIN2(n687), .Q(n1584) );
  nnd2s1 U1379 ( .DIN1(\IR[18] ), .DIN2(n662), .Q(n1583) );
  nnd2s1 U1380 ( .DIN1(n1585), .DIN2(n1586), .Q(\IFinst/n681 ) );
  nnd2s1 U1381 ( .DIN1(n662), .DIN2(n278), .Q(n1586) );
  nnd2s1 U1382 ( .DIN1(n9551), .DIN2(n686), .Q(n1585) );
  nnd2s1 U1383 ( .DIN1(n1587), .DIN2(n1588), .Q(\IFinst/n679 ) );
  nnd2s1 U1384 ( .DIN1(n9552), .DIN2(n684), .Q(n1588) );
  nnd2s1 U1385 ( .DIN1(\IR[17] ), .DIN2(n663), .Q(n1587) );
  nnd2s1 U1386 ( .DIN1(n1589), .DIN2(n1590), .Q(\IFinst/n676 ) );
  nnd2s1 U1387 ( .DIN1(n661), .DIN2(n274), .Q(n1590) );
  nnd2s1 U1388 ( .DIN1(n9553), .DIN2(n685), .Q(n1589) );
  nnd2s1 U1389 ( .DIN1(n1591), .DIN2(n1592), .Q(\IFinst/n674 ) );
  nnd2s1 U1390 ( .DIN1(n9554), .DIN2(n684), .Q(n1592) );
  nnd2s1 U1391 ( .DIN1(\IR[16] ), .DIN2(n661), .Q(n1591) );
  nnd2s1 U1392 ( .DIN1(n1593), .DIN2(n1594), .Q(\IFinst/n671 ) );
  nnd2s1 U1393 ( .DIN1(n664), .DIN2(n272), .Q(n1594) );
  nnd2s1 U1394 ( .DIN1(n9555), .DIN2(n687), .Q(n1593) );
  nnd2s1 U1395 ( .DIN1(n1595), .DIN2(n1596), .Q(\IFinst/n669 ) );
  nnd2s1 U1396 ( .DIN1(n9556), .DIN2(n686), .Q(n1596) );
  nnd2s1 U1397 ( .DIN1(\IR[15] ), .DIN2(n664), .Q(n1595) );
  nnd2s1 U1398 ( .DIN1(n1597), .DIN2(n1598), .Q(\IFinst/n666 ) );
  nnd2s1 U1399 ( .DIN1(n663), .DIN2(n92), .Q(n1598) );
  nnd2s1 U1400 ( .DIN1(n9557), .DIN2(n685), .Q(n1597) );
  nnd2s1 U1401 ( .DIN1(n1599), .DIN2(n1600), .Q(\IFinst/n664 ) );
  nnd2s1 U1402 ( .DIN1(n9558), .DIN2(n684), .Q(n1600) );
  nnd2s1 U1403 ( .DIN1(\IR[14] ), .DIN2(n662), .Q(n1599) );
  nnd2s1 U1404 ( .DIN1(n1601), .DIN2(n1602), .Q(\IFinst/n661 ) );
  nnd2s1 U1405 ( .DIN1(n662), .DIN2(n97), .Q(n1602) );
  nnd2s1 U1406 ( .DIN1(n9559), .DIN2(n687), .Q(n1601) );
  nnd2s1 U1407 ( .DIN1(n1603), .DIN2(n1604), .Q(\IFinst/n659 ) );
  nnd2s1 U1408 ( .DIN1(n9560), .DIN2(n686), .Q(n1604) );
  nnd2s1 U1409 ( .DIN1(\IR[13] ), .DIN2(n663), .Q(n1603) );
  nnd2s1 U1410 ( .DIN1(n1605), .DIN2(n1606), .Q(\IFinst/n656 ) );
  nnd2s1 U1411 ( .DIN1(n661), .DIN2(n113), .Q(n1606) );
  nnd2s1 U1412 ( .DIN1(n9561), .DIN2(n685), .Q(n1605) );
  nnd2s1 U1413 ( .DIN1(n1607), .DIN2(n1608), .Q(\IFinst/n654 ) );
  nnd2s1 U1414 ( .DIN1(n9562), .DIN2(n684), .Q(n1608) );
  nnd2s1 U1415 ( .DIN1(\IR[12] ), .DIN2(n661), .Q(n1607) );
  nnd2s1 U1416 ( .DIN1(n1609), .DIN2(n1610), .Q(\IFinst/n651 ) );
  nnd2s1 U1417 ( .DIN1(n664), .DIN2(n98), .Q(n1610) );
  nnd2s1 U1418 ( .DIN1(n9563), .DIN2(n687), .Q(n1609) );
  nnd2s1 U1419 ( .DIN1(n1611), .DIN2(n1612), .Q(\IFinst/n649 ) );
  nnd2s1 U1420 ( .DIN1(n9564), .DIN2(n686), .Q(n1612) );
  nnd2s1 U1421 ( .DIN1(\IR[11] ), .DIN2(n664), .Q(n1611) );
  nnd2s1 U1422 ( .DIN1(n1613), .DIN2(n1614), .Q(\IFinst/n646 ) );
  nnd2s1 U1423 ( .DIN1(n663), .DIN2(n114), .Q(n1614) );
  nnd2s1 U1424 ( .DIN1(n9565), .DIN2(n685), .Q(n1613) );
  nnd2s1 U1425 ( .DIN1(n1615), .DIN2(n1616), .Q(\IFinst/n644 ) );
  nnd2s1 U1426 ( .DIN1(n9566), .DIN2(n684), .Q(n1616) );
  nnd2s1 U1427 ( .DIN1(\IR[10] ), .DIN2(n662), .Q(n1615) );
  nnd2s1 U1428 ( .DIN1(n1617), .DIN2(n1618), .Q(\IFinst/n641 ) );
  nnd2s1 U1429 ( .DIN1(n662), .DIN2(n110), .Q(n1618) );
  nnd2s1 U1430 ( .DIN1(n9567), .DIN2(n687), .Q(n1617) );
  nnd2s1 U1431 ( .DIN1(n1619), .DIN2(n1620), .Q(\IFinst/n639 ) );
  nnd2s1 U1432 ( .DIN1(n9568), .DIN2(n686), .Q(n1620) );
  nnd2s1 U1433 ( .DIN1(\IR[9] ), .DIN2(n663), .Q(n1619) );
  nnd2s1 U1434 ( .DIN1(n1621), .DIN2(n1622), .Q(\IFinst/n636 ) );
  nnd2s1 U1435 ( .DIN1(n661), .DIN2(n125), .Q(n1622) );
  nnd2s1 U1436 ( .DIN1(n9569), .DIN2(n685), .Q(n1621) );
  nnd2s1 U1437 ( .DIN1(n1623), .DIN2(n1624), .Q(\IFinst/n634 ) );
  nnd2s1 U1438 ( .DIN1(n9570), .DIN2(n684), .Q(n1624) );
  nnd2s1 U1439 ( .DIN1(\IR[8] ), .DIN2(n661), .Q(n1623) );
  nnd2s1 U1440 ( .DIN1(n1625), .DIN2(n1626), .Q(\IFinst/n631 ) );
  nnd2s1 U1441 ( .DIN1(n664), .DIN2(n111), .Q(n1626) );
  nnd2s1 U1442 ( .DIN1(n9571), .DIN2(n687), .Q(n1625) );
  nnd2s1 U1443 ( .DIN1(n1627), .DIN2(n1628), .Q(\IFinst/n629 ) );
  nnd2s1 U1444 ( .DIN1(n9572), .DIN2(n686), .Q(n1628) );
  nnd2s1 U1445 ( .DIN1(\IR[7] ), .DIN2(n664), .Q(n1627) );
  nnd2s1 U1446 ( .DIN1(n1629), .DIN2(n1630), .Q(\IFinst/n626 ) );
  nnd2s1 U1447 ( .DIN1(n663), .DIN2(n126), .Q(n1630) );
  nnd2s1 U1448 ( .DIN1(n9573), .DIN2(n685), .Q(n1629) );
  nnd2s1 U1449 ( .DIN1(n1631), .DIN2(n1632), .Q(\IFinst/n624 ) );
  nnd2s1 U1450 ( .DIN1(n9574), .DIN2(n684), .Q(n1632) );
  nnd2s1 U1451 ( .DIN1(\IR[6] ), .DIN2(n662), .Q(n1631) );
  nnd2s1 U1452 ( .DIN1(n1633), .DIN2(n1634), .Q(\IFinst/n621 ) );
  nnd2s1 U1453 ( .DIN1(n662), .DIN2(n112), .Q(n1634) );
  nnd2s1 U1454 ( .DIN1(n9575), .DIN2(n687), .Q(n1633) );
  nnd2s1 U1455 ( .DIN1(n1635), .DIN2(n1636), .Q(\IFinst/n619 ) );
  nnd2s1 U1456 ( .DIN1(n9576), .DIN2(n686), .Q(n1636) );
  nnd2s1 U1457 ( .DIN1(\IR[5] ), .DIN2(n663), .Q(n1635) );
  nnd2s1 U1458 ( .DIN1(n1637), .DIN2(n1638), .Q(\IFinst/n616 ) );
  nnd2s1 U1459 ( .DIN1(n661), .DIN2(n115), .Q(n1638) );
  nnd2s1 U1460 ( .DIN1(n9577), .DIN2(n685), .Q(n1637) );
  nnd2s1 U1461 ( .DIN1(n1639), .DIN2(n1640), .Q(\IFinst/n614 ) );
  nnd2s1 U1462 ( .DIN1(n9578), .DIN2(n684), .Q(n1640) );
  nnd2s1 U1463 ( .DIN1(\IR[4] ), .DIN2(n661), .Q(n1639) );
  nnd2s1 U1464 ( .DIN1(n1641), .DIN2(n1642), .Q(\IFinst/n611 ) );
  nnd2s1 U1465 ( .DIN1(n664), .DIN2(n99), .Q(n1642) );
  nnd2s1 U1466 ( .DIN1(n9579), .DIN2(n687), .Q(n1641) );
  nnd2s1 U1467 ( .DIN1(n1643), .DIN2(n1644), .Q(\IFinst/n609 ) );
  nnd2s1 U1468 ( .DIN1(n9580), .DIN2(n686), .Q(n1644) );
  nnd2s1 U1469 ( .DIN1(\IR[3] ), .DIN2(n664), .Q(n1643) );
  nnd2s1 U1470 ( .DIN1(n1645), .DIN2(n1646), .Q(\IFinst/n606 ) );
  nnd2s1 U1471 ( .DIN1(n663), .DIN2(n116), .Q(n1646) );
  nnd2s1 U1472 ( .DIN1(n9581), .DIN2(n685), .Q(n1645) );
  nnd2s1 U1473 ( .DIN1(n1647), .DIN2(n1648), .Q(\IFinst/n604 ) );
  nnd2s1 U1474 ( .DIN1(n9582), .DIN2(n684), .Q(n1648) );
  nnd2s1 U1475 ( .DIN1(\IR[2] ), .DIN2(n662), .Q(n1647) );
  nnd2s1 U1476 ( .DIN1(n1649), .DIN2(n1650), .Q(\IFinst/n601 ) );
  nnd2s1 U1477 ( .DIN1(n661), .DIN2(n100), .Q(n1650) );
  nnd2s1 U1478 ( .DIN1(n9583), .DIN2(n687), .Q(n1649) );
  nnd2s1 U1479 ( .DIN1(n1651), .DIN2(n1652), .Q(\IFinst/n599 ) );
  nnd2s1 U1480 ( .DIN1(n9584), .DIN2(n686), .Q(n1652) );
  nnd2s1 U1481 ( .DIN1(\IR[1] ), .DIN2(n661), .Q(n1651) );
  nnd2s1 U1482 ( .DIN1(n1653), .DIN2(n1654), .Q(\IFinst/n596 ) );
  nnd2s1 U1483 ( .DIN1(n664), .DIN2(n42), .Q(n1654) );
  nnd2s1 U1484 ( .DIN1(n9585), .DIN2(n684), .Q(n1653) );
  nnd2s1 U1485 ( .DIN1(n1655), .DIN2(n1656), .Q(\IFinst/n594 ) );
  nnd2s1 U1486 ( .DIN1(n9586), .DIN2(n687), .Q(n1656) );
  nnd2s1 U1487 ( .DIN1(\IR[0] ), .DIN2(n664), .Q(n1655) );
  nnd2s1 U1488 ( .DIN1(n1657), .DIN2(n1658), .Q(\IFinst/n591 ) );
  nnd2s1 U1489 ( .DIN1(n663), .DIN2(n41), .Q(n1658) );
  nnd2s1 U1490 ( .DIN1(n9587), .DIN2(n686), .Q(n1657) );
  nnd3s1 U1491 ( .DIN1(n1659), .DIN2(n1660), .DIN3(n1661), .Q(\IFinst/N99 ) );
  nnd2s1 U1492 ( .DIN1(n804), .DIN2(n260), .Q(n1661) );
  nnd2s1 U1493 ( .DIN1(n1663), .DIN2(n645), .Q(n1660) );
  xnr2s1 U1494 ( .DIN1(n1664), .DIN2(\NPC[27] ), .Q(n1663) );
  nnd2s1 U1495 ( .DIN1(n657), .DIN2(n9517), .Q(n1659) );
  nnd3s1 U1496 ( .DIN1(n1665), .DIN2(n1666), .DIN3(n1667), .Q(\IFinst/N98 ) );
  nnd2s1 U1497 ( .DIN1(n804), .DIN2(n259), .Q(n1667) );
  nnd2s1 U1498 ( .DIN1(n1668), .DIN2(n648), .Q(n1666) );
  xnr2s1 U1499 ( .DIN1(n9428), .DIN2(n1669), .Q(n1668) );
  nnd2s1 U1500 ( .DIN1(n660), .DIN2(n9516), .Q(n1665) );
  nnd3s1 U1501 ( .DIN1(n1670), .DIN2(n1671), .DIN3(n1672), .Q(\IFinst/N97 ) );
  nnd2s1 U1502 ( .DIN1(n804), .DIN2(n258), .Q(n1672) );
  nnd2s1 U1503 ( .DIN1(n1673), .DIN2(n647), .Q(n1671) );
  xnr2s1 U1504 ( .DIN1(n1674), .DIN2(\NPC[25] ), .Q(n1673) );
  nnd2s1 U1505 ( .DIN1(n659), .DIN2(n9515), .Q(n1670) );
  nnd3s1 U1506 ( .DIN1(n1675), .DIN2(n1676), .DIN3(n1677), .Q(\IFinst/N96 ) );
  nnd2s1 U1507 ( .DIN1(n804), .DIN2(n257), .Q(n1677) );
  nnd2s1 U1508 ( .DIN1(n1678), .DIN2(n646), .Q(n1676) );
  xnr2s1 U1509 ( .DIN1(n9430), .DIN2(n1679), .Q(n1678) );
  nnd2s1 U1510 ( .DIN1(n658), .DIN2(n9514), .Q(n1675) );
  nnd3s1 U1511 ( .DIN1(n1680), .DIN2(n1681), .DIN3(n1682), .Q(\IFinst/N95 ) );
  nnd2s1 U1512 ( .DIN1(n804), .DIN2(n256), .Q(n1682) );
  nnd2s1 U1513 ( .DIN1(n1683), .DIN2(n645), .Q(n1681) );
  xnr2s1 U1514 ( .DIN1(n1684), .DIN2(\NPC[23] ), .Q(n1683) );
  nnd2s1 U1515 ( .DIN1(n657), .DIN2(n9513), .Q(n1680) );
  nnd3s1 U1516 ( .DIN1(n1685), .DIN2(n1686), .DIN3(n1687), .Q(\IFinst/N94 ) );
  nnd2s1 U1517 ( .DIN1(n804), .DIN2(n255), .Q(n1687) );
  nnd2s1 U1518 ( .DIN1(n1688), .DIN2(n648), .Q(n1686) );
  xnr2s1 U1519 ( .DIN1(n9432), .DIN2(n1689), .Q(n1688) );
  nnd2s1 U1520 ( .DIN1(n660), .DIN2(n9512), .Q(n1685) );
  nnd3s1 U1521 ( .DIN1(n1690), .DIN2(n1691), .DIN3(n1692), .Q(\IFinst/N93 ) );
  nnd2s1 U1522 ( .DIN1(n804), .DIN2(n254), .Q(n1692) );
  nnd2s1 U1523 ( .DIN1(n1693), .DIN2(n647), .Q(n1691) );
  xnr2s1 U1524 ( .DIN1(n1694), .DIN2(\NPC[21] ), .Q(n1693) );
  nnd2s1 U1525 ( .DIN1(n659), .DIN2(n9511), .Q(n1690) );
  nnd3s1 U1526 ( .DIN1(n1695), .DIN2(n1696), .DIN3(n1697), .Q(\IFinst/N92 ) );
  nnd2s1 U1527 ( .DIN1(n804), .DIN2(n253), .Q(n1697) );
  nnd2s1 U1528 ( .DIN1(n1698), .DIN2(n646), .Q(n1696) );
  xnr2s1 U1529 ( .DIN1(n9434), .DIN2(n1699), .Q(n1698) );
  nnd2s1 U1530 ( .DIN1(n658), .DIN2(n9510), .Q(n1695) );
  nnd3s1 U1531 ( .DIN1(n1700), .DIN2(n1701), .DIN3(n1702), .Q(\IFinst/N91 ) );
  nnd2s1 U1532 ( .DIN1(n804), .DIN2(n252), .Q(n1702) );
  nnd2s1 U1533 ( .DIN1(n1703), .DIN2(n645), .Q(n1701) );
  xnr2s1 U1534 ( .DIN1(n1704), .DIN2(\NPC[19] ), .Q(n1703) );
  nnd2s1 U1535 ( .DIN1(n657), .DIN2(n9509), .Q(n1700) );
  nnd3s1 U1536 ( .DIN1(n1705), .DIN2(n1706), .DIN3(n1707), .Q(\IFinst/N90 ) );
  nnd2s1 U1537 ( .DIN1(n804), .DIN2(n251), .Q(n1707) );
  nnd2s1 U1538 ( .DIN1(n1708), .DIN2(n648), .Q(n1706) );
  xnr2s1 U1539 ( .DIN1(n9436), .DIN2(n1709), .Q(n1708) );
  nnd2s1 U1540 ( .DIN1(n660), .DIN2(n9508), .Q(n1705) );
  nnd3s1 U1541 ( .DIN1(n1710), .DIN2(n1711), .DIN3(n1712), .Q(\IFinst/N89 ) );
  nnd2s1 U1542 ( .DIN1(n804), .DIN2(n250), .Q(n1712) );
  nnd2s1 U1543 ( .DIN1(n1713), .DIN2(n647), .Q(n1711) );
  xnr2s1 U1544 ( .DIN1(n1714), .DIN2(\NPC[17] ), .Q(n1713) );
  nnd2s1 U1545 ( .DIN1(n659), .DIN2(n9507), .Q(n1710) );
  nnd3s1 U1546 ( .DIN1(n1715), .DIN2(n1716), .DIN3(n1717), .Q(\IFinst/N88 ) );
  nnd2s1 U1547 ( .DIN1(n804), .DIN2(n249), .Q(n1717) );
  nnd2s1 U1548 ( .DIN1(n1718), .DIN2(n646), .Q(n1716) );
  xnr2s1 U1549 ( .DIN1(n9438), .DIN2(n1719), .Q(n1718) );
  nnd2s1 U1550 ( .DIN1(n658), .DIN2(n9506), .Q(n1715) );
  nnd3s1 U1551 ( .DIN1(n1720), .DIN2(n1721), .DIN3(n1722), .Q(\IFinst/N87 ) );
  nnd2s1 U1552 ( .DIN1(n804), .DIN2(n248), .Q(n1722) );
  nnd2s1 U1553 ( .DIN1(n1723), .DIN2(n645), .Q(n1721) );
  xnr2s1 U1554 ( .DIN1(n1724), .DIN2(\NPC[15] ), .Q(n1723) );
  nnd2s1 U1555 ( .DIN1(n657), .DIN2(n9505), .Q(n1720) );
  nnd3s1 U1556 ( .DIN1(n1725), .DIN2(n1726), .DIN3(n1727), .Q(\IFinst/N86 ) );
  nnd2s1 U1557 ( .DIN1(n804), .DIN2(n247), .Q(n1727) );
  nnd2s1 U1558 ( .DIN1(n1728), .DIN2(n648), .Q(n1726) );
  xnr2s1 U1559 ( .DIN1(n9440), .DIN2(n1729), .Q(n1728) );
  nnd2s1 U1560 ( .DIN1(n660), .DIN2(n9504), .Q(n1725) );
  nnd3s1 U1561 ( .DIN1(n1730), .DIN2(n1731), .DIN3(n1732), .Q(\IFinst/N85 ) );
  nnd2s1 U1562 ( .DIN1(n804), .DIN2(n246), .Q(n1732) );
  nnd2s1 U1563 ( .DIN1(n1733), .DIN2(n647), .Q(n1731) );
  xnr2s1 U1564 ( .DIN1(n1734), .DIN2(\NPC[13] ), .Q(n1733) );
  nnd2s1 U1565 ( .DIN1(n659), .DIN2(n9503), .Q(n1730) );
  nnd3s1 U1566 ( .DIN1(n1735), .DIN2(n1736), .DIN3(n1737), .Q(\IFinst/N84 ) );
  nnd2s1 U1567 ( .DIN1(n804), .DIN2(n245), .Q(n1737) );
  nnd2s1 U1568 ( .DIN1(n1738), .DIN2(n646), .Q(n1736) );
  xnr2s1 U1569 ( .DIN1(n9442), .DIN2(n1739), .Q(n1738) );
  nnd2s1 U1570 ( .DIN1(n658), .DIN2(n9502), .Q(n1735) );
  nnd3s1 U1571 ( .DIN1(n1740), .DIN2(n1741), .DIN3(n1742), .Q(\IFinst/N83 ) );
  nnd2s1 U1572 ( .DIN1(n804), .DIN2(n244), .Q(n1742) );
  nnd2s1 U1573 ( .DIN1(n1743), .DIN2(n645), .Q(n1741) );
  xnr2s1 U1574 ( .DIN1(n1744), .DIN2(\NPC[11] ), .Q(n1743) );
  nnd2s1 U1575 ( .DIN1(n657), .DIN2(n9501), .Q(n1740) );
  nnd3s1 U1576 ( .DIN1(n1745), .DIN2(n1746), .DIN3(n1747), .Q(\IFinst/N82 ) );
  nnd2s1 U1577 ( .DIN1(n1662), .DIN2(n243), .Q(n1747) );
  nnd2s1 U1578 ( .DIN1(n1748), .DIN2(n648), .Q(n1746) );
  xnr2s1 U1579 ( .DIN1(n9444), .DIN2(n1749), .Q(n1748) );
  nnd2s1 U1580 ( .DIN1(n660), .DIN2(n9500), .Q(n1745) );
  nnd3s1 U1581 ( .DIN1(n1750), .DIN2(n1751), .DIN3(n1752), .Q(\IFinst/N81 ) );
  nnd2s1 U1582 ( .DIN1(n1662), .DIN2(n242), .Q(n1752) );
  nnd2s1 U1583 ( .DIN1(n1753), .DIN2(n647), .Q(n1751) );
  xnr2s1 U1584 ( .DIN1(n1754), .DIN2(\NPC[9] ), .Q(n1753) );
  nnd2s1 U1585 ( .DIN1(n659), .DIN2(n9499), .Q(n1750) );
  nnd3s1 U1586 ( .DIN1(n1755), .DIN2(n1756), .DIN3(n1757), .Q(\IFinst/N80 ) );
  nnd2s1 U1587 ( .DIN1(n1662), .DIN2(n241), .Q(n1757) );
  nnd2s1 U1588 ( .DIN1(n1758), .DIN2(n646), .Q(n1756) );
  xnr2s1 U1589 ( .DIN1(n9446), .DIN2(n1759), .Q(n1758) );
  nnd2s1 U1590 ( .DIN1(n658), .DIN2(n9498), .Q(n1755) );
  nnd3s1 U1591 ( .DIN1(n1760), .DIN2(n1761), .DIN3(n1762), .Q(\IFinst/N79 ) );
  nnd2s1 U1592 ( .DIN1(n1662), .DIN2(n240), .Q(n1762) );
  nnd2s1 U1593 ( .DIN1(n1763), .DIN2(n645), .Q(n1761) );
  xnr2s1 U1594 ( .DIN1(n1764), .DIN2(\NPC[7] ), .Q(n1763) );
  nnd2s1 U1595 ( .DIN1(n657), .DIN2(n9497), .Q(n1760) );
  nnd3s1 U1596 ( .DIN1(n1765), .DIN2(n1766), .DIN3(n1767), .Q(\IFinst/N78 ) );
  nnd2s1 U1597 ( .DIN1(n1662), .DIN2(n239), .Q(n1767) );
  nnd2s1 U1598 ( .DIN1(n1768), .DIN2(n648), .Q(n1766) );
  xnr2s1 U1599 ( .DIN1(n9448), .DIN2(n1769), .Q(n1768) );
  nnd2s1 U1600 ( .DIN1(n660), .DIN2(n9496), .Q(n1765) );
  nnd3s1 U1601 ( .DIN1(n1770), .DIN2(n1771), .DIN3(n1772), .Q(\IFinst/N77 ) );
  nnd2s1 U1602 ( .DIN1(n1662), .DIN2(n238), .Q(n1772) );
  nnd2s1 U1603 ( .DIN1(n1773), .DIN2(n647), .Q(n1771) );
  xnr2s1 U1604 ( .DIN1(n1774), .DIN2(\NPC[5] ), .Q(n1773) );
  nnd2s1 U1605 ( .DIN1(n659), .DIN2(n9495), .Q(n1770) );
  nnd3s1 U1606 ( .DIN1(n1775), .DIN2(n1776), .DIN3(n1777), .Q(\IFinst/N76 ) );
  nnd2s1 U1607 ( .DIN1(n1662), .DIN2(n237), .Q(n1777) );
  nnd2s1 U1608 ( .DIN1(n1778), .DIN2(n646), .Q(n1776) );
  xnr2s1 U1609 ( .DIN1(n9450), .DIN2(n1779), .Q(n1778) );
  nnd2s1 U1610 ( .DIN1(n658), .DIN2(n9494), .Q(n1775) );
  nnd3s1 U1611 ( .DIN1(n1780), .DIN2(n1781), .DIN3(n1782), .Q(\IFinst/N75 ) );
  nnd2s1 U1612 ( .DIN1(n1662), .DIN2(n236), .Q(n1782) );
  nnd2s1 U1613 ( .DIN1(n648), .DIN2(n1783), .Q(n1781) );
  xnr2s1 U1614 ( .DIN1(\NPC[3] ), .DIN2(n9491), .Q(n1783) );
  nnd2s1 U1615 ( .DIN1(n657), .DIN2(n9493), .Q(n1780) );
  nnd3s1 U1616 ( .DIN1(n1784), .DIN2(n1785), .DIN3(n1786), .Q(\IFinst/N74 ) );
  nnd2s1 U1617 ( .DIN1(n1662), .DIN2(n235), .Q(n1786) );
  nnd2s1 U1618 ( .DIN1(n9491), .DIN2(n645), .Q(n1785) );
  nnd2s1 U1619 ( .DIN1(n660), .DIN2(n9492), .Q(n1784) );
  nnd3s1 U1620 ( .DIN1(n1787), .DIN2(n1470), .DIN3(n1788), .Q(\IFinst/N73 ) );
  nnd2s1 U1621 ( .DIN1(n1662), .DIN2(n234), .Q(n1788) );
  nnd2s1 U1622 ( .DIN1(n647), .DIN2(\IFinst/N8 ), .Q(n1470) );
  nnd2s1 U1623 ( .DIN1(n659), .DIN2(n9490), .Q(n1787) );
  nnd3s1 U1624 ( .DIN1(n1789), .DIN2(n1468), .DIN3(n1790), .Q(\IFinst/N72 ) );
  nnd2s1 U1625 ( .DIN1(n1662), .DIN2(n233), .Q(n1790) );
  nnd2s1 U1626 ( .DIN1(n646), .DIN2(\IFinst/N7 ), .Q(n1468) );
  nnd2s1 U1627 ( .DIN1(n658), .DIN2(n9523), .Q(n1789) );
  nnd3s1 U1628 ( .DIN1(n1791), .DIN2(n1792), .DIN3(n1793), .Q(\IFinst/N135 )
         );
  nnd2s1 U1629 ( .DIN1(n657), .DIN2(n9525), .Q(n1793) );
  nnd2s1 U1630 ( .DIN1(n780), .DIN2(n9524), .Q(n1792) );
  nnd2s1 U1631 ( .DIN1(\IR[31] ), .DIN2(n443), .Q(n1791) );
  nnd3s1 U1632 ( .DIN1(n1795), .DIN2(n1796), .DIN3(n1797), .Q(\IFinst/N134 )
         );
  nnd2s1 U1633 ( .DIN1(n660), .DIN2(n9527), .Q(n1797) );
  nnd2s1 U1634 ( .DIN1(n779), .DIN2(n9526), .Q(n1796) );
  nnd2s1 U1635 ( .DIN1(\IR[30] ), .DIN2(n442), .Q(n1795) );
  nnd3s1 U1636 ( .DIN1(n1798), .DIN2(n1799), .DIN3(n1800), .Q(\IFinst/N133 )
         );
  nnd2s1 U1637 ( .DIN1(n659), .DIN2(n9529), .Q(n1800) );
  nnd2s1 U1638 ( .DIN1(n780), .DIN2(n9528), .Q(n1799) );
  nnd2s1 U1639 ( .DIN1(\IR[29] ), .DIN2(n443), .Q(n1798) );
  nnd3s1 U1640 ( .DIN1(n1801), .DIN2(n1802), .DIN3(n1803), .Q(\IFinst/N132 )
         );
  nnd2s1 U1641 ( .DIN1(n658), .DIN2(n9531), .Q(n1803) );
  nnd2s1 U1642 ( .DIN1(n779), .DIN2(n9530), .Q(n1802) );
  nnd2s1 U1643 ( .DIN1(\IR[28] ), .DIN2(n442), .Q(n1801) );
  nnd3s1 U1644 ( .DIN1(n1804), .DIN2(n1805), .DIN3(n1806), .Q(\IFinst/N131 )
         );
  nnd2s1 U1645 ( .DIN1(n657), .DIN2(n9533), .Q(n1806) );
  nnd2s1 U1646 ( .DIN1(n780), .DIN2(n9532), .Q(n1805) );
  nnd2s1 U1647 ( .DIN1(\IR[27] ), .DIN2(n443), .Q(n1804) );
  nnd3s1 U1648 ( .DIN1(n1807), .DIN2(n1808), .DIN3(n1809), .Q(\IFinst/N130 )
         );
  nnd2s1 U1649 ( .DIN1(n660), .DIN2(n9535), .Q(n1809) );
  nnd2s1 U1650 ( .DIN1(n779), .DIN2(n9534), .Q(n1808) );
  nnd2s1 U1651 ( .DIN1(\IR[26] ), .DIN2(n442), .Q(n1807) );
  nnd3s1 U1652 ( .DIN1(n1810), .DIN2(n1811), .DIN3(n1812), .Q(\IFinst/N129 )
         );
  nnd2s1 U1653 ( .DIN1(n659), .DIN2(n9537), .Q(n1812) );
  nnd2s1 U1654 ( .DIN1(n780), .DIN2(n9536), .Q(n1811) );
  nnd2s1 U1655 ( .DIN1(\IR[25] ), .DIN2(n443), .Q(n1810) );
  nnd3s1 U1656 ( .DIN1(n1813), .DIN2(n1814), .DIN3(n1815), .Q(\IFinst/N128 )
         );
  nnd2s1 U1657 ( .DIN1(n658), .DIN2(n9539), .Q(n1815) );
  nnd2s1 U1658 ( .DIN1(n779), .DIN2(n9538), .Q(n1814) );
  nnd2s1 U1659 ( .DIN1(\IR[24] ), .DIN2(n442), .Q(n1813) );
  nnd3s1 U1660 ( .DIN1(n1816), .DIN2(n1817), .DIN3(n1818), .Q(\IFinst/N127 )
         );
  nnd2s1 U1661 ( .DIN1(n657), .DIN2(n9541), .Q(n1818) );
  nnd2s1 U1662 ( .DIN1(n780), .DIN2(n9540), .Q(n1817) );
  nnd2s1 U1663 ( .DIN1(\IR[23] ), .DIN2(n443), .Q(n1816) );
  nnd3s1 U1664 ( .DIN1(n1819), .DIN2(n1820), .DIN3(n1821), .Q(\IFinst/N126 )
         );
  nnd2s1 U1665 ( .DIN1(n660), .DIN2(n9543), .Q(n1821) );
  nnd2s1 U1666 ( .DIN1(n779), .DIN2(n9542), .Q(n1820) );
  nnd2s1 U1667 ( .DIN1(\IR[22] ), .DIN2(n442), .Q(n1819) );
  nnd3s1 U1668 ( .DIN1(n1822), .DIN2(n1823), .DIN3(n1824), .Q(\IFinst/N125 )
         );
  nnd2s1 U1669 ( .DIN1(n659), .DIN2(n9545), .Q(n1824) );
  nnd2s1 U1670 ( .DIN1(n780), .DIN2(n9544), .Q(n1823) );
  nnd2s1 U1671 ( .DIN1(\IR[21] ), .DIN2(n443), .Q(n1822) );
  nnd3s1 U1672 ( .DIN1(n1825), .DIN2(n1826), .DIN3(n1827), .Q(\IFinst/N124 )
         );
  nnd2s1 U1673 ( .DIN1(n658), .DIN2(n9547), .Q(n1827) );
  nnd2s1 U1674 ( .DIN1(n779), .DIN2(n9546), .Q(n1826) );
  nnd2s1 U1675 ( .DIN1(\IR[20] ), .DIN2(n442), .Q(n1825) );
  nnd3s1 U1676 ( .DIN1(n1828), .DIN2(n1829), .DIN3(n1830), .Q(\IFinst/N123 )
         );
  nnd2s1 U1677 ( .DIN1(n657), .DIN2(n9549), .Q(n1830) );
  nnd2s1 U1678 ( .DIN1(n780), .DIN2(n9548), .Q(n1829) );
  nnd2s1 U1679 ( .DIN1(\IR[19] ), .DIN2(n443), .Q(n1828) );
  nnd3s1 U1680 ( .DIN1(n1831), .DIN2(n1832), .DIN3(n1833), .Q(\IFinst/N122 )
         );
  nnd2s1 U1681 ( .DIN1(n660), .DIN2(n9551), .Q(n1833) );
  nnd2s1 U1682 ( .DIN1(n779), .DIN2(n9550), .Q(n1832) );
  nnd2s1 U1683 ( .DIN1(\IR[18] ), .DIN2(n442), .Q(n1831) );
  nnd3s1 U1684 ( .DIN1(n1834), .DIN2(n1835), .DIN3(n1836), .Q(\IFinst/N121 )
         );
  nnd2s1 U1685 ( .DIN1(n659), .DIN2(n9553), .Q(n1836) );
  nnd2s1 U1686 ( .DIN1(n780), .DIN2(n9552), .Q(n1835) );
  nnd2s1 U1687 ( .DIN1(\IR[17] ), .DIN2(n443), .Q(n1834) );
  nnd3s1 U1688 ( .DIN1(n1837), .DIN2(n1838), .DIN3(n1839), .Q(\IFinst/N120 )
         );
  nnd2s1 U1689 ( .DIN1(n658), .DIN2(n9555), .Q(n1839) );
  nnd2s1 U1690 ( .DIN1(n779), .DIN2(n9554), .Q(n1838) );
  nnd2s1 U1691 ( .DIN1(\IR[16] ), .DIN2(n442), .Q(n1837) );
  nnd3s1 U1692 ( .DIN1(n1840), .DIN2(n1841), .DIN3(n1842), .Q(\IFinst/N119 )
         );
  nnd2s1 U1693 ( .DIN1(n657), .DIN2(n9557), .Q(n1842) );
  nnd2s1 U1694 ( .DIN1(n780), .DIN2(n9556), .Q(n1841) );
  nnd2s1 U1695 ( .DIN1(\IR[15] ), .DIN2(n443), .Q(n1840) );
  nnd3s1 U1696 ( .DIN1(n1843), .DIN2(n1844), .DIN3(n1845), .Q(\IFinst/N118 )
         );
  nnd2s1 U1697 ( .DIN1(n660), .DIN2(n9559), .Q(n1845) );
  nnd2s1 U1698 ( .DIN1(n779), .DIN2(n9558), .Q(n1844) );
  nnd2s1 U1699 ( .DIN1(\IR[14] ), .DIN2(n442), .Q(n1843) );
  nnd3s1 U1700 ( .DIN1(n1846), .DIN2(n1847), .DIN3(n1848), .Q(\IFinst/N117 )
         );
  nnd2s1 U1701 ( .DIN1(n659), .DIN2(n9561), .Q(n1848) );
  nnd2s1 U1702 ( .DIN1(n780), .DIN2(n9560), .Q(n1847) );
  nnd2s1 U1703 ( .DIN1(\IR[13] ), .DIN2(n443), .Q(n1846) );
  nnd3s1 U1704 ( .DIN1(n1849), .DIN2(n1850), .DIN3(n1851), .Q(\IFinst/N116 )
         );
  nnd2s1 U1705 ( .DIN1(n658), .DIN2(n9563), .Q(n1851) );
  nnd2s1 U1706 ( .DIN1(n779), .DIN2(n9562), .Q(n1850) );
  nnd2s1 U1707 ( .DIN1(\IR[12] ), .DIN2(n442), .Q(n1849) );
  nnd3s1 U1708 ( .DIN1(n1852), .DIN2(n1853), .DIN3(n1854), .Q(\IFinst/N115 )
         );
  nnd2s1 U1709 ( .DIN1(n657), .DIN2(n9565), .Q(n1854) );
  nnd2s1 U1710 ( .DIN1(n780), .DIN2(n9564), .Q(n1853) );
  nnd2s1 U1711 ( .DIN1(\IR[11] ), .DIN2(n443), .Q(n1852) );
  nnd3s1 U1712 ( .DIN1(n1855), .DIN2(n1856), .DIN3(n1857), .Q(\IFinst/N114 )
         );
  nnd2s1 U1713 ( .DIN1(n660), .DIN2(n9567), .Q(n1857) );
  nnd2s1 U1714 ( .DIN1(n779), .DIN2(n9566), .Q(n1856) );
  nnd2s1 U1715 ( .DIN1(\IR[10] ), .DIN2(n442), .Q(n1855) );
  nnd3s1 U1716 ( .DIN1(n1858), .DIN2(n1859), .DIN3(n1860), .Q(\IFinst/N113 )
         );
  nnd2s1 U1717 ( .DIN1(n659), .DIN2(n9569), .Q(n1860) );
  nnd2s1 U1718 ( .DIN1(n780), .DIN2(n9568), .Q(n1859) );
  nnd2s1 U1719 ( .DIN1(\IR[9] ), .DIN2(n443), .Q(n1858) );
  nnd3s1 U1720 ( .DIN1(n1861), .DIN2(n1862), .DIN3(n1863), .Q(\IFinst/N112 )
         );
  nnd2s1 U1721 ( .DIN1(n658), .DIN2(n9571), .Q(n1863) );
  nnd2s1 U1722 ( .DIN1(n779), .DIN2(n9570), .Q(n1862) );
  nnd2s1 U1723 ( .DIN1(\IR[8] ), .DIN2(n442), .Q(n1861) );
  nnd3s1 U1724 ( .DIN1(n1864), .DIN2(n1865), .DIN3(n1866), .Q(\IFinst/N111 )
         );
  nnd2s1 U1725 ( .DIN1(n657), .DIN2(n9573), .Q(n1866) );
  nnd2s1 U1726 ( .DIN1(n780), .DIN2(n9572), .Q(n1865) );
  nnd2s1 U1727 ( .DIN1(\IR[7] ), .DIN2(n443), .Q(n1864) );
  nnd3s1 U1728 ( .DIN1(n1867), .DIN2(n1868), .DIN3(n1869), .Q(\IFinst/N110 )
         );
  nnd2s1 U1729 ( .DIN1(n660), .DIN2(n9575), .Q(n1869) );
  nnd2s1 U1730 ( .DIN1(n779), .DIN2(n9574), .Q(n1868) );
  nnd2s1 U1731 ( .DIN1(\IR[6] ), .DIN2(n442), .Q(n1867) );
  nnd3s1 U1732 ( .DIN1(n1870), .DIN2(n1871), .DIN3(n1872), .Q(\IFinst/N109 )
         );
  nnd2s1 U1733 ( .DIN1(n659), .DIN2(n9577), .Q(n1872) );
  nnd2s1 U1734 ( .DIN1(n780), .DIN2(n9576), .Q(n1871) );
  nnd2s1 U1735 ( .DIN1(\IR[5] ), .DIN2(n443), .Q(n1870) );
  nnd3s1 U1736 ( .DIN1(n1873), .DIN2(n1874), .DIN3(n1875), .Q(\IFinst/N108 )
         );
  nnd2s1 U1737 ( .DIN1(n658), .DIN2(n9579), .Q(n1875) );
  nnd2s1 U1738 ( .DIN1(n779), .DIN2(n9578), .Q(n1874) );
  nnd2s1 U1739 ( .DIN1(\IR[4] ), .DIN2(n442), .Q(n1873) );
  nnd3s1 U1740 ( .DIN1(n1876), .DIN2(n1877), .DIN3(n1878), .Q(\IFinst/N107 )
         );
  nnd2s1 U1741 ( .DIN1(n657), .DIN2(n9581), .Q(n1878) );
  nnd2s1 U1742 ( .DIN1(n780), .DIN2(n9580), .Q(n1877) );
  nnd2s1 U1743 ( .DIN1(\IR[3] ), .DIN2(n443), .Q(n1876) );
  nnd3s1 U1744 ( .DIN1(n1879), .DIN2(n1880), .DIN3(n1881), .Q(\IFinst/N106 )
         );
  nnd2s1 U1745 ( .DIN1(n660), .DIN2(n9583), .Q(n1881) );
  nnd2s1 U1746 ( .DIN1(n779), .DIN2(n9582), .Q(n1880) );
  nnd2s1 U1747 ( .DIN1(\IR[2] ), .DIN2(n442), .Q(n1879) );
  nnd3s1 U1748 ( .DIN1(n1882), .DIN2(n1883), .DIN3(n1884), .Q(\IFinst/N105 )
         );
  nnd2s1 U1749 ( .DIN1(n659), .DIN2(n9585), .Q(n1884) );
  nnd2s1 U1750 ( .DIN1(n780), .DIN2(n9584), .Q(n1883) );
  nnd2s1 U1751 ( .DIN1(\IR[1] ), .DIN2(n443), .Q(n1882) );
  nnd3s1 U1752 ( .DIN1(n1885), .DIN2(n1886), .DIN3(n1887), .Q(\IFinst/N104 )
         );
  nnd2s1 U1753 ( .DIN1(n658), .DIN2(n9587), .Q(n1887) );
  nnd2s1 U1754 ( .DIN1(n779), .DIN2(n9586), .Q(n1886) );
  nnd2s1 U1755 ( .DIN1(\IR[0] ), .DIN2(n442), .Q(n1885) );
  nnd2s1 U1756 ( .DIN1(n9383), .DIN2(n648), .Q(n1888) );
  nnd3s1 U1757 ( .DIN1(n1889), .DIN2(n1890), .DIN3(n1891), .Q(\IFinst/N103 )
         );
  or2s1 U1758 ( .DIN1(n9459), .DIN2(n9406), .Q(n1891) );
  nnd2s1 U1759 ( .DIN1(n1892), .DIN2(n647), .Q(n1890) );
  xnr2s1 U1760 ( .DIN1(n1893), .DIN2(\NPC[31] ), .Q(n1892) );
  nnd2s1 U1761 ( .DIN1(n1894), .DIN2(\NPC[30] ), .Q(n1893) );
  nnd2s1 U1762 ( .DIN1(n657), .DIN2(n9522), .Q(n1889) );
  nnd3s1 U1763 ( .DIN1(n1895), .DIN2(n1896), .DIN3(n1897), .Q(\IFinst/N102 )
         );
  nnd2s1 U1764 ( .DIN1(n1662), .DIN2(n263), .Q(n1897) );
  nnd2s1 U1765 ( .DIN1(n1898), .DIN2(n645), .Q(n1896) );
  xnr2s1 U1766 ( .DIN1(n9520), .DIN2(n1894), .Q(n1898) );
  nor2s1 U1767 ( .DIN1(n1899), .DIN2(n9425), .Q(n1894) );
  nnd2s1 U1768 ( .DIN1(n660), .DIN2(n9521), .Q(n1895) );
  nnd3s1 U1769 ( .DIN1(n1900), .DIN2(n1901), .DIN3(n1902), .Q(\IFinst/N101 )
         );
  nnd2s1 U1770 ( .DIN1(n1662), .DIN2(n262), .Q(n1902) );
  nnd2s1 U1771 ( .DIN1(n1903), .DIN2(n648), .Q(n1901) );
  xnr2s1 U1772 ( .DIN1(n1899), .DIN2(\NPC[29] ), .Q(n1903) );
  nnd2s1 U1773 ( .DIN1(n1904), .DIN2(\NPC[28] ), .Q(n1899) );
  nnd2s1 U1774 ( .DIN1(n659), .DIN2(n9519), .Q(n1900) );
  nnd3s1 U1775 ( .DIN1(n1905), .DIN2(n1906), .DIN3(n1907), .Q(\IFinst/N100 )
         );
  nnd2s1 U1776 ( .DIN1(n1662), .DIN2(n261), .Q(n1907) );
  nnd2s1 U1777 ( .DIN1(n1908), .DIN2(n647), .Q(n1906) );
  nor2s1 U1778 ( .DIN1(n1662), .DIN2(n685), .Q(n1466) );
  xnr2s1 U1779 ( .DIN1(n9426), .DIN2(n1904), .Q(n1908) );
  nor2s1 U1780 ( .DIN1(n1664), .DIN2(n9427), .Q(n1904) );
  nnd2s1 U1781 ( .DIN1(n1669), .DIN2(\NPC[26] ), .Q(n1664) );
  nor2s1 U1782 ( .DIN1(n1674), .DIN2(n9429), .Q(n1669) );
  nnd2s1 U1783 ( .DIN1(n1679), .DIN2(\NPC[24] ), .Q(n1674) );
  nor2s1 U1784 ( .DIN1(n1684), .DIN2(n9431), .Q(n1679) );
  nnd2s1 U1785 ( .DIN1(n1689), .DIN2(\NPC[22] ), .Q(n1684) );
  nor2s1 U1786 ( .DIN1(n1694), .DIN2(n9433), .Q(n1689) );
  nnd2s1 U1787 ( .DIN1(n1699), .DIN2(\NPC[20] ), .Q(n1694) );
  nor2s1 U1788 ( .DIN1(n1704), .DIN2(n9435), .Q(n1699) );
  nnd2s1 U1789 ( .DIN1(n1709), .DIN2(\NPC[18] ), .Q(n1704) );
  nor2s1 U1790 ( .DIN1(n1714), .DIN2(n9437), .Q(n1709) );
  nnd2s1 U1791 ( .DIN1(n1719), .DIN2(\NPC[16] ), .Q(n1714) );
  nor2s1 U1792 ( .DIN1(n1724), .DIN2(n9439), .Q(n1719) );
  nnd2s1 U1793 ( .DIN1(n1729), .DIN2(\NPC[14] ), .Q(n1724) );
  nor2s1 U1794 ( .DIN1(n1734), .DIN2(n9441), .Q(n1729) );
  nnd2s1 U1795 ( .DIN1(n1739), .DIN2(\NPC[12] ), .Q(n1734) );
  nor2s1 U1796 ( .DIN1(n1744), .DIN2(n9443), .Q(n1739) );
  nnd2s1 U1797 ( .DIN1(n1749), .DIN2(\NPC[10] ), .Q(n1744) );
  nor2s1 U1798 ( .DIN1(n1754), .DIN2(n9445), .Q(n1749) );
  nnd2s1 U1799 ( .DIN1(n1759), .DIN2(\NPC[8] ), .Q(n1754) );
  nor2s1 U1800 ( .DIN1(n1764), .DIN2(n9447), .Q(n1759) );
  nnd2s1 U1801 ( .DIN1(n1769), .DIN2(\NPC[6] ), .Q(n1764) );
  nor2s1 U1802 ( .DIN1(n1774), .DIN2(n9449), .Q(n1769) );
  nnd2s1 U1803 ( .DIN1(n1779), .DIN2(\NPC[4] ), .Q(n1774) );
  nor2s1 U1804 ( .DIN1(n9451), .DIN2(n9491), .Q(n1779) );
  nnd2s1 U1805 ( .DIN1(n658), .DIN2(n9518), .Q(n1905) );
  nnd2s1 U1806 ( .DIN1(n675), .DIN2(n1909), .Q(\IDinst/n5947 ) );
  nnd2s1 U1807 ( .DIN1(n1910), .DIN2(CLI), .Q(n1909) );
  nnd3s1 U1808 ( .DIN1(n677), .DIN2(n1910), .DIN3(n1911), .Q(\IDinst/n5946 )
         );
  nnd2s1 U1809 ( .DIN1(n1912), .DIN2(n215), .Q(n1911) );
  nnd2s1 U1810 ( .DIN1(n1913), .DIN2(n1914), .Q(n1912) );
  hi1s1 U1811 ( .DIN(n1915), .Q(n1913) );
  nnd2s1 U1812 ( .DIN1(n1916), .DIN2(n1917), .Q(\IDinst/n5945 ) );
  nnd4s1 U1813 ( .DIN1(n1914), .DIN2(n1918), .DIN3(n1919), .DIN4(n1920), 
        .Q(n1917) );
  and2s1 U1814 ( .DIN1(FREEZE), .DIN2(\IDinst/n1445 ), .Q(n1920) );
  nnd2s1 U1815 ( .DIN1(n441), .DIN2(n1921), .Q(n1916) );
  nor2s1 U1816 ( .DIN1(n1922), .DIN2(n383), .Q(\IDinst/n5944 ) );
  and2s1 U1817 ( .DIN1(n1923), .DIN2(n1924), .Q(n1922) );
  nnd2s1 U1818 ( .DIN1(n1925), .DIN2(n1926), .Q(\IDinst/n5943 ) );
  nnd2s1 U1819 ( .DIN1(n383), .DIN2(n323), .Q(n1926) );
  nnd2s1 U1820 ( .DIN1(n1927), .DIN2(n441), .Q(n1925) );
  nnd2s1 U1821 ( .DIN1(n1928), .DIN2(n1929), .Q(\IDinst/n5926 ) );
  nnd2s1 U1822 ( .DIN1(n382), .DIN2(n273), .Q(n1929) );
  nnd2s1 U1823 ( .DIN1(n1198), .DIN2(n329), .Q(n1928) );
  nnd2s1 U1824 ( .DIN1(n1930), .DIN2(n1931), .Q(\IDinst/n5925 ) );
  nnd2s1 U1825 ( .DIN1(n383), .DIN2(n275), .Q(n1931) );
  nnd2s1 U1826 ( .DIN1(n1312), .DIN2(n441), .Q(n1930) );
  nnd2s1 U1827 ( .DIN1(n1932), .DIN2(n1933), .Q(\IDinst/n5924 ) );
  nnd2s1 U1828 ( .DIN1(n382), .DIN2(n279), .Q(n1933) );
  nnd2s1 U1829 ( .DIN1(n1372), .DIN2(n329), .Q(n1932) );
  nnd2s1 U1830 ( .DIN1(n1934), .DIN2(n1935), .Q(\IDinst/n5923 ) );
  nnd2s1 U1831 ( .DIN1(n383), .DIN2(n281), .Q(n1935) );
  nnd2s1 U1832 ( .DIN1(n667), .DIN2(n441), .Q(n1934) );
  nnd2s1 U1833 ( .DIN1(n1936), .DIN2(n1937), .Q(\IDinst/n5922 ) );
  nnd2s1 U1834 ( .DIN1(n382), .DIN2(n277), .Q(n1937) );
  nnd2s1 U1835 ( .DIN1(n535), .DIN2(n329), .Q(n1936) );
  nnd2s1 U1836 ( .DIN1(n1938), .DIN2(n1939), .Q(\IDinst/n5921 ) );
  nnd2s1 U1837 ( .DIN1(n383), .DIN2(n309), .Q(n1939) );
  nnd2s1 U1838 ( .DIN1(n1065), .DIN2(n441), .Q(n1938) );
  nnd2s1 U1839 ( .DIN1(n1940), .DIN2(n1941), .Q(\IDinst/n5920 ) );
  nnd2s1 U1840 ( .DIN1(n382), .DIN2(n307), .Q(n1941) );
  nnd2s1 U1841 ( .DIN1(n1153), .DIN2(n329), .Q(n1940) );
  nnd2s1 U1842 ( .DIN1(n1942), .DIN2(n1943), .Q(\IDinst/n5919 ) );
  nnd2s1 U1843 ( .DIN1(n383), .DIN2(n313), .Q(n1943) );
  nnd2s1 U1844 ( .DIN1(n1194), .DIN2(n441), .Q(n1942) );
  nnd2s1 U1845 ( .DIN1(n1944), .DIN2(n1945), .Q(\IDinst/n5918 ) );
  nnd2s1 U1846 ( .DIN1(n382), .DIN2(n315), .Q(n1945) );
  nnd2s1 U1847 ( .DIN1(n642), .DIN2(n329), .Q(n1944) );
  nnd2s1 U1848 ( .DIN1(n1946), .DIN2(n1947), .Q(\IDinst/n5917 ) );
  nnd2s1 U1849 ( .DIN1(n383), .DIN2(n311), .Q(n1947) );
  nnd2s1 U1850 ( .DIN1(n539), .DIN2(n441), .Q(n1946) );
  nnd2s1 U1851 ( .DIN1(n1948), .DIN2(n1949), .Q(\IDinst/n5916 ) );
  nnd2s1 U1852 ( .DIN1(n382), .DIN2(n319), .Q(n1949) );
  nnd2s1 U1853 ( .DIN1(n1950), .DIN2(n329), .Q(n1948) );
  nnd2s1 U1854 ( .DIN1(n1951), .DIN2(n1952), .Q(\IDinst/n5915 ) );
  nnd2s1 U1855 ( .DIN1(n383), .DIN2(n321), .Q(n1952) );
  nnd2s1 U1856 ( .DIN1(n1953), .DIN2(n441), .Q(n1951) );
  nnd2s1 U1857 ( .DIN1(n1954), .DIN2(n1955), .Q(\IDinst/n5914 ) );
  nnd2s1 U1858 ( .DIN1(n382), .DIN2(n325), .Q(n1955) );
  nnd2s1 U1859 ( .DIN1(n1956), .DIN2(n329), .Q(n1954) );
  nnd2s1 U1860 ( .DIN1(n1957), .DIN2(n1958), .Q(\IDinst/n5913 ) );
  nnd2s1 U1861 ( .DIN1(n383), .DIN2(n327), .Q(n1958) );
  nnd2s1 U1862 ( .DIN1(n1959), .DIN2(n441), .Q(n1957) );
  nnd2s1 U1863 ( .DIN1(n1960), .DIN2(n1961), .Q(\IDinst/n5912 ) );
  nnd2s1 U1864 ( .DIN1(n382), .DIN2(n317), .Q(n1961) );
  nnd2s1 U1865 ( .DIN1(n1962), .DIN2(n329), .Q(n1960) );
  nnd3s1 U1866 ( .DIN1(n1963), .DIN2(n1964), .DIN3(n1965), .Q(\IDinst/n5911 )
         );
  nnd2s1 U1867 ( .DIN1(n649), .DIN2(n232), .Q(n1965) );
  nnd2s1 U1868 ( .DIN1(n1966), .DIN2(n114), .Q(n1963) );
  nnd3s1 U1869 ( .DIN1(n1967), .DIN2(n1964), .DIN3(n1968), .Q(\IDinst/n5910 )
         );
  nnd2s1 U1870 ( .DIN1(n652), .DIN2(n231), .Q(n1968) );
  nnd2s1 U1871 ( .DIN1(n1966), .DIN2(n98), .Q(n1967) );
  nnd3s1 U1872 ( .DIN1(n1969), .DIN2(n1964), .DIN3(n1970), .Q(\IDinst/n5909 )
         );
  nnd2s1 U1873 ( .DIN1(n651), .DIN2(n230), .Q(n1970) );
  nnd2s1 U1874 ( .DIN1(n1966), .DIN2(n113), .Q(n1969) );
  nnd3s1 U1875 ( .DIN1(n1971), .DIN2(n1964), .DIN3(n1972), .Q(\IDinst/n5908 )
         );
  nnd2s1 U1876 ( .DIN1(n650), .DIN2(n50), .Q(n1972) );
  nnd2s1 U1877 ( .DIN1(n1966), .DIN2(n97), .Q(n1971) );
  nnd3s1 U1878 ( .DIN1(n1973), .DIN2(n1964), .DIN3(n1974), .Q(\IDinst/n5907 )
         );
  nnd2s1 U1879 ( .DIN1(n649), .DIN2(n142), .Q(n1974) );
  nnd2s1 U1880 ( .DIN1(n1966), .DIN2(n92), .Q(n1973) );
  nnd2s1 U1881 ( .DIN1(n1975), .DIN2(n1976), .Q(\IDinst/n5906 ) );
  nnd2s1 U1882 ( .DIN1(n563), .DIN2(n799), .Q(n1976) );
  nnd2s1 U1883 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][0] ), .Q(n1975) );
  nnd2s1 U1884 ( .DIN1(n1978), .DIN2(n1979), .Q(\IDinst/n5905 ) );
  nnd2s1 U1885 ( .DIN1(n562), .DIN2(n798), .Q(n1979) );
  nnd2s1 U1886 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][1] ), .Q(n1978) );
  nnd2s1 U1887 ( .DIN1(n1981), .DIN2(n1982), .Q(\IDinst/n5904 ) );
  nnd2s1 U1888 ( .DIN1(n563), .DIN2(n800), .Q(n1982) );
  nnd2s1 U1889 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][2] ), .Q(n1981) );
  nnd2s1 U1890 ( .DIN1(n1984), .DIN2(n1985), .Q(\IDinst/n5903 ) );
  nnd2s1 U1891 ( .DIN1(n562), .DIN2(n797), .Q(n1985) );
  nnd2s1 U1892 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][3] ), .Q(n1984) );
  nnd2s1 U1893 ( .DIN1(n1987), .DIN2(n1988), .Q(\IDinst/n5902 ) );
  nnd2s1 U1894 ( .DIN1(n563), .DIN2(n796), .Q(n1988) );
  nnd2s1 U1895 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][4] ), .Q(n1987) );
  nnd2s1 U1896 ( .DIN1(n1990), .DIN2(n1991), .Q(\IDinst/n5901 ) );
  nnd2s1 U1897 ( .DIN1(n562), .DIN2(n795), .Q(n1991) );
  nnd2s1 U1898 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][5] ), .Q(n1990) );
  nnd2s1 U1899 ( .DIN1(n1993), .DIN2(n1994), .Q(\IDinst/n5900 ) );
  nnd2s1 U1900 ( .DIN1(n563), .DIN2(n794), .Q(n1994) );
  nnd2s1 U1901 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][6] ), .Q(n1993) );
  nnd2s1 U1902 ( .DIN1(n1996), .DIN2(n1997), .Q(\IDinst/n5899 ) );
  nnd2s1 U1903 ( .DIN1(n562), .DIN2(n793), .Q(n1997) );
  nnd2s1 U1904 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][7] ), .Q(n1996) );
  nnd2s1 U1905 ( .DIN1(n1999), .DIN2(n2000), .Q(\IDinst/n5898 ) );
  nnd2s1 U1906 ( .DIN1(n561), .DIN2(n799), .Q(n2000) );
  nnd2s1 U1907 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][0] ), .Q(n1999) );
  nnd2s1 U1908 ( .DIN1(n2001), .DIN2(n2002), .Q(\IDinst/n5897 ) );
  nnd2s1 U1909 ( .DIN1(n560), .DIN2(n798), .Q(n2002) );
  nnd2s1 U1910 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][1] ), .Q(n2001) );
  nnd2s1 U1911 ( .DIN1(n2003), .DIN2(n2004), .Q(\IDinst/n5896 ) );
  nnd2s1 U1912 ( .DIN1(n561), .DIN2(n800), .Q(n2004) );
  nnd2s1 U1913 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][2] ), .Q(n2003) );
  nnd2s1 U1914 ( .DIN1(n2005), .DIN2(n2006), .Q(\IDinst/n5895 ) );
  nnd2s1 U1915 ( .DIN1(n560), .DIN2(n797), .Q(n2006) );
  nnd2s1 U1916 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][3] ), .Q(n2005) );
  nnd2s1 U1917 ( .DIN1(n2007), .DIN2(n2008), .Q(\IDinst/n5894 ) );
  nnd2s1 U1918 ( .DIN1(n561), .DIN2(n796), .Q(n2008) );
  nnd2s1 U1919 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][4] ), .Q(n2007) );
  nnd2s1 U1920 ( .DIN1(n2009), .DIN2(n2010), .Q(\IDinst/n5893 ) );
  nnd2s1 U1921 ( .DIN1(n560), .DIN2(n795), .Q(n2010) );
  nnd2s1 U1922 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][5] ), .Q(n2009) );
  nnd2s1 U1923 ( .DIN1(n2011), .DIN2(n2012), .Q(\IDinst/n5892 ) );
  nnd2s1 U1924 ( .DIN1(n561), .DIN2(n794), .Q(n2012) );
  nnd2s1 U1925 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][6] ), .Q(n2011) );
  nnd2s1 U1926 ( .DIN1(n2013), .DIN2(n2014), .Q(\IDinst/n5891 ) );
  nnd2s1 U1927 ( .DIN1(n560), .DIN2(n793), .Q(n2014) );
  nnd2s1 U1928 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][7] ), .Q(n2013) );
  nnd2s1 U1929 ( .DIN1(n2015), .DIN2(n2016), .Q(\IDinst/n5890 ) );
  nnd2s1 U1930 ( .DIN1(n559), .DIN2(n799), .Q(n2016) );
  nnd2s1 U1931 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][0] ), .Q(n2015) );
  nnd2s1 U1932 ( .DIN1(n2017), .DIN2(n2018), .Q(\IDinst/n5889 ) );
  nnd2s1 U1933 ( .DIN1(n558), .DIN2(n798), .Q(n2018) );
  nnd2s1 U1934 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][1] ), .Q(n2017) );
  nnd2s1 U1935 ( .DIN1(n2019), .DIN2(n2020), .Q(\IDinst/n5888 ) );
  nnd2s1 U1936 ( .DIN1(n559), .DIN2(n800), .Q(n2020) );
  nnd2s1 U1937 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][2] ), .Q(n2019) );
  nnd2s1 U1938 ( .DIN1(n2021), .DIN2(n2022), .Q(\IDinst/n5887 ) );
  nnd2s1 U1939 ( .DIN1(n558), .DIN2(n797), .Q(n2022) );
  nnd2s1 U1940 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][3] ), .Q(n2021) );
  nnd2s1 U1941 ( .DIN1(n2023), .DIN2(n2024), .Q(\IDinst/n5886 ) );
  nnd2s1 U1942 ( .DIN1(n559), .DIN2(n796), .Q(n2024) );
  nnd2s1 U1943 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][4] ), .Q(n2023) );
  nnd2s1 U1944 ( .DIN1(n2025), .DIN2(n2026), .Q(\IDinst/n5885 ) );
  nnd2s1 U1945 ( .DIN1(n558), .DIN2(n795), .Q(n2026) );
  nnd2s1 U1946 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][5] ), .Q(n2025) );
  nnd2s1 U1947 ( .DIN1(n2027), .DIN2(n2028), .Q(\IDinst/n5884 ) );
  nnd2s1 U1948 ( .DIN1(n559), .DIN2(n794), .Q(n2028) );
  nnd2s1 U1949 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][6] ), .Q(n2027) );
  nnd2s1 U1950 ( .DIN1(n2029), .DIN2(n2030), .Q(\IDinst/n5883 ) );
  nnd2s1 U1951 ( .DIN1(n558), .DIN2(n793), .Q(n2030) );
  nnd2s1 U1952 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][7] ), .Q(n2029) );
  nnd2s1 U1953 ( .DIN1(n2031), .DIN2(n2032), .Q(\IDinst/n5882 ) );
  nnd2s1 U1954 ( .DIN1(n557), .DIN2(n799), .Q(n2032) );
  nnd2s1 U1955 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][0] ), .Q(n2031) );
  nnd2s1 U1956 ( .DIN1(n2033), .DIN2(n2034), .Q(\IDinst/n5881 ) );
  nnd2s1 U1957 ( .DIN1(n556), .DIN2(n798), .Q(n2034) );
  nnd2s1 U1958 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][1] ), .Q(n2033) );
  nnd2s1 U1959 ( .DIN1(n2035), .DIN2(n2036), .Q(\IDinst/n5880 ) );
  nnd2s1 U1960 ( .DIN1(n557), .DIN2(n800), .Q(n2036) );
  nnd2s1 U1961 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][2] ), .Q(n2035) );
  nnd2s1 U1962 ( .DIN1(n2037), .DIN2(n2038), .Q(\IDinst/n5879 ) );
  nnd2s1 U1963 ( .DIN1(n556), .DIN2(n797), .Q(n2038) );
  nnd2s1 U1964 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][3] ), .Q(n2037) );
  nnd2s1 U1965 ( .DIN1(n2039), .DIN2(n2040), .Q(\IDinst/n5878 ) );
  nnd2s1 U1966 ( .DIN1(n557), .DIN2(n796), .Q(n2040) );
  nnd2s1 U1967 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][4] ), .Q(n2039) );
  nnd2s1 U1968 ( .DIN1(n2041), .DIN2(n2042), .Q(\IDinst/n5877 ) );
  nnd2s1 U1969 ( .DIN1(n556), .DIN2(n795), .Q(n2042) );
  nnd2s1 U1970 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][5] ), .Q(n2041) );
  nnd2s1 U1971 ( .DIN1(n2043), .DIN2(n2044), .Q(\IDinst/n5876 ) );
  nnd2s1 U1972 ( .DIN1(n557), .DIN2(n794), .Q(n2044) );
  nnd2s1 U1973 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][6] ), .Q(n2043) );
  nnd2s1 U1974 ( .DIN1(n2045), .DIN2(n2046), .Q(\IDinst/n5875 ) );
  nnd2s1 U1975 ( .DIN1(n556), .DIN2(n793), .Q(n2046) );
  nnd2s1 U1976 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][7] ), .Q(n2045) );
  nnd2s1 U1977 ( .DIN1(n2047), .DIN2(n2048), .Q(\IDinst/n5874 ) );
  nnd2s1 U1978 ( .DIN1(n571), .DIN2(n799), .Q(n2048) );
  nnd2s1 U1979 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][0] ), .Q(n2047) );
  nnd2s1 U1980 ( .DIN1(n2049), .DIN2(n2050), .Q(\IDinst/n5873 ) );
  nnd2s1 U1981 ( .DIN1(n570), .DIN2(n798), .Q(n2050) );
  nnd2s1 U1982 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][1] ), .Q(n2049) );
  nnd2s1 U1983 ( .DIN1(n2051), .DIN2(n2052), .Q(\IDinst/n5872 ) );
  nnd2s1 U1984 ( .DIN1(n571), .DIN2(n800), .Q(n2052) );
  nnd2s1 U1985 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][2] ), .Q(n2051) );
  nnd2s1 U1986 ( .DIN1(n2053), .DIN2(n2054), .Q(\IDinst/n5871 ) );
  nnd2s1 U1987 ( .DIN1(n570), .DIN2(n797), .Q(n2054) );
  nnd2s1 U1988 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][3] ), .Q(n2053) );
  nnd2s1 U1989 ( .DIN1(n2055), .DIN2(n2056), .Q(\IDinst/n5870 ) );
  nnd2s1 U1990 ( .DIN1(n571), .DIN2(n796), .Q(n2056) );
  nnd2s1 U1991 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][4] ), .Q(n2055) );
  nnd2s1 U1992 ( .DIN1(n2057), .DIN2(n2058), .Q(\IDinst/n5869 ) );
  nnd2s1 U1993 ( .DIN1(n570), .DIN2(n795), .Q(n2058) );
  nnd2s1 U1994 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][5] ), .Q(n2057) );
  nnd2s1 U1995 ( .DIN1(n2059), .DIN2(n2060), .Q(\IDinst/n5868 ) );
  nnd2s1 U1996 ( .DIN1(n571), .DIN2(n794), .Q(n2060) );
  nnd2s1 U1997 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][6] ), .Q(n2059) );
  nnd2s1 U1998 ( .DIN1(n2061), .DIN2(n2062), .Q(\IDinst/n5867 ) );
  nnd2s1 U1999 ( .DIN1(n570), .DIN2(n793), .Q(n2062) );
  nnd2s1 U2000 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][7] ), .Q(n2061) );
  nnd2s1 U2001 ( .DIN1(n2063), .DIN2(n2064), .Q(\IDinst/n5866 ) );
  nnd2s1 U2002 ( .DIN1(n569), .DIN2(n799), .Q(n2064) );
  nnd2s1 U2003 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][0] ), .Q(n2063) );
  nnd2s1 U2004 ( .DIN1(n2065), .DIN2(n2066), .Q(\IDinst/n5865 ) );
  nnd2s1 U2005 ( .DIN1(n568), .DIN2(n798), .Q(n2066) );
  nnd2s1 U2006 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][1] ), .Q(n2065) );
  nnd2s1 U2007 ( .DIN1(n2067), .DIN2(n2068), .Q(\IDinst/n5864 ) );
  nnd2s1 U2008 ( .DIN1(n569), .DIN2(n800), .Q(n2068) );
  nnd2s1 U2009 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][2] ), .Q(n2067) );
  nnd2s1 U2010 ( .DIN1(n2069), .DIN2(n2070), .Q(\IDinst/n5863 ) );
  nnd2s1 U2011 ( .DIN1(n568), .DIN2(n797), .Q(n2070) );
  nnd2s1 U2012 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][3] ), .Q(n2069) );
  nnd2s1 U2013 ( .DIN1(n2071), .DIN2(n2072), .Q(\IDinst/n5862 ) );
  nnd2s1 U2014 ( .DIN1(n569), .DIN2(n796), .Q(n2072) );
  nnd2s1 U2015 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][4] ), .Q(n2071) );
  nnd2s1 U2016 ( .DIN1(n2073), .DIN2(n2074), .Q(\IDinst/n5861 ) );
  nnd2s1 U2017 ( .DIN1(n568), .DIN2(n795), .Q(n2074) );
  nnd2s1 U2018 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][5] ), .Q(n2073) );
  nnd2s1 U2019 ( .DIN1(n2075), .DIN2(n2076), .Q(\IDinst/n5860 ) );
  nnd2s1 U2020 ( .DIN1(n569), .DIN2(n794), .Q(n2076) );
  nnd2s1 U2021 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][6] ), .Q(n2075) );
  nnd2s1 U2022 ( .DIN1(n2077), .DIN2(n2078), .Q(\IDinst/n5859 ) );
  nnd2s1 U2023 ( .DIN1(n568), .DIN2(n793), .Q(n2078) );
  nnd2s1 U2024 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][7] ), .Q(n2077) );
  nnd2s1 U2025 ( .DIN1(n2079), .DIN2(n2080), .Q(\IDinst/n5858 ) );
  nnd2s1 U2026 ( .DIN1(n567), .DIN2(n799), .Q(n2080) );
  nnd2s1 U2027 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][0] ), .Q(n2079) );
  nnd2s1 U2028 ( .DIN1(n2081), .DIN2(n2082), .Q(\IDinst/n5857 ) );
  nnd2s1 U2029 ( .DIN1(n566), .DIN2(n798), .Q(n2082) );
  nnd2s1 U2030 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][1] ), .Q(n2081) );
  nnd2s1 U2031 ( .DIN1(n2083), .DIN2(n2084), .Q(\IDinst/n5856 ) );
  nnd2s1 U2032 ( .DIN1(n567), .DIN2(n800), .Q(n2084) );
  nnd2s1 U2033 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][2] ), .Q(n2083) );
  nnd2s1 U2034 ( .DIN1(n2085), .DIN2(n2086), .Q(\IDinst/n5855 ) );
  nnd2s1 U2035 ( .DIN1(n566), .DIN2(n797), .Q(n2086) );
  nnd2s1 U2036 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][3] ), .Q(n2085) );
  nnd2s1 U2037 ( .DIN1(n2087), .DIN2(n2088), .Q(\IDinst/n5854 ) );
  nnd2s1 U2038 ( .DIN1(n567), .DIN2(n796), .Q(n2088) );
  nnd2s1 U2039 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][4] ), .Q(n2087) );
  nnd2s1 U2040 ( .DIN1(n2089), .DIN2(n2090), .Q(\IDinst/n5853 ) );
  nnd2s1 U2041 ( .DIN1(n566), .DIN2(n795), .Q(n2090) );
  nnd2s1 U2042 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][5] ), .Q(n2089) );
  nnd2s1 U2043 ( .DIN1(n2091), .DIN2(n2092), .Q(\IDinst/n5852 ) );
  nnd2s1 U2044 ( .DIN1(n567), .DIN2(n794), .Q(n2092) );
  nnd2s1 U2045 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][6] ), .Q(n2091) );
  nnd2s1 U2046 ( .DIN1(n2093), .DIN2(n2094), .Q(\IDinst/n5851 ) );
  nnd2s1 U2047 ( .DIN1(n566), .DIN2(n793), .Q(n2094) );
  nnd2s1 U2048 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][7] ), .Q(n2093) );
  nnd2s1 U2049 ( .DIN1(n2095), .DIN2(n2096), .Q(\IDinst/n5850 ) );
  nnd2s1 U2050 ( .DIN1(n565), .DIN2(n799), .Q(n2096) );
  nnd2s1 U2051 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][0] ), .Q(n2095) );
  nnd2s1 U2052 ( .DIN1(n2097), .DIN2(n2098), .Q(\IDinst/n5849 ) );
  nnd2s1 U2053 ( .DIN1(n564), .DIN2(n798), .Q(n2098) );
  nnd2s1 U2054 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][1] ), .Q(n2097) );
  nnd2s1 U2055 ( .DIN1(n2099), .DIN2(n2100), .Q(\IDinst/n5848 ) );
  nnd2s1 U2056 ( .DIN1(n565), .DIN2(n800), .Q(n2100) );
  nnd2s1 U2057 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][2] ), .Q(n2099) );
  nnd2s1 U2058 ( .DIN1(n2101), .DIN2(n2102), .Q(\IDinst/n5847 ) );
  nnd2s1 U2059 ( .DIN1(n564), .DIN2(n797), .Q(n2102) );
  nnd2s1 U2060 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][3] ), .Q(n2101) );
  nnd2s1 U2061 ( .DIN1(n2103), .DIN2(n2104), .Q(\IDinst/n5846 ) );
  nnd2s1 U2062 ( .DIN1(n565), .DIN2(n796), .Q(n2104) );
  nnd2s1 U2063 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][4] ), .Q(n2103) );
  nnd2s1 U2064 ( .DIN1(n2105), .DIN2(n2106), .Q(\IDinst/n5845 ) );
  nnd2s1 U2065 ( .DIN1(n564), .DIN2(n795), .Q(n2106) );
  nnd2s1 U2066 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][5] ), .Q(n2105) );
  nnd2s1 U2067 ( .DIN1(n2107), .DIN2(n2108), .Q(\IDinst/n5844 ) );
  nnd2s1 U2068 ( .DIN1(n565), .DIN2(n794), .Q(n2108) );
  nnd2s1 U2069 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][6] ), .Q(n2107) );
  nnd2s1 U2070 ( .DIN1(n2109), .DIN2(n2110), .Q(\IDinst/n5843 ) );
  nnd2s1 U2071 ( .DIN1(n564), .DIN2(n793), .Q(n2110) );
  nnd2s1 U2072 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][7] ), .Q(n2109) );
  nnd2s1 U2073 ( .DIN1(n2111), .DIN2(n2112), .Q(\IDinst/n5842 ) );
  nnd2s1 U2074 ( .DIN1(n579), .DIN2(n799), .Q(n2112) );
  nnd2s1 U2075 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][0] ), .Q(n2111) );
  nnd2s1 U2076 ( .DIN1(n2113), .DIN2(n2114), .Q(\IDinst/n5841 ) );
  nnd2s1 U2077 ( .DIN1(n578), .DIN2(n798), .Q(n2114) );
  nnd2s1 U2078 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][1] ), .Q(n2113) );
  nnd2s1 U2079 ( .DIN1(n2115), .DIN2(n2116), .Q(\IDinst/n5840 ) );
  nnd2s1 U2080 ( .DIN1(n579), .DIN2(n800), .Q(n2116) );
  nnd2s1 U2081 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][2] ), .Q(n2115) );
  nnd2s1 U2082 ( .DIN1(n2117), .DIN2(n2118), .Q(\IDinst/n5839 ) );
  nnd2s1 U2083 ( .DIN1(n578), .DIN2(n797), .Q(n2118) );
  nnd2s1 U2084 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][3] ), .Q(n2117) );
  nnd2s1 U2085 ( .DIN1(n2119), .DIN2(n2120), .Q(\IDinst/n5838 ) );
  nnd2s1 U2086 ( .DIN1(n579), .DIN2(n796), .Q(n2120) );
  nnd2s1 U2087 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][4] ), .Q(n2119) );
  nnd2s1 U2088 ( .DIN1(n2121), .DIN2(n2122), .Q(\IDinst/n5837 ) );
  nnd2s1 U2089 ( .DIN1(n578), .DIN2(n795), .Q(n2122) );
  nnd2s1 U2090 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][5] ), .Q(n2121) );
  nnd2s1 U2091 ( .DIN1(n2123), .DIN2(n2124), .Q(\IDinst/n5836 ) );
  nnd2s1 U2092 ( .DIN1(n579), .DIN2(n794), .Q(n2124) );
  nnd2s1 U2093 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][6] ), .Q(n2123) );
  nnd2s1 U2094 ( .DIN1(n2125), .DIN2(n2126), .Q(\IDinst/n5835 ) );
  nnd2s1 U2095 ( .DIN1(n578), .DIN2(n793), .Q(n2126) );
  nnd2s1 U2096 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][7] ), .Q(n2125) );
  nnd2s1 U2097 ( .DIN1(n2127), .DIN2(n2128), .Q(\IDinst/n5834 ) );
  nnd2s1 U2098 ( .DIN1(n577), .DIN2(n799), .Q(n2128) );
  nnd2s1 U2099 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][0] ), .Q(n2127) );
  nnd2s1 U2100 ( .DIN1(n2129), .DIN2(n2130), .Q(\IDinst/n5833 ) );
  nnd2s1 U2101 ( .DIN1(n576), .DIN2(n798), .Q(n2130) );
  nnd2s1 U2102 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][1] ), .Q(n2129) );
  nnd2s1 U2103 ( .DIN1(n2131), .DIN2(n2132), .Q(\IDinst/n5832 ) );
  nnd2s1 U2104 ( .DIN1(n577), .DIN2(n800), .Q(n2132) );
  nnd2s1 U2105 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][2] ), .Q(n2131) );
  nnd2s1 U2106 ( .DIN1(n2133), .DIN2(n2134), .Q(\IDinst/n5831 ) );
  nnd2s1 U2107 ( .DIN1(n576), .DIN2(n797), .Q(n2134) );
  nnd2s1 U2108 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][3] ), .Q(n2133) );
  nnd2s1 U2109 ( .DIN1(n2135), .DIN2(n2136), .Q(\IDinst/n5830 ) );
  nnd2s1 U2110 ( .DIN1(n577), .DIN2(n796), .Q(n2136) );
  nnd2s1 U2111 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][4] ), .Q(n2135) );
  nnd2s1 U2112 ( .DIN1(n2137), .DIN2(n2138), .Q(\IDinst/n5829 ) );
  nnd2s1 U2113 ( .DIN1(n576), .DIN2(n795), .Q(n2138) );
  nnd2s1 U2114 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][5] ), .Q(n2137) );
  nnd2s1 U2115 ( .DIN1(n2139), .DIN2(n2140), .Q(\IDinst/n5828 ) );
  nnd2s1 U2116 ( .DIN1(n577), .DIN2(n794), .Q(n2140) );
  nnd2s1 U2117 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][6] ), .Q(n2139) );
  nnd2s1 U2118 ( .DIN1(n2141), .DIN2(n2142), .Q(\IDinst/n5827 ) );
  nnd2s1 U2119 ( .DIN1(n576), .DIN2(n793), .Q(n2142) );
  nnd2s1 U2120 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][7] ), .Q(n2141) );
  nnd2s1 U2121 ( .DIN1(n2143), .DIN2(n2144), .Q(\IDinst/n5826 ) );
  nnd2s1 U2122 ( .DIN1(n575), .DIN2(n799), .Q(n2144) );
  nnd2s1 U2123 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][0] ), .Q(n2143) );
  nnd2s1 U2124 ( .DIN1(n2145), .DIN2(n2146), .Q(\IDinst/n5825 ) );
  nnd2s1 U2125 ( .DIN1(n574), .DIN2(n798), .Q(n2146) );
  nnd2s1 U2126 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][1] ), .Q(n2145) );
  nnd2s1 U2127 ( .DIN1(n2147), .DIN2(n2148), .Q(\IDinst/n5824 ) );
  nnd2s1 U2128 ( .DIN1(n575), .DIN2(n800), .Q(n2148) );
  nnd2s1 U2129 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][2] ), .Q(n2147) );
  nnd2s1 U2130 ( .DIN1(n2149), .DIN2(n2150), .Q(\IDinst/n5823 ) );
  nnd2s1 U2131 ( .DIN1(n574), .DIN2(n797), .Q(n2150) );
  nnd2s1 U2132 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][3] ), .Q(n2149) );
  nnd2s1 U2133 ( .DIN1(n2151), .DIN2(n2152), .Q(\IDinst/n5822 ) );
  nnd2s1 U2134 ( .DIN1(n575), .DIN2(n796), .Q(n2152) );
  nnd2s1 U2135 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][4] ), .Q(n2151) );
  nnd2s1 U2136 ( .DIN1(n2153), .DIN2(n2154), .Q(\IDinst/n5821 ) );
  nnd2s1 U2137 ( .DIN1(n574), .DIN2(n795), .Q(n2154) );
  nnd2s1 U2138 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][5] ), .Q(n2153) );
  nnd2s1 U2139 ( .DIN1(n2155), .DIN2(n2156), .Q(\IDinst/n5820 ) );
  nnd2s1 U2140 ( .DIN1(n575), .DIN2(n794), .Q(n2156) );
  nnd2s1 U2141 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][6] ), .Q(n2155) );
  nnd2s1 U2142 ( .DIN1(n2157), .DIN2(n2158), .Q(\IDinst/n5819 ) );
  nnd2s1 U2143 ( .DIN1(n574), .DIN2(n793), .Q(n2158) );
  nnd2s1 U2144 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][7] ), .Q(n2157) );
  nnd2s1 U2145 ( .DIN1(n2159), .DIN2(n2160), .Q(\IDinst/n5818 ) );
  nnd2s1 U2146 ( .DIN1(n573), .DIN2(n799), .Q(n2160) );
  nnd2s1 U2147 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][0] ), .Q(n2159) );
  nnd2s1 U2148 ( .DIN1(n2161), .DIN2(n2162), .Q(\IDinst/n5817 ) );
  nnd2s1 U2149 ( .DIN1(n572), .DIN2(n798), .Q(n2162) );
  nnd2s1 U2150 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][1] ), .Q(n2161) );
  nnd2s1 U2151 ( .DIN1(n2163), .DIN2(n2164), .Q(\IDinst/n5816 ) );
  nnd2s1 U2152 ( .DIN1(n573), .DIN2(n800), .Q(n2164) );
  nnd2s1 U2153 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][2] ), .Q(n2163) );
  nnd2s1 U2154 ( .DIN1(n2165), .DIN2(n2166), .Q(\IDinst/n5815 ) );
  nnd2s1 U2155 ( .DIN1(n572), .DIN2(n797), .Q(n2166) );
  nnd2s1 U2156 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][3] ), .Q(n2165) );
  nnd2s1 U2157 ( .DIN1(n2167), .DIN2(n2168), .Q(\IDinst/n5814 ) );
  nnd2s1 U2158 ( .DIN1(n573), .DIN2(n796), .Q(n2168) );
  nnd2s1 U2159 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][4] ), .Q(n2167) );
  nnd2s1 U2160 ( .DIN1(n2169), .DIN2(n2170), .Q(\IDinst/n5813 ) );
  nnd2s1 U2161 ( .DIN1(n572), .DIN2(n795), .Q(n2170) );
  nnd2s1 U2162 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][5] ), .Q(n2169) );
  nnd2s1 U2163 ( .DIN1(n2171), .DIN2(n2172), .Q(\IDinst/n5812 ) );
  nnd2s1 U2164 ( .DIN1(n573), .DIN2(n794), .Q(n2172) );
  nnd2s1 U2165 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][6] ), .Q(n2171) );
  nnd2s1 U2166 ( .DIN1(n2173), .DIN2(n2174), .Q(\IDinst/n5811 ) );
  nnd2s1 U2167 ( .DIN1(n572), .DIN2(n793), .Q(n2174) );
  nnd2s1 U2168 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][7] ), .Q(n2173) );
  nnd2s1 U2169 ( .DIN1(n2175), .DIN2(n2176), .Q(\IDinst/n5810 ) );
  nnd2s1 U2170 ( .DIN1(n587), .DIN2(n799), .Q(n2176) );
  nnd2s1 U2171 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][0] ), .Q(n2175) );
  nnd2s1 U2172 ( .DIN1(n2177), .DIN2(n2178), .Q(\IDinst/n5809 ) );
  nnd2s1 U2173 ( .DIN1(n586), .DIN2(n798), .Q(n2178) );
  nnd2s1 U2174 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][1] ), .Q(n2177) );
  nnd2s1 U2175 ( .DIN1(n2179), .DIN2(n2180), .Q(\IDinst/n5808 ) );
  nnd2s1 U2176 ( .DIN1(n587), .DIN2(n800), .Q(n2180) );
  nnd2s1 U2177 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][2] ), .Q(n2179) );
  nnd2s1 U2178 ( .DIN1(n2181), .DIN2(n2182), .Q(\IDinst/n5807 ) );
  nnd2s1 U2179 ( .DIN1(n586), .DIN2(n797), .Q(n2182) );
  nnd2s1 U2180 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][3] ), .Q(n2181) );
  nnd2s1 U2181 ( .DIN1(n2183), .DIN2(n2184), .Q(\IDinst/n5806 ) );
  nnd2s1 U2182 ( .DIN1(n587), .DIN2(n796), .Q(n2184) );
  nnd2s1 U2183 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][4] ), .Q(n2183) );
  nnd2s1 U2184 ( .DIN1(n2185), .DIN2(n2186), .Q(\IDinst/n5805 ) );
  nnd2s1 U2185 ( .DIN1(n586), .DIN2(n795), .Q(n2186) );
  nnd2s1 U2186 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][5] ), .Q(n2185) );
  nnd2s1 U2187 ( .DIN1(n2187), .DIN2(n2188), .Q(\IDinst/n5804 ) );
  nnd2s1 U2188 ( .DIN1(n587), .DIN2(n794), .Q(n2188) );
  nnd2s1 U2189 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][6] ), .Q(n2187) );
  nnd2s1 U2190 ( .DIN1(n2189), .DIN2(n2190), .Q(\IDinst/n5803 ) );
  nnd2s1 U2191 ( .DIN1(n586), .DIN2(n793), .Q(n2190) );
  nnd2s1 U2192 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][7] ), .Q(n2189) );
  nnd2s1 U2193 ( .DIN1(n2191), .DIN2(n2192), .Q(\IDinst/n5802 ) );
  nnd2s1 U2194 ( .DIN1(n585), .DIN2(n799), .Q(n2192) );
  nnd2s1 U2195 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][0] ), .Q(n2191) );
  nnd2s1 U2196 ( .DIN1(n2193), .DIN2(n2194), .Q(\IDinst/n5801 ) );
  nnd2s1 U2197 ( .DIN1(n584), .DIN2(n798), .Q(n2194) );
  nnd2s1 U2198 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][1] ), .Q(n2193) );
  nnd2s1 U2199 ( .DIN1(n2195), .DIN2(n2196), .Q(\IDinst/n5800 ) );
  nnd2s1 U2200 ( .DIN1(n585), .DIN2(n800), .Q(n2196) );
  nnd2s1 U2201 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][2] ), .Q(n2195) );
  nnd2s1 U2202 ( .DIN1(n2197), .DIN2(n2198), .Q(\IDinst/n5799 ) );
  nnd2s1 U2203 ( .DIN1(n584), .DIN2(n797), .Q(n2198) );
  nnd2s1 U2204 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][3] ), .Q(n2197) );
  nnd2s1 U2205 ( .DIN1(n2199), .DIN2(n2200), .Q(\IDinst/n5798 ) );
  nnd2s1 U2206 ( .DIN1(n585), .DIN2(n796), .Q(n2200) );
  nnd2s1 U2207 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][4] ), .Q(n2199) );
  nnd2s1 U2208 ( .DIN1(n2201), .DIN2(n2202), .Q(\IDinst/n5797 ) );
  nnd2s1 U2209 ( .DIN1(n584), .DIN2(n795), .Q(n2202) );
  nnd2s1 U2210 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][5] ), .Q(n2201) );
  nnd2s1 U2211 ( .DIN1(n2203), .DIN2(n2204), .Q(\IDinst/n5796 ) );
  nnd2s1 U2212 ( .DIN1(n585), .DIN2(n794), .Q(n2204) );
  nnd2s1 U2213 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][6] ), .Q(n2203) );
  nnd2s1 U2214 ( .DIN1(n2205), .DIN2(n2206), .Q(\IDinst/n5795 ) );
  nnd2s1 U2215 ( .DIN1(n584), .DIN2(n793), .Q(n2206) );
  nnd2s1 U2216 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][7] ), .Q(n2205) );
  nnd2s1 U2217 ( .DIN1(n2207), .DIN2(n2208), .Q(\IDinst/n5794 ) );
  nnd2s1 U2218 ( .DIN1(n583), .DIN2(n799), .Q(n2208) );
  nnd2s1 U2219 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][0] ), .Q(n2207) );
  nnd2s1 U2220 ( .DIN1(n2209), .DIN2(n2210), .Q(\IDinst/n5793 ) );
  nnd2s1 U2221 ( .DIN1(n582), .DIN2(n798), .Q(n2210) );
  nnd2s1 U2222 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][1] ), .Q(n2209) );
  nnd2s1 U2223 ( .DIN1(n2211), .DIN2(n2212), .Q(\IDinst/n5792 ) );
  nnd2s1 U2224 ( .DIN1(n583), .DIN2(n800), .Q(n2212) );
  nnd2s1 U2225 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][2] ), .Q(n2211) );
  nnd2s1 U2226 ( .DIN1(n2213), .DIN2(n2214), .Q(\IDinst/n5791 ) );
  nnd2s1 U2227 ( .DIN1(n582), .DIN2(n797), .Q(n2214) );
  nnd2s1 U2228 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][3] ), .Q(n2213) );
  nnd2s1 U2229 ( .DIN1(n2215), .DIN2(n2216), .Q(\IDinst/n5790 ) );
  nnd2s1 U2230 ( .DIN1(n583), .DIN2(n796), .Q(n2216) );
  nnd2s1 U2231 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][4] ), .Q(n2215) );
  nnd2s1 U2232 ( .DIN1(n2217), .DIN2(n2218), .Q(\IDinst/n5789 ) );
  nnd2s1 U2233 ( .DIN1(n582), .DIN2(n795), .Q(n2218) );
  nnd2s1 U2234 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][5] ), .Q(n2217) );
  nnd2s1 U2235 ( .DIN1(n2219), .DIN2(n2220), .Q(\IDinst/n5788 ) );
  nnd2s1 U2236 ( .DIN1(n583), .DIN2(n794), .Q(n2220) );
  nnd2s1 U2237 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][6] ), .Q(n2219) );
  nnd2s1 U2238 ( .DIN1(n2221), .DIN2(n2222), .Q(\IDinst/n5787 ) );
  nnd2s1 U2239 ( .DIN1(n582), .DIN2(n793), .Q(n2222) );
  nnd2s1 U2240 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][7] ), .Q(n2221) );
  nnd2s1 U2241 ( .DIN1(n2223), .DIN2(n2224), .Q(\IDinst/n5786 ) );
  nnd2s1 U2242 ( .DIN1(n581), .DIN2(n799), .Q(n2224) );
  nnd2s1 U2243 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][0] ), .Q(n2223) );
  nnd2s1 U2244 ( .DIN1(n2225), .DIN2(n2226), .Q(\IDinst/n5785 ) );
  nnd2s1 U2245 ( .DIN1(n580), .DIN2(n798), .Q(n2226) );
  nnd2s1 U2246 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][1] ), .Q(n2225) );
  nnd2s1 U2247 ( .DIN1(n2227), .DIN2(n2228), .Q(\IDinst/n5784 ) );
  nnd2s1 U2248 ( .DIN1(n581), .DIN2(n800), .Q(n2228) );
  nnd2s1 U2249 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][2] ), .Q(n2227) );
  nnd2s1 U2250 ( .DIN1(n2229), .DIN2(n2230), .Q(\IDinst/n5783 ) );
  nnd2s1 U2251 ( .DIN1(n580), .DIN2(n797), .Q(n2230) );
  nnd2s1 U2252 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][3] ), .Q(n2229) );
  nnd2s1 U2253 ( .DIN1(n2231), .DIN2(n2232), .Q(\IDinst/n5782 ) );
  nnd2s1 U2254 ( .DIN1(n581), .DIN2(n796), .Q(n2232) );
  nnd2s1 U2255 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][4] ), .Q(n2231) );
  nnd2s1 U2256 ( .DIN1(n2233), .DIN2(n2234), .Q(\IDinst/n5781 ) );
  nnd2s1 U2257 ( .DIN1(n580), .DIN2(n795), .Q(n2234) );
  nnd2s1 U2258 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][5] ), .Q(n2233) );
  nnd2s1 U2259 ( .DIN1(n2235), .DIN2(n2236), .Q(\IDinst/n5780 ) );
  nnd2s1 U2260 ( .DIN1(n581), .DIN2(n794), .Q(n2236) );
  nnd2s1 U2261 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][6] ), .Q(n2235) );
  nnd2s1 U2262 ( .DIN1(n2237), .DIN2(n2238), .Q(\IDinst/n5779 ) );
  nnd2s1 U2263 ( .DIN1(n580), .DIN2(n793), .Q(n2238) );
  nnd2s1 U2264 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][7] ), .Q(n2237) );
  nnd2s1 U2265 ( .DIN1(n2239), .DIN2(n2240), .Q(\IDinst/n5778 ) );
  nnd2s1 U2266 ( .DIN1(n611), .DIN2(n799), .Q(n2240) );
  nnd2s1 U2267 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][0] ), .Q(n2239) );
  nnd2s1 U2268 ( .DIN1(n2241), .DIN2(n2242), .Q(\IDinst/n5777 ) );
  nnd2s1 U2269 ( .DIN1(n610), .DIN2(n798), .Q(n2242) );
  nnd2s1 U2270 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][1] ), .Q(n2241) );
  nnd2s1 U2271 ( .DIN1(n2243), .DIN2(n2244), .Q(\IDinst/n5776 ) );
  nnd2s1 U2272 ( .DIN1(n611), .DIN2(n800), .Q(n2244) );
  nnd2s1 U2273 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][2] ), .Q(n2243) );
  nnd2s1 U2274 ( .DIN1(n2245), .DIN2(n2246), .Q(\IDinst/n5775 ) );
  nnd2s1 U2275 ( .DIN1(n610), .DIN2(n797), .Q(n2246) );
  nnd2s1 U2276 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][3] ), .Q(n2245) );
  nnd2s1 U2277 ( .DIN1(n2247), .DIN2(n2248), .Q(\IDinst/n5774 ) );
  nnd2s1 U2278 ( .DIN1(n611), .DIN2(n796), .Q(n2248) );
  nnd2s1 U2279 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][4] ), .Q(n2247) );
  nnd2s1 U2280 ( .DIN1(n2249), .DIN2(n2250), .Q(\IDinst/n5773 ) );
  nnd2s1 U2281 ( .DIN1(n610), .DIN2(n795), .Q(n2250) );
  nnd2s1 U2282 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][5] ), .Q(n2249) );
  nnd2s1 U2283 ( .DIN1(n2251), .DIN2(n2252), .Q(\IDinst/n5772 ) );
  nnd2s1 U2284 ( .DIN1(n611), .DIN2(n794), .Q(n2252) );
  nnd2s1 U2285 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][6] ), .Q(n2251) );
  nnd2s1 U2286 ( .DIN1(n2253), .DIN2(n2254), .Q(\IDinst/n5771 ) );
  nnd2s1 U2287 ( .DIN1(n610), .DIN2(n793), .Q(n2254) );
  nnd2s1 U2288 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][7] ), .Q(n2253) );
  nnd2s1 U2289 ( .DIN1(n2255), .DIN2(n2256), .Q(\IDinst/n5770 ) );
  nnd2s1 U2290 ( .DIN1(n609), .DIN2(n1977), .Q(n2256) );
  nnd2s1 U2291 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][0] ), .Q(n2255) );
  nnd2s1 U2292 ( .DIN1(n2257), .DIN2(n2258), .Q(\IDinst/n5769 ) );
  nnd2s1 U2293 ( .DIN1(n608), .DIN2(n1980), .Q(n2258) );
  nnd2s1 U2294 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][1] ), .Q(n2257) );
  nnd2s1 U2295 ( .DIN1(n2259), .DIN2(n2260), .Q(\IDinst/n5768 ) );
  nnd2s1 U2296 ( .DIN1(n609), .DIN2(n1983), .Q(n2260) );
  nnd2s1 U2297 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][2] ), .Q(n2259) );
  nnd2s1 U2298 ( .DIN1(n2261), .DIN2(n2262), .Q(\IDinst/n5767 ) );
  nnd2s1 U2299 ( .DIN1(n608), .DIN2(n1986), .Q(n2262) );
  nnd2s1 U2300 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][3] ), .Q(n2261) );
  nnd2s1 U2301 ( .DIN1(n2263), .DIN2(n2264), .Q(\IDinst/n5766 ) );
  nnd2s1 U2302 ( .DIN1(n609), .DIN2(n1989), .Q(n2264) );
  nnd2s1 U2303 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][4] ), .Q(n2263) );
  nnd2s1 U2304 ( .DIN1(n2265), .DIN2(n2266), .Q(\IDinst/n5765 ) );
  nnd2s1 U2305 ( .DIN1(n608), .DIN2(n1992), .Q(n2266) );
  nnd2s1 U2306 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][5] ), .Q(n2265) );
  nnd2s1 U2307 ( .DIN1(n2267), .DIN2(n2268), .Q(\IDinst/n5764 ) );
  nnd2s1 U2308 ( .DIN1(n609), .DIN2(n1995), .Q(n2268) );
  nnd2s1 U2309 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][6] ), .Q(n2267) );
  nnd2s1 U2310 ( .DIN1(n2269), .DIN2(n2270), .Q(\IDinst/n5763 ) );
  nnd2s1 U2311 ( .DIN1(n608), .DIN2(n1998), .Q(n2270) );
  nnd2s1 U2312 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][7] ), .Q(n2269) );
  nnd2s1 U2313 ( .DIN1(n2271), .DIN2(n2272), .Q(\IDinst/n5762 ) );
  nnd2s1 U2314 ( .DIN1(n607), .DIN2(n1977), .Q(n2272) );
  nnd2s1 U2315 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][0] ), .Q(n2271) );
  nnd2s1 U2316 ( .DIN1(n2273), .DIN2(n2274), .Q(\IDinst/n5761 ) );
  nnd2s1 U2317 ( .DIN1(n606), .DIN2(n1980), .Q(n2274) );
  nnd2s1 U2318 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][1] ), .Q(n2273) );
  nnd2s1 U2319 ( .DIN1(n2275), .DIN2(n2276), .Q(\IDinst/n5760 ) );
  nnd2s1 U2320 ( .DIN1(n607), .DIN2(n1983), .Q(n2276) );
  nnd2s1 U2321 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][2] ), .Q(n2275) );
  nnd2s1 U2322 ( .DIN1(n2277), .DIN2(n2278), .Q(\IDinst/n5759 ) );
  nnd2s1 U2323 ( .DIN1(n606), .DIN2(n1986), .Q(n2278) );
  nnd2s1 U2324 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][3] ), .Q(n2277) );
  nnd2s1 U2325 ( .DIN1(n2279), .DIN2(n2280), .Q(\IDinst/n5758 ) );
  nnd2s1 U2326 ( .DIN1(n607), .DIN2(n1989), .Q(n2280) );
  nnd2s1 U2327 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][4] ), .Q(n2279) );
  nnd2s1 U2328 ( .DIN1(n2281), .DIN2(n2282), .Q(\IDinst/n5757 ) );
  nnd2s1 U2329 ( .DIN1(n606), .DIN2(n1992), .Q(n2282) );
  nnd2s1 U2330 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][5] ), .Q(n2281) );
  nnd2s1 U2331 ( .DIN1(n2283), .DIN2(n2284), .Q(\IDinst/n5756 ) );
  nnd2s1 U2332 ( .DIN1(n607), .DIN2(n1995), .Q(n2284) );
  nnd2s1 U2333 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][6] ), .Q(n2283) );
  nnd2s1 U2334 ( .DIN1(n2285), .DIN2(n2286), .Q(\IDinst/n5755 ) );
  nnd2s1 U2335 ( .DIN1(n606), .DIN2(n1998), .Q(n2286) );
  nnd2s1 U2336 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][7] ), .Q(n2285) );
  nnd2s1 U2337 ( .DIN1(n2287), .DIN2(n2288), .Q(\IDinst/n5754 ) );
  nnd2s1 U2338 ( .DIN1(n605), .DIN2(n1977), .Q(n2288) );
  nnd2s1 U2339 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][0] ), .Q(n2287) );
  nnd2s1 U2340 ( .DIN1(n2289), .DIN2(n2290), .Q(\IDinst/n5753 ) );
  nnd2s1 U2341 ( .DIN1(n604), .DIN2(n1980), .Q(n2290) );
  nnd2s1 U2342 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][1] ), .Q(n2289) );
  nnd2s1 U2343 ( .DIN1(n2291), .DIN2(n2292), .Q(\IDinst/n5752 ) );
  nnd2s1 U2344 ( .DIN1(n605), .DIN2(n1983), .Q(n2292) );
  nnd2s1 U2345 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][2] ), .Q(n2291) );
  nnd2s1 U2346 ( .DIN1(n2293), .DIN2(n2294), .Q(\IDinst/n5751 ) );
  nnd2s1 U2347 ( .DIN1(n604), .DIN2(n1986), .Q(n2294) );
  nnd2s1 U2348 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][3] ), .Q(n2293) );
  nnd2s1 U2349 ( .DIN1(n2295), .DIN2(n2296), .Q(\IDinst/n5750 ) );
  nnd2s1 U2350 ( .DIN1(n605), .DIN2(n1989), .Q(n2296) );
  nnd2s1 U2351 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][4] ), .Q(n2295) );
  nnd2s1 U2352 ( .DIN1(n2297), .DIN2(n2298), .Q(\IDinst/n5749 ) );
  nnd2s1 U2353 ( .DIN1(n604), .DIN2(n1992), .Q(n2298) );
  nnd2s1 U2354 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][5] ), .Q(n2297) );
  nnd2s1 U2355 ( .DIN1(n2299), .DIN2(n2300), .Q(\IDinst/n5748 ) );
  nnd2s1 U2356 ( .DIN1(n605), .DIN2(n1995), .Q(n2300) );
  nnd2s1 U2357 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][6] ), .Q(n2299) );
  nnd2s1 U2358 ( .DIN1(n2301), .DIN2(n2302), .Q(\IDinst/n5747 ) );
  nnd2s1 U2359 ( .DIN1(n604), .DIN2(n1998), .Q(n2302) );
  nnd2s1 U2360 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][7] ), .Q(n2301) );
  nnd2s1 U2361 ( .DIN1(n2303), .DIN2(n2304), .Q(\IDinst/n5746 ) );
  nnd2s1 U2362 ( .DIN1(n619), .DIN2(n1977), .Q(n2304) );
  nnd2s1 U2363 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][0] ), .Q(n2303) );
  nnd2s1 U2364 ( .DIN1(n2305), .DIN2(n2306), .Q(\IDinst/n5745 ) );
  nnd2s1 U2365 ( .DIN1(n618), .DIN2(n1980), .Q(n2306) );
  nnd2s1 U2366 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][1] ), .Q(n2305) );
  nnd2s1 U2367 ( .DIN1(n2307), .DIN2(n2308), .Q(\IDinst/n5744 ) );
  nnd2s1 U2368 ( .DIN1(n619), .DIN2(n1983), .Q(n2308) );
  nnd2s1 U2369 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][2] ), .Q(n2307) );
  nnd2s1 U2370 ( .DIN1(n2309), .DIN2(n2310), .Q(\IDinst/n5743 ) );
  nnd2s1 U2371 ( .DIN1(n618), .DIN2(n1986), .Q(n2310) );
  nnd2s1 U2372 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][3] ), .Q(n2309) );
  nnd2s1 U2373 ( .DIN1(n2311), .DIN2(n2312), .Q(\IDinst/n5742 ) );
  nnd2s1 U2374 ( .DIN1(n619), .DIN2(n1989), .Q(n2312) );
  nnd2s1 U2375 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][4] ), .Q(n2311) );
  nnd2s1 U2376 ( .DIN1(n2313), .DIN2(n2314), .Q(\IDinst/n5741 ) );
  nnd2s1 U2377 ( .DIN1(n618), .DIN2(n1992), .Q(n2314) );
  nnd2s1 U2378 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][5] ), .Q(n2313) );
  nnd2s1 U2379 ( .DIN1(n2315), .DIN2(n2316), .Q(\IDinst/n5740 ) );
  nnd2s1 U2380 ( .DIN1(n619), .DIN2(n1995), .Q(n2316) );
  nnd2s1 U2381 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][6] ), .Q(n2315) );
  nnd2s1 U2382 ( .DIN1(n2317), .DIN2(n2318), .Q(\IDinst/n5739 ) );
  nnd2s1 U2383 ( .DIN1(n618), .DIN2(n1998), .Q(n2318) );
  nnd2s1 U2384 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][7] ), .Q(n2317) );
  nnd2s1 U2385 ( .DIN1(n2319), .DIN2(n2320), .Q(\IDinst/n5738 ) );
  nnd2s1 U2386 ( .DIN1(n617), .DIN2(n1977), .Q(n2320) );
  nnd2s1 U2387 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][0] ), .Q(n2319) );
  nnd2s1 U2388 ( .DIN1(n2321), .DIN2(n2322), .Q(\IDinst/n5737 ) );
  nnd2s1 U2389 ( .DIN1(n616), .DIN2(n1980), .Q(n2322) );
  nnd2s1 U2390 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][1] ), .Q(n2321) );
  nnd2s1 U2391 ( .DIN1(n2323), .DIN2(n2324), .Q(\IDinst/n5736 ) );
  nnd2s1 U2392 ( .DIN1(n617), .DIN2(n1983), .Q(n2324) );
  nnd2s1 U2393 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][2] ), .Q(n2323) );
  nnd2s1 U2394 ( .DIN1(n2325), .DIN2(n2326), .Q(\IDinst/n5735 ) );
  nnd2s1 U2395 ( .DIN1(n616), .DIN2(n1986), .Q(n2326) );
  nnd2s1 U2396 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][3] ), .Q(n2325) );
  nnd2s1 U2397 ( .DIN1(n2327), .DIN2(n2328), .Q(\IDinst/n5734 ) );
  nnd2s1 U2398 ( .DIN1(n617), .DIN2(n1989), .Q(n2328) );
  nnd2s1 U2399 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][4] ), .Q(n2327) );
  nnd2s1 U2400 ( .DIN1(n2329), .DIN2(n2330), .Q(\IDinst/n5733 ) );
  nnd2s1 U2401 ( .DIN1(n616), .DIN2(n1992), .Q(n2330) );
  nnd2s1 U2402 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][5] ), .Q(n2329) );
  nnd2s1 U2403 ( .DIN1(n2331), .DIN2(n2332), .Q(\IDinst/n5732 ) );
  nnd2s1 U2404 ( .DIN1(n617), .DIN2(n1995), .Q(n2332) );
  nnd2s1 U2405 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][6] ), .Q(n2331) );
  nnd2s1 U2406 ( .DIN1(n2333), .DIN2(n2334), .Q(\IDinst/n5731 ) );
  nnd2s1 U2407 ( .DIN1(n616), .DIN2(n1998), .Q(n2334) );
  nnd2s1 U2408 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][7] ), .Q(n2333) );
  nnd2s1 U2409 ( .DIN1(n2335), .DIN2(n2336), .Q(\IDinst/n5730 ) );
  nnd2s1 U2410 ( .DIN1(n615), .DIN2(n1977), .Q(n2336) );
  nnd2s1 U2411 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][0] ), .Q(n2335) );
  nnd2s1 U2412 ( .DIN1(n2337), .DIN2(n2338), .Q(\IDinst/n5729 ) );
  nnd2s1 U2413 ( .DIN1(n614), .DIN2(n1980), .Q(n2338) );
  nnd2s1 U2414 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][1] ), .Q(n2337) );
  nnd2s1 U2415 ( .DIN1(n2339), .DIN2(n2340), .Q(\IDinst/n5728 ) );
  nnd2s1 U2416 ( .DIN1(n615), .DIN2(n1983), .Q(n2340) );
  nnd2s1 U2417 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][2] ), .Q(n2339) );
  nnd2s1 U2418 ( .DIN1(n2341), .DIN2(n2342), .Q(\IDinst/n5727 ) );
  nnd2s1 U2419 ( .DIN1(n614), .DIN2(n1986), .Q(n2342) );
  nnd2s1 U2420 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][3] ), .Q(n2341) );
  nnd2s1 U2421 ( .DIN1(n2343), .DIN2(n2344), .Q(\IDinst/n5726 ) );
  nnd2s1 U2422 ( .DIN1(n615), .DIN2(n1989), .Q(n2344) );
  nnd2s1 U2423 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][4] ), .Q(n2343) );
  nnd2s1 U2424 ( .DIN1(n2345), .DIN2(n2346), .Q(\IDinst/n5725 ) );
  nnd2s1 U2425 ( .DIN1(n614), .DIN2(n1992), .Q(n2346) );
  nnd2s1 U2426 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][5] ), .Q(n2345) );
  nnd2s1 U2427 ( .DIN1(n2347), .DIN2(n2348), .Q(\IDinst/n5724 ) );
  nnd2s1 U2428 ( .DIN1(n615), .DIN2(n1995), .Q(n2348) );
  nnd2s1 U2429 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][6] ), .Q(n2347) );
  nnd2s1 U2430 ( .DIN1(n2349), .DIN2(n2350), .Q(\IDinst/n5723 ) );
  nnd2s1 U2431 ( .DIN1(n614), .DIN2(n1998), .Q(n2350) );
  nnd2s1 U2432 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][7] ), .Q(n2349) );
  nnd2s1 U2433 ( .DIN1(n2351), .DIN2(n2352), .Q(\IDinst/n5722 ) );
  nnd2s1 U2434 ( .DIN1(n613), .DIN2(n1977), .Q(n2352) );
  nnd2s1 U2435 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][0] ), .Q(n2351) );
  nnd2s1 U2436 ( .DIN1(n2353), .DIN2(n2354), .Q(\IDinst/n5721 ) );
  nnd2s1 U2437 ( .DIN1(n612), .DIN2(n1980), .Q(n2354) );
  nnd2s1 U2438 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][1] ), .Q(n2353) );
  nnd2s1 U2439 ( .DIN1(n2355), .DIN2(n2356), .Q(\IDinst/n5720 ) );
  nnd2s1 U2440 ( .DIN1(n613), .DIN2(n1983), .Q(n2356) );
  nnd2s1 U2441 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][2] ), .Q(n2355) );
  nnd2s1 U2442 ( .DIN1(n2357), .DIN2(n2358), .Q(\IDinst/n5719 ) );
  nnd2s1 U2443 ( .DIN1(n612), .DIN2(n1986), .Q(n2358) );
  nnd2s1 U2444 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][3] ), .Q(n2357) );
  nnd2s1 U2445 ( .DIN1(n2359), .DIN2(n2360), .Q(\IDinst/n5718 ) );
  nnd2s1 U2446 ( .DIN1(n613), .DIN2(n1989), .Q(n2360) );
  nnd2s1 U2447 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][4] ), .Q(n2359) );
  nnd2s1 U2448 ( .DIN1(n2361), .DIN2(n2362), .Q(\IDinst/n5717 ) );
  nnd2s1 U2449 ( .DIN1(n612), .DIN2(n1992), .Q(n2362) );
  nnd2s1 U2450 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][5] ), .Q(n2361) );
  nnd2s1 U2451 ( .DIN1(n2363), .DIN2(n2364), .Q(\IDinst/n5716 ) );
  nnd2s1 U2452 ( .DIN1(n613), .DIN2(n1995), .Q(n2364) );
  nnd2s1 U2453 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][6] ), .Q(n2363) );
  nnd2s1 U2454 ( .DIN1(n2365), .DIN2(n2366), .Q(\IDinst/n5715 ) );
  nnd2s1 U2455 ( .DIN1(n612), .DIN2(n1998), .Q(n2366) );
  nnd2s1 U2456 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][7] ), .Q(n2365) );
  nnd2s1 U2457 ( .DIN1(n2367), .DIN2(n2368), .Q(\IDinst/n5714 ) );
  nnd2s1 U2458 ( .DIN1(n595), .DIN2(n1977), .Q(n2368) );
  nnd2s1 U2459 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][0] ), .Q(n2367) );
  nnd2s1 U2460 ( .DIN1(n2369), .DIN2(n2370), .Q(\IDinst/n5713 ) );
  nnd2s1 U2461 ( .DIN1(n594), .DIN2(n1980), .Q(n2370) );
  nnd2s1 U2462 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][1] ), .Q(n2369) );
  nnd2s1 U2463 ( .DIN1(n2371), .DIN2(n2372), .Q(\IDinst/n5712 ) );
  nnd2s1 U2464 ( .DIN1(n595), .DIN2(n1983), .Q(n2372) );
  nnd2s1 U2465 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][2] ), .Q(n2371) );
  nnd2s1 U2466 ( .DIN1(n2373), .DIN2(n2374), .Q(\IDinst/n5711 ) );
  nnd2s1 U2467 ( .DIN1(n594), .DIN2(n1986), .Q(n2374) );
  nnd2s1 U2468 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][3] ), .Q(n2373) );
  nnd2s1 U2469 ( .DIN1(n2375), .DIN2(n2376), .Q(\IDinst/n5710 ) );
  nnd2s1 U2470 ( .DIN1(n595), .DIN2(n1989), .Q(n2376) );
  nnd2s1 U2471 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][4] ), .Q(n2375) );
  nnd2s1 U2472 ( .DIN1(n2377), .DIN2(n2378), .Q(\IDinst/n5709 ) );
  nnd2s1 U2473 ( .DIN1(n594), .DIN2(n1992), .Q(n2378) );
  nnd2s1 U2474 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][5] ), .Q(n2377) );
  nnd2s1 U2475 ( .DIN1(n2379), .DIN2(n2380), .Q(\IDinst/n5708 ) );
  nnd2s1 U2476 ( .DIN1(n595), .DIN2(n1995), .Q(n2380) );
  nnd2s1 U2477 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][6] ), .Q(n2379) );
  nnd2s1 U2478 ( .DIN1(n2381), .DIN2(n2382), .Q(\IDinst/n5707 ) );
  nnd2s1 U2479 ( .DIN1(n594), .DIN2(n1998), .Q(n2382) );
  nnd2s1 U2480 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][7] ), .Q(n2381) );
  nnd2s1 U2481 ( .DIN1(n2383), .DIN2(n2384), .Q(\IDinst/n5706 ) );
  nnd2s1 U2482 ( .DIN1(n593), .DIN2(n1977), .Q(n2384) );
  nnd2s1 U2483 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][0] ), .Q(n2383) );
  nnd2s1 U2484 ( .DIN1(n2385), .DIN2(n2386), .Q(\IDinst/n5705 ) );
  nnd2s1 U2485 ( .DIN1(n592), .DIN2(n1980), .Q(n2386) );
  nnd2s1 U2486 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][1] ), .Q(n2385) );
  nnd2s1 U2487 ( .DIN1(n2387), .DIN2(n2388), .Q(\IDinst/n5704 ) );
  nnd2s1 U2488 ( .DIN1(n593), .DIN2(n1983), .Q(n2388) );
  nnd2s1 U2489 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][2] ), .Q(n2387) );
  nnd2s1 U2490 ( .DIN1(n2389), .DIN2(n2390), .Q(\IDinst/n5703 ) );
  nnd2s1 U2491 ( .DIN1(n592), .DIN2(n1986), .Q(n2390) );
  nnd2s1 U2492 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][3] ), .Q(n2389) );
  nnd2s1 U2493 ( .DIN1(n2391), .DIN2(n2392), .Q(\IDinst/n5702 ) );
  nnd2s1 U2494 ( .DIN1(n593), .DIN2(n1989), .Q(n2392) );
  nnd2s1 U2495 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][4] ), .Q(n2391) );
  nnd2s1 U2496 ( .DIN1(n2393), .DIN2(n2394), .Q(\IDinst/n5701 ) );
  nnd2s1 U2497 ( .DIN1(n592), .DIN2(n1992), .Q(n2394) );
  nnd2s1 U2498 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][5] ), .Q(n2393) );
  nnd2s1 U2499 ( .DIN1(n2395), .DIN2(n2396), .Q(\IDinst/n5700 ) );
  nnd2s1 U2500 ( .DIN1(n593), .DIN2(n1995), .Q(n2396) );
  nnd2s1 U2501 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][6] ), .Q(n2395) );
  nnd2s1 U2502 ( .DIN1(n2397), .DIN2(n2398), .Q(\IDinst/n5699 ) );
  nnd2s1 U2503 ( .DIN1(n592), .DIN2(n1998), .Q(n2398) );
  nnd2s1 U2504 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][7] ), .Q(n2397) );
  nnd2s1 U2505 ( .DIN1(n2399), .DIN2(n2400), .Q(\IDinst/n5698 ) );
  nnd2s1 U2506 ( .DIN1(n591), .DIN2(n1977), .Q(n2400) );
  nnd2s1 U2507 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][0] ), .Q(n2399) );
  nnd2s1 U2508 ( .DIN1(n2401), .DIN2(n2402), .Q(\IDinst/n5697 ) );
  nnd2s1 U2509 ( .DIN1(n590), .DIN2(n1980), .Q(n2402) );
  nnd2s1 U2510 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][1] ), .Q(n2401) );
  nnd2s1 U2511 ( .DIN1(n2403), .DIN2(n2404), .Q(\IDinst/n5696 ) );
  nnd2s1 U2512 ( .DIN1(n591), .DIN2(n1983), .Q(n2404) );
  nnd2s1 U2513 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][2] ), .Q(n2403) );
  nnd2s1 U2514 ( .DIN1(n2405), .DIN2(n2406), .Q(\IDinst/n5695 ) );
  nnd2s1 U2515 ( .DIN1(n590), .DIN2(n1986), .Q(n2406) );
  nnd2s1 U2516 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][3] ), .Q(n2405) );
  nnd2s1 U2517 ( .DIN1(n2407), .DIN2(n2408), .Q(\IDinst/n5694 ) );
  nnd2s1 U2518 ( .DIN1(n591), .DIN2(n1989), .Q(n2408) );
  nnd2s1 U2519 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][4] ), .Q(n2407) );
  nnd2s1 U2520 ( .DIN1(n2409), .DIN2(n2410), .Q(\IDinst/n5693 ) );
  nnd2s1 U2521 ( .DIN1(n590), .DIN2(n1992), .Q(n2410) );
  nnd2s1 U2522 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][5] ), .Q(n2409) );
  nnd2s1 U2523 ( .DIN1(n2411), .DIN2(n2412), .Q(\IDinst/n5692 ) );
  nnd2s1 U2524 ( .DIN1(n591), .DIN2(n1995), .Q(n2412) );
  nnd2s1 U2525 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][6] ), .Q(n2411) );
  nnd2s1 U2526 ( .DIN1(n2413), .DIN2(n2414), .Q(\IDinst/n5691 ) );
  nnd2s1 U2527 ( .DIN1(n590), .DIN2(n1998), .Q(n2414) );
  nnd2s1 U2528 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][7] ), .Q(n2413) );
  nnd2s1 U2529 ( .DIN1(n2415), .DIN2(n2416), .Q(\IDinst/n5690 ) );
  nnd2s1 U2530 ( .DIN1(n589), .DIN2(n1977), .Q(n2416) );
  nnd2s1 U2531 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][0] ), .Q(n2415) );
  nnd2s1 U2532 ( .DIN1(n2417), .DIN2(n2418), .Q(\IDinst/n5689 ) );
  nnd2s1 U2533 ( .DIN1(n588), .DIN2(n1980), .Q(n2418) );
  nnd2s1 U2534 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][1] ), .Q(n2417) );
  nnd2s1 U2535 ( .DIN1(n2419), .DIN2(n2420), .Q(\IDinst/n5688 ) );
  nnd2s1 U2536 ( .DIN1(n589), .DIN2(n1983), .Q(n2420) );
  nnd2s1 U2537 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][2] ), .Q(n2419) );
  nnd2s1 U2538 ( .DIN1(n2421), .DIN2(n2422), .Q(\IDinst/n5687 ) );
  nnd2s1 U2539 ( .DIN1(n588), .DIN2(n1986), .Q(n2422) );
  nnd2s1 U2540 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][3] ), .Q(n2421) );
  nnd2s1 U2541 ( .DIN1(n2423), .DIN2(n2424), .Q(\IDinst/n5686 ) );
  nnd2s1 U2542 ( .DIN1(n589), .DIN2(n1989), .Q(n2424) );
  nnd2s1 U2543 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][4] ), .Q(n2423) );
  nnd2s1 U2544 ( .DIN1(n2425), .DIN2(n2426), .Q(\IDinst/n5685 ) );
  nnd2s1 U2545 ( .DIN1(n588), .DIN2(n1992), .Q(n2426) );
  nnd2s1 U2546 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][5] ), .Q(n2425) );
  nnd2s1 U2547 ( .DIN1(n2427), .DIN2(n2428), .Q(\IDinst/n5684 ) );
  nnd2s1 U2548 ( .DIN1(n589), .DIN2(n1995), .Q(n2428) );
  nnd2s1 U2549 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][6] ), .Q(n2427) );
  nnd2s1 U2550 ( .DIN1(n2429), .DIN2(n2430), .Q(\IDinst/n5683 ) );
  nnd2s1 U2551 ( .DIN1(n588), .DIN2(n1998), .Q(n2430) );
  nnd2s1 U2552 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][7] ), .Q(n2429) );
  nnd2s1 U2553 ( .DIN1(n2431), .DIN2(n2432), .Q(\IDinst/n5682 ) );
  nnd2s1 U2554 ( .DIN1(n603), .DIN2(n1977), .Q(n2432) );
  nnd2s1 U2555 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][0] ), .Q(n2431) );
  nnd2s1 U2556 ( .DIN1(n2433), .DIN2(n2434), .Q(\IDinst/n5681 ) );
  nnd2s1 U2557 ( .DIN1(n602), .DIN2(n1980), .Q(n2434) );
  nnd2s1 U2558 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][1] ), .Q(n2433) );
  nnd2s1 U2559 ( .DIN1(n2435), .DIN2(n2436), .Q(\IDinst/n5680 ) );
  nnd2s1 U2560 ( .DIN1(n603), .DIN2(n1983), .Q(n2436) );
  nnd2s1 U2561 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][2] ), .Q(n2435) );
  nnd2s1 U2562 ( .DIN1(n2437), .DIN2(n2438), .Q(\IDinst/n5679 ) );
  nnd2s1 U2563 ( .DIN1(n602), .DIN2(n1986), .Q(n2438) );
  nnd2s1 U2564 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][3] ), .Q(n2437) );
  nnd2s1 U2565 ( .DIN1(n2439), .DIN2(n2440), .Q(\IDinst/n5678 ) );
  nnd2s1 U2566 ( .DIN1(n603), .DIN2(n1989), .Q(n2440) );
  nnd2s1 U2567 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][4] ), .Q(n2439) );
  nnd2s1 U2568 ( .DIN1(n2441), .DIN2(n2442), .Q(\IDinst/n5677 ) );
  nnd2s1 U2569 ( .DIN1(n602), .DIN2(n1992), .Q(n2442) );
  nnd2s1 U2570 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][5] ), .Q(n2441) );
  nnd2s1 U2571 ( .DIN1(n2443), .DIN2(n2444), .Q(\IDinst/n5676 ) );
  nnd2s1 U2572 ( .DIN1(n603), .DIN2(n1995), .Q(n2444) );
  nnd2s1 U2573 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][6] ), .Q(n2443) );
  nnd2s1 U2574 ( .DIN1(n2445), .DIN2(n2446), .Q(\IDinst/n5675 ) );
  nnd2s1 U2575 ( .DIN1(n602), .DIN2(n1998), .Q(n2446) );
  nnd2s1 U2576 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][7] ), .Q(n2445) );
  nnd2s1 U2577 ( .DIN1(n2447), .DIN2(n2448), .Q(\IDinst/n5674 ) );
  nnd2s1 U2578 ( .DIN1(n601), .DIN2(n1977), .Q(n2448) );
  nnd2s1 U2579 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][0] ), .Q(n2447) );
  nnd2s1 U2580 ( .DIN1(n2449), .DIN2(n2450), .Q(\IDinst/n5673 ) );
  nnd2s1 U2581 ( .DIN1(n600), .DIN2(n1980), .Q(n2450) );
  nnd2s1 U2582 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][1] ), .Q(n2449) );
  nnd2s1 U2583 ( .DIN1(n2451), .DIN2(n2452), .Q(\IDinst/n5672 ) );
  nnd2s1 U2584 ( .DIN1(n601), .DIN2(n1983), .Q(n2452) );
  nnd2s1 U2585 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][2] ), .Q(n2451) );
  nnd2s1 U2586 ( .DIN1(n2453), .DIN2(n2454), .Q(\IDinst/n5671 ) );
  nnd2s1 U2587 ( .DIN1(n600), .DIN2(n1986), .Q(n2454) );
  nnd2s1 U2588 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][3] ), .Q(n2453) );
  nnd2s1 U2589 ( .DIN1(n2455), .DIN2(n2456), .Q(\IDinst/n5670 ) );
  nnd2s1 U2590 ( .DIN1(n601), .DIN2(n1989), .Q(n2456) );
  nnd2s1 U2591 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][4] ), .Q(n2455) );
  nnd2s1 U2592 ( .DIN1(n2457), .DIN2(n2458), .Q(\IDinst/n5669 ) );
  nnd2s1 U2593 ( .DIN1(n600), .DIN2(n1992), .Q(n2458) );
  nnd2s1 U2594 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][5] ), .Q(n2457) );
  nnd2s1 U2595 ( .DIN1(n2459), .DIN2(n2460), .Q(\IDinst/n5668 ) );
  nnd2s1 U2596 ( .DIN1(n601), .DIN2(n1995), .Q(n2460) );
  nnd2s1 U2597 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][6] ), .Q(n2459) );
  nnd2s1 U2598 ( .DIN1(n2461), .DIN2(n2462), .Q(\IDinst/n5667 ) );
  nnd2s1 U2599 ( .DIN1(n600), .DIN2(n1998), .Q(n2462) );
  nnd2s1 U2600 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][7] ), .Q(n2461) );
  nnd2s1 U2601 ( .DIN1(n2463), .DIN2(n2464), .Q(\IDinst/n5666 ) );
  nnd2s1 U2602 ( .DIN1(n599), .DIN2(n1977), .Q(n2464) );
  nnd2s1 U2603 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][0] ), .Q(n2463) );
  nnd2s1 U2604 ( .DIN1(n2465), .DIN2(n2466), .Q(\IDinst/n5665 ) );
  nnd2s1 U2605 ( .DIN1(n598), .DIN2(n1980), .Q(n2466) );
  nnd2s1 U2606 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][1] ), .Q(n2465) );
  nnd2s1 U2607 ( .DIN1(n2467), .DIN2(n2468), .Q(\IDinst/n5664 ) );
  nnd2s1 U2608 ( .DIN1(n599), .DIN2(n1983), .Q(n2468) );
  nnd2s1 U2609 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][2] ), .Q(n2467) );
  nnd2s1 U2610 ( .DIN1(n2469), .DIN2(n2470), .Q(\IDinst/n5663 ) );
  nnd2s1 U2611 ( .DIN1(n598), .DIN2(n1986), .Q(n2470) );
  nnd2s1 U2612 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][3] ), .Q(n2469) );
  nnd2s1 U2613 ( .DIN1(n2471), .DIN2(n2472), .Q(\IDinst/n5662 ) );
  nnd2s1 U2614 ( .DIN1(n599), .DIN2(n1989), .Q(n2472) );
  nnd2s1 U2615 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][4] ), .Q(n2471) );
  nnd2s1 U2616 ( .DIN1(n2473), .DIN2(n2474), .Q(\IDinst/n5661 ) );
  nnd2s1 U2617 ( .DIN1(n598), .DIN2(n1992), .Q(n2474) );
  nnd2s1 U2618 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][5] ), .Q(n2473) );
  nnd2s1 U2619 ( .DIN1(n2475), .DIN2(n2476), .Q(\IDinst/n5660 ) );
  nnd2s1 U2620 ( .DIN1(n599), .DIN2(n1995), .Q(n2476) );
  nnd2s1 U2621 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][6] ), .Q(n2475) );
  nnd2s1 U2622 ( .DIN1(n2477), .DIN2(n2478), .Q(\IDinst/n5659 ) );
  nnd2s1 U2623 ( .DIN1(n598), .DIN2(n1998), .Q(n2478) );
  nnd2s1 U2624 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][7] ), .Q(n2477) );
  nnd2s1 U2625 ( .DIN1(n2479), .DIN2(n2480), .Q(\IDinst/n5658 ) );
  nnd2s1 U2626 ( .DIN1(n597), .DIN2(n1977), .Q(n2480) );
  nnd2s1 U2627 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][0] ), .Q(n2479) );
  nnd2s1 U2628 ( .DIN1(n2481), .DIN2(n2482), .Q(\IDinst/n5657 ) );
  nnd2s1 U2629 ( .DIN1(n596), .DIN2(n1980), .Q(n2482) );
  nnd2s1 U2630 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][1] ), .Q(n2481) );
  nnd2s1 U2631 ( .DIN1(n2483), .DIN2(n2484), .Q(\IDinst/n5656 ) );
  nnd2s1 U2632 ( .DIN1(n597), .DIN2(n1983), .Q(n2484) );
  nnd2s1 U2633 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][2] ), .Q(n2483) );
  nnd2s1 U2634 ( .DIN1(n2485), .DIN2(n2486), .Q(\IDinst/n5655 ) );
  nnd2s1 U2635 ( .DIN1(n596), .DIN2(n1986), .Q(n2486) );
  nnd2s1 U2636 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][3] ), .Q(n2485) );
  nnd2s1 U2637 ( .DIN1(n2487), .DIN2(n2488), .Q(\IDinst/n5654 ) );
  nnd2s1 U2638 ( .DIN1(n597), .DIN2(n1989), .Q(n2488) );
  nnd2s1 U2639 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][4] ), .Q(n2487) );
  nnd2s1 U2640 ( .DIN1(n2489), .DIN2(n2490), .Q(\IDinst/n5653 ) );
  nnd2s1 U2641 ( .DIN1(n596), .DIN2(n1992), .Q(n2490) );
  nnd2s1 U2642 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][5] ), .Q(n2489) );
  nnd2s1 U2643 ( .DIN1(n2491), .DIN2(n2492), .Q(\IDinst/n5652 ) );
  nnd2s1 U2644 ( .DIN1(n597), .DIN2(n1995), .Q(n2492) );
  nnd2s1 U2645 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][6] ), .Q(n2491) );
  nnd2s1 U2646 ( .DIN1(n2493), .DIN2(n2494), .Q(\IDinst/n5651 ) );
  nnd2s1 U2647 ( .DIN1(n596), .DIN2(n1998), .Q(n2494) );
  nnd2s1 U2648 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][7] ), .Q(n2493) );
  nnd2s1 U2649 ( .DIN1(n2495), .DIN2(n2496), .Q(\IDinst/n5650 ) );
  nnd2s1 U2650 ( .DIN1(n1950), .DIN2(n396), .Q(n2496) );
  nnd2s1 U2651 ( .DIN1(n652), .DIN2(IR_opcode_field[0]), .Q(n2495) );
  nnd2s1 U2652 ( .DIN1(n2497), .DIN2(n2498), .Q(\IDinst/n5649 ) );
  nnd2s1 U2653 ( .DIN1(n1953), .DIN2(n396), .Q(n2498) );
  nnd2s1 U2654 ( .DIN1(n651), .DIN2(IR_opcode_field[1]), .Q(n2497) );
  nnd2s1 U2655 ( .DIN1(n2499), .DIN2(n2500), .Q(\IDinst/n5648 ) );
  nnd2s1 U2656 ( .DIN1(n1956), .DIN2(n396), .Q(n2500) );
  nnd2s1 U2657 ( .DIN1(n650), .DIN2(IR_opcode_field[2]), .Q(n2499) );
  nnd2s1 U2658 ( .DIN1(n2501), .DIN2(n2502), .Q(\IDinst/n5647 ) );
  nnd2s1 U2659 ( .DIN1(n1959), .DIN2(n396), .Q(n2502) );
  nnd2s1 U2660 ( .DIN1(n649), .DIN2(IR_opcode_field[3]), .Q(n2501) );
  nnd2s1 U2661 ( .DIN1(n2503), .DIN2(n2504), .Q(\IDinst/n5646 ) );
  nnd2s1 U2662 ( .DIN1(n1962), .DIN2(n396), .Q(n2504) );
  nnd2s1 U2663 ( .DIN1(n652), .DIN2(IR_opcode_field[4]), .Q(n2503) );
  nnd2s1 U2664 ( .DIN1(n2505), .DIN2(n2506), .Q(\IDinst/n5645 ) );
  nnd2s1 U2665 ( .DIN1(n1927), .DIN2(n396), .Q(n2506) );
  nnd2s1 U2666 ( .DIN1(IR_opcode_field[5]), .DIN2(n651), .Q(n2505) );
  nnd2s1 U2667 ( .DIN1(n2507), .DIN2(n2508), .Q(\IDinst/n5644 ) );
  nnd2s1 U2668 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][8] ), .Q(n2508) );
  nnd2s1 U2669 ( .DIN1(n597), .DIN2(n693), .Q(n2507) );
  nnd2s1 U2670 ( .DIN1(n2510), .DIN2(n2511), .Q(\IDinst/n5643 ) );
  nnd2s1 U2671 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][8] ), .Q(n2511) );
  nnd2s1 U2672 ( .DIN1(n599), .DIN2(n693), .Q(n2510) );
  nnd2s1 U2673 ( .DIN1(n2512), .DIN2(n2513), .Q(\IDinst/n5642 ) );
  nnd2s1 U2674 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][8] ), .Q(n2513) );
  nnd2s1 U2675 ( .DIN1(n601), .DIN2(n693), .Q(n2512) );
  nnd2s1 U2676 ( .DIN1(n2514), .DIN2(n2515), .Q(\IDinst/n5641 ) );
  nnd2s1 U2677 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][8] ), .Q(n2515) );
  nnd2s1 U2678 ( .DIN1(n603), .DIN2(n693), .Q(n2514) );
  nnd2s1 U2679 ( .DIN1(n2516), .DIN2(n2517), .Q(\IDinst/n5640 ) );
  nnd2s1 U2680 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][8] ), .Q(n2517) );
  nnd2s1 U2681 ( .DIN1(n589), .DIN2(n693), .Q(n2516) );
  nnd2s1 U2682 ( .DIN1(n2518), .DIN2(n2519), .Q(\IDinst/n5639 ) );
  nnd2s1 U2683 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][8] ), .Q(n2519) );
  nnd2s1 U2684 ( .DIN1(n591), .DIN2(n693), .Q(n2518) );
  nnd2s1 U2685 ( .DIN1(n2520), .DIN2(n2521), .Q(\IDinst/n5638 ) );
  nnd2s1 U2686 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][8] ), .Q(n2521) );
  nnd2s1 U2687 ( .DIN1(n593), .DIN2(n693), .Q(n2520) );
  nnd2s1 U2688 ( .DIN1(n2522), .DIN2(n2523), .Q(\IDinst/n5637 ) );
  nnd2s1 U2689 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][8] ), .Q(n2523) );
  nnd2s1 U2690 ( .DIN1(n595), .DIN2(n693), .Q(n2522) );
  nnd2s1 U2691 ( .DIN1(n2524), .DIN2(n2525), .Q(\IDinst/n5636 ) );
  nnd2s1 U2692 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][8] ), .Q(n2525) );
  nnd2s1 U2693 ( .DIN1(n613), .DIN2(n693), .Q(n2524) );
  nnd2s1 U2694 ( .DIN1(n2526), .DIN2(n2527), .Q(\IDinst/n5635 ) );
  nnd2s1 U2695 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][8] ), .Q(n2527) );
  nnd2s1 U2696 ( .DIN1(n615), .DIN2(n693), .Q(n2526) );
  nnd2s1 U2697 ( .DIN1(n2528), .DIN2(n2529), .Q(\IDinst/n5634 ) );
  nnd2s1 U2698 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][8] ), .Q(n2529) );
  nnd2s1 U2699 ( .DIN1(n617), .DIN2(n693), .Q(n2528) );
  nnd2s1 U2700 ( .DIN1(n2530), .DIN2(n2531), .Q(\IDinst/n5633 ) );
  nnd2s1 U2701 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][8] ), .Q(n2531) );
  nnd2s1 U2702 ( .DIN1(n619), .DIN2(n693), .Q(n2530) );
  nnd2s1 U2703 ( .DIN1(n2532), .DIN2(n2533), .Q(\IDinst/n5632 ) );
  nnd2s1 U2704 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][8] ), .Q(n2533) );
  nnd2s1 U2705 ( .DIN1(n605), .DIN2(n693), .Q(n2532) );
  nnd2s1 U2706 ( .DIN1(n2534), .DIN2(n2535), .Q(\IDinst/n5631 ) );
  nnd2s1 U2707 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][8] ), .Q(n2535) );
  nnd2s1 U2708 ( .DIN1(n607), .DIN2(n2509), .Q(n2534) );
  nnd2s1 U2709 ( .DIN1(n2536), .DIN2(n2537), .Q(\IDinst/n5630 ) );
  nnd2s1 U2710 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][8] ), .Q(n2537) );
  nnd2s1 U2711 ( .DIN1(n609), .DIN2(n2509), .Q(n2536) );
  nnd2s1 U2712 ( .DIN1(n2538), .DIN2(n2539), .Q(\IDinst/n5629 ) );
  nnd2s1 U2713 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][8] ), .Q(n2539) );
  nnd2s1 U2714 ( .DIN1(n611), .DIN2(n2509), .Q(n2538) );
  nnd2s1 U2715 ( .DIN1(n2540), .DIN2(n2541), .Q(\IDinst/n5628 ) );
  nnd2s1 U2716 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][8] ), .Q(n2541) );
  nnd2s1 U2717 ( .DIN1(n581), .DIN2(n2509), .Q(n2540) );
  nnd2s1 U2718 ( .DIN1(n2542), .DIN2(n2543), .Q(\IDinst/n5627 ) );
  nnd2s1 U2719 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][8] ), .Q(n2543) );
  nnd2s1 U2720 ( .DIN1(n583), .DIN2(n2509), .Q(n2542) );
  nnd2s1 U2721 ( .DIN1(n2544), .DIN2(n2545), .Q(\IDinst/n5626 ) );
  nnd2s1 U2722 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][8] ), .Q(n2545) );
  nnd2s1 U2723 ( .DIN1(n585), .DIN2(n2509), .Q(n2544) );
  nnd2s1 U2724 ( .DIN1(n2546), .DIN2(n2547), .Q(\IDinst/n5625 ) );
  nnd2s1 U2725 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][8] ), .Q(n2547) );
  nnd2s1 U2726 ( .DIN1(n587), .DIN2(n2509), .Q(n2546) );
  nnd2s1 U2727 ( .DIN1(n2548), .DIN2(n2549), .Q(\IDinst/n5624 ) );
  nnd2s1 U2728 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][8] ), .Q(n2549) );
  nnd2s1 U2729 ( .DIN1(n573), .DIN2(n2509), .Q(n2548) );
  nnd2s1 U2730 ( .DIN1(n2550), .DIN2(n2551), .Q(\IDinst/n5623 ) );
  nnd2s1 U2731 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][8] ), .Q(n2551) );
  nnd2s1 U2732 ( .DIN1(n575), .DIN2(n2509), .Q(n2550) );
  nnd2s1 U2733 ( .DIN1(n2552), .DIN2(n2553), .Q(\IDinst/n5622 ) );
  nnd2s1 U2734 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][8] ), .Q(n2553) );
  nnd2s1 U2735 ( .DIN1(n577), .DIN2(n2509), .Q(n2552) );
  nnd2s1 U2736 ( .DIN1(n2554), .DIN2(n2555), .Q(\IDinst/n5621 ) );
  nnd2s1 U2737 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][8] ), .Q(n2555) );
  nnd2s1 U2738 ( .DIN1(n579), .DIN2(n2509), .Q(n2554) );
  nnd2s1 U2739 ( .DIN1(n2556), .DIN2(n2557), .Q(\IDinst/n5620 ) );
  nnd2s1 U2740 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][8] ), .Q(n2557) );
  nnd2s1 U2741 ( .DIN1(n565), .DIN2(n2509), .Q(n2556) );
  nnd2s1 U2742 ( .DIN1(n2558), .DIN2(n2559), .Q(\IDinst/n5619 ) );
  nnd2s1 U2743 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][8] ), .Q(n2559) );
  nnd2s1 U2744 ( .DIN1(n567), .DIN2(n2509), .Q(n2558) );
  nnd2s1 U2745 ( .DIN1(n2560), .DIN2(n2561), .Q(\IDinst/n5618 ) );
  nnd2s1 U2746 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][8] ), .Q(n2561) );
  nnd2s1 U2747 ( .DIN1(n569), .DIN2(n2509), .Q(n2560) );
  nnd2s1 U2748 ( .DIN1(n2562), .DIN2(n2563), .Q(\IDinst/n5617 ) );
  nnd2s1 U2749 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][8] ), .Q(n2563) );
  nnd2s1 U2750 ( .DIN1(n571), .DIN2(n2509), .Q(n2562) );
  nnd2s1 U2751 ( .DIN1(n2564), .DIN2(n2565), .Q(\IDinst/n5616 ) );
  nnd2s1 U2752 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][8] ), .Q(n2565) );
  nnd2s1 U2753 ( .DIN1(n557), .DIN2(n2509), .Q(n2564) );
  nnd2s1 U2754 ( .DIN1(n2566), .DIN2(n2567), .Q(\IDinst/n5615 ) );
  nnd2s1 U2755 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][8] ), .Q(n2567) );
  nnd2s1 U2756 ( .DIN1(n559), .DIN2(n2509), .Q(n2566) );
  nnd2s1 U2757 ( .DIN1(n2568), .DIN2(n2569), .Q(\IDinst/n5614 ) );
  nnd2s1 U2758 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][8] ), .Q(n2569) );
  nnd2s1 U2759 ( .DIN1(n561), .DIN2(n2509), .Q(n2568) );
  nnd2s1 U2760 ( .DIN1(n2570), .DIN2(n2571), .Q(\IDinst/n5613 ) );
  nnd2s1 U2761 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][8] ), .Q(n2571) );
  nnd2s1 U2762 ( .DIN1(n563), .DIN2(n2509), .Q(n2570) );
  nnd2s1 U2763 ( .DIN1(n2572), .DIN2(n2573), .Q(n2509) );
  nnd2s1 U2764 ( .DIN1(n2574), .DIN2(n200), .Q(n2573) );
  nnd2s1 U2765 ( .DIN1(n2575), .DIN2(n2576), .Q(\IDinst/n5612 ) );
  nnd2s1 U2766 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][9] ), .Q(n2576) );
  nnd2s1 U2767 ( .DIN1(n596), .DIN2(n697), .Q(n2575) );
  nnd2s1 U2768 ( .DIN1(n2578), .DIN2(n2579), .Q(\IDinst/n5611 ) );
  nnd2s1 U2769 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][9] ), .Q(n2579) );
  nnd2s1 U2770 ( .DIN1(n598), .DIN2(n697), .Q(n2578) );
  nnd2s1 U2771 ( .DIN1(n2580), .DIN2(n2581), .Q(\IDinst/n5610 ) );
  nnd2s1 U2772 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][9] ), .Q(n2581) );
  nnd2s1 U2773 ( .DIN1(n600), .DIN2(n697), .Q(n2580) );
  nnd2s1 U2774 ( .DIN1(n2582), .DIN2(n2583), .Q(\IDinst/n5609 ) );
  nnd2s1 U2775 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][9] ), .Q(n2583) );
  nnd2s1 U2776 ( .DIN1(n602), .DIN2(n697), .Q(n2582) );
  nnd2s1 U2777 ( .DIN1(n2584), .DIN2(n2585), .Q(\IDinst/n5608 ) );
  nnd2s1 U2778 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][9] ), .Q(n2585) );
  nnd2s1 U2779 ( .DIN1(n588), .DIN2(n697), .Q(n2584) );
  nnd2s1 U2780 ( .DIN1(n2586), .DIN2(n2587), .Q(\IDinst/n5607 ) );
  nnd2s1 U2781 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][9] ), .Q(n2587) );
  nnd2s1 U2782 ( .DIN1(n590), .DIN2(n697), .Q(n2586) );
  nnd2s1 U2783 ( .DIN1(n2588), .DIN2(n2589), .Q(\IDinst/n5606 ) );
  nnd2s1 U2784 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][9] ), .Q(n2589) );
  nnd2s1 U2785 ( .DIN1(n592), .DIN2(n697), .Q(n2588) );
  nnd2s1 U2786 ( .DIN1(n2590), .DIN2(n2591), .Q(\IDinst/n5605 ) );
  nnd2s1 U2787 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][9] ), .Q(n2591) );
  nnd2s1 U2788 ( .DIN1(n594), .DIN2(n697), .Q(n2590) );
  nnd2s1 U2789 ( .DIN1(n2592), .DIN2(n2593), .Q(\IDinst/n5604 ) );
  nnd2s1 U2790 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][9] ), .Q(n2593) );
  nnd2s1 U2791 ( .DIN1(n612), .DIN2(n697), .Q(n2592) );
  nnd2s1 U2792 ( .DIN1(n2594), .DIN2(n2595), .Q(\IDinst/n5603 ) );
  nnd2s1 U2793 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][9] ), .Q(n2595) );
  nnd2s1 U2794 ( .DIN1(n614), .DIN2(n697), .Q(n2594) );
  nnd2s1 U2795 ( .DIN1(n2596), .DIN2(n2597), .Q(\IDinst/n5602 ) );
  nnd2s1 U2796 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][9] ), .Q(n2597) );
  nnd2s1 U2797 ( .DIN1(n616), .DIN2(n697), .Q(n2596) );
  nnd2s1 U2798 ( .DIN1(n2598), .DIN2(n2599), .Q(\IDinst/n5601 ) );
  nnd2s1 U2799 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][9] ), .Q(n2599) );
  nnd2s1 U2800 ( .DIN1(n618), .DIN2(n697), .Q(n2598) );
  nnd2s1 U2801 ( .DIN1(n2600), .DIN2(n2601), .Q(\IDinst/n5600 ) );
  nnd2s1 U2802 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][9] ), .Q(n2601) );
  nnd2s1 U2803 ( .DIN1(n604), .DIN2(n697), .Q(n2600) );
  nnd2s1 U2804 ( .DIN1(n2602), .DIN2(n2603), .Q(\IDinst/n5599 ) );
  nnd2s1 U2805 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][9] ), .Q(n2603) );
  nnd2s1 U2806 ( .DIN1(n606), .DIN2(n2577), .Q(n2602) );
  nnd2s1 U2807 ( .DIN1(n2604), .DIN2(n2605), .Q(\IDinst/n5598 ) );
  nnd2s1 U2808 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][9] ), .Q(n2605) );
  nnd2s1 U2809 ( .DIN1(n608), .DIN2(n2577), .Q(n2604) );
  nnd2s1 U2810 ( .DIN1(n2606), .DIN2(n2607), .Q(\IDinst/n5597 ) );
  nnd2s1 U2811 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][9] ), .Q(n2607) );
  nnd2s1 U2812 ( .DIN1(n610), .DIN2(n2577), .Q(n2606) );
  nnd2s1 U2813 ( .DIN1(n2608), .DIN2(n2609), .Q(\IDinst/n5596 ) );
  nnd2s1 U2814 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][9] ), .Q(n2609) );
  nnd2s1 U2815 ( .DIN1(n580), .DIN2(n2577), .Q(n2608) );
  nnd2s1 U2816 ( .DIN1(n2610), .DIN2(n2611), .Q(\IDinst/n5595 ) );
  nnd2s1 U2817 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][9] ), .Q(n2611) );
  nnd2s1 U2818 ( .DIN1(n582), .DIN2(n2577), .Q(n2610) );
  nnd2s1 U2819 ( .DIN1(n2612), .DIN2(n2613), .Q(\IDinst/n5594 ) );
  nnd2s1 U2820 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][9] ), .Q(n2613) );
  nnd2s1 U2821 ( .DIN1(n584), .DIN2(n2577), .Q(n2612) );
  nnd2s1 U2822 ( .DIN1(n2614), .DIN2(n2615), .Q(\IDinst/n5593 ) );
  nnd2s1 U2823 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][9] ), .Q(n2615) );
  nnd2s1 U2824 ( .DIN1(n586), .DIN2(n2577), .Q(n2614) );
  nnd2s1 U2825 ( .DIN1(n2616), .DIN2(n2617), .Q(\IDinst/n5592 ) );
  nnd2s1 U2826 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][9] ), .Q(n2617) );
  nnd2s1 U2827 ( .DIN1(n572), .DIN2(n2577), .Q(n2616) );
  nnd2s1 U2828 ( .DIN1(n2618), .DIN2(n2619), .Q(\IDinst/n5591 ) );
  nnd2s1 U2829 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][9] ), .Q(n2619) );
  nnd2s1 U2830 ( .DIN1(n574), .DIN2(n2577), .Q(n2618) );
  nnd2s1 U2831 ( .DIN1(n2620), .DIN2(n2621), .Q(\IDinst/n5590 ) );
  nnd2s1 U2832 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][9] ), .Q(n2621) );
  nnd2s1 U2833 ( .DIN1(n576), .DIN2(n2577), .Q(n2620) );
  nnd2s1 U2834 ( .DIN1(n2622), .DIN2(n2623), .Q(\IDinst/n5589 ) );
  nnd2s1 U2835 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][9] ), .Q(n2623) );
  nnd2s1 U2836 ( .DIN1(n578), .DIN2(n2577), .Q(n2622) );
  nnd2s1 U2837 ( .DIN1(n2624), .DIN2(n2625), .Q(\IDinst/n5588 ) );
  nnd2s1 U2838 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][9] ), .Q(n2625) );
  nnd2s1 U2839 ( .DIN1(n564), .DIN2(n2577), .Q(n2624) );
  nnd2s1 U2840 ( .DIN1(n2626), .DIN2(n2627), .Q(\IDinst/n5587 ) );
  nnd2s1 U2841 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][9] ), .Q(n2627) );
  nnd2s1 U2842 ( .DIN1(n566), .DIN2(n2577), .Q(n2626) );
  nnd2s1 U2843 ( .DIN1(n2628), .DIN2(n2629), .Q(\IDinst/n5586 ) );
  nnd2s1 U2844 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][9] ), .Q(n2629) );
  nnd2s1 U2845 ( .DIN1(n568), .DIN2(n2577), .Q(n2628) );
  nnd2s1 U2846 ( .DIN1(n2630), .DIN2(n2631), .Q(\IDinst/n5585 ) );
  nnd2s1 U2847 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][9] ), .Q(n2631) );
  nnd2s1 U2848 ( .DIN1(n570), .DIN2(n2577), .Q(n2630) );
  nnd2s1 U2849 ( .DIN1(n2632), .DIN2(n2633), .Q(\IDinst/n5584 ) );
  nnd2s1 U2850 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][9] ), .Q(n2633) );
  nnd2s1 U2851 ( .DIN1(n556), .DIN2(n2577), .Q(n2632) );
  nnd2s1 U2852 ( .DIN1(n2634), .DIN2(n2635), .Q(\IDinst/n5583 ) );
  nnd2s1 U2853 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][9] ), .Q(n2635) );
  nnd2s1 U2854 ( .DIN1(n558), .DIN2(n2577), .Q(n2634) );
  nnd2s1 U2855 ( .DIN1(n2636), .DIN2(n2637), .Q(\IDinst/n5582 ) );
  nnd2s1 U2856 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][9] ), .Q(n2637) );
  nnd2s1 U2857 ( .DIN1(n560), .DIN2(n2577), .Q(n2636) );
  nnd2s1 U2858 ( .DIN1(n2638), .DIN2(n2639), .Q(\IDinst/n5581 ) );
  nnd2s1 U2859 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][9] ), .Q(n2639) );
  nnd2s1 U2860 ( .DIN1(n562), .DIN2(n2577), .Q(n2638) );
  nnd2s1 U2861 ( .DIN1(n2572), .DIN2(n2640), .Q(n2577) );
  nnd2s1 U2862 ( .DIN1(n2574), .DIN2(n198), .Q(n2640) );
  nnd2s1 U2863 ( .DIN1(n2641), .DIN2(n2642), .Q(\IDinst/n5580 ) );
  nnd2s1 U2864 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][10] ), .Q(n2642) );
  nnd2s1 U2865 ( .DIN1(n597), .DIN2(n702), .Q(n2641) );
  nnd2s1 U2866 ( .DIN1(n2644), .DIN2(n2645), .Q(\IDinst/n5579 ) );
  nnd2s1 U2867 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][10] ), .Q(n2645) );
  nnd2s1 U2868 ( .DIN1(n599), .DIN2(n702), .Q(n2644) );
  nnd2s1 U2869 ( .DIN1(n2646), .DIN2(n2647), .Q(\IDinst/n5578 ) );
  nnd2s1 U2870 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][10] ), .Q(n2647) );
  nnd2s1 U2871 ( .DIN1(n601), .DIN2(n702), .Q(n2646) );
  nnd2s1 U2872 ( .DIN1(n2648), .DIN2(n2649), .Q(\IDinst/n5577 ) );
  nnd2s1 U2873 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][10] ), .Q(n2649) );
  nnd2s1 U2874 ( .DIN1(n603), .DIN2(n702), .Q(n2648) );
  nnd2s1 U2875 ( .DIN1(n2650), .DIN2(n2651), .Q(\IDinst/n5576 ) );
  nnd2s1 U2876 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][10] ), .Q(n2651) );
  nnd2s1 U2877 ( .DIN1(n589), .DIN2(n702), .Q(n2650) );
  nnd2s1 U2878 ( .DIN1(n2652), .DIN2(n2653), .Q(\IDinst/n5575 ) );
  nnd2s1 U2879 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][10] ), .Q(n2653) );
  nnd2s1 U2880 ( .DIN1(n591), .DIN2(n702), .Q(n2652) );
  nnd2s1 U2881 ( .DIN1(n2654), .DIN2(n2655), .Q(\IDinst/n5574 ) );
  nnd2s1 U2882 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][10] ), .Q(n2655) );
  nnd2s1 U2883 ( .DIN1(n593), .DIN2(n702), .Q(n2654) );
  nnd2s1 U2884 ( .DIN1(n2656), .DIN2(n2657), .Q(\IDinst/n5573 ) );
  nnd2s1 U2885 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][10] ), .Q(n2657) );
  nnd2s1 U2886 ( .DIN1(n595), .DIN2(n702), .Q(n2656) );
  nnd2s1 U2887 ( .DIN1(n2658), .DIN2(n2659), .Q(\IDinst/n5572 ) );
  nnd2s1 U2888 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][10] ), .Q(n2659) );
  nnd2s1 U2889 ( .DIN1(n613), .DIN2(n702), .Q(n2658) );
  nnd2s1 U2890 ( .DIN1(n2660), .DIN2(n2661), .Q(\IDinst/n5571 ) );
  nnd2s1 U2891 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][10] ), .Q(n2661) );
  nnd2s1 U2892 ( .DIN1(n615), .DIN2(n702), .Q(n2660) );
  nnd2s1 U2893 ( .DIN1(n2662), .DIN2(n2663), .Q(\IDinst/n5570 ) );
  nnd2s1 U2894 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][10] ), .Q(n2663) );
  nnd2s1 U2895 ( .DIN1(n617), .DIN2(n702), .Q(n2662) );
  nnd2s1 U2896 ( .DIN1(n2664), .DIN2(n2665), .Q(\IDinst/n5569 ) );
  nnd2s1 U2897 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][10] ), .Q(n2665) );
  nnd2s1 U2898 ( .DIN1(n619), .DIN2(n702), .Q(n2664) );
  nnd2s1 U2899 ( .DIN1(n2666), .DIN2(n2667), .Q(\IDinst/n5568 ) );
  nnd2s1 U2900 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][10] ), .Q(n2667) );
  nnd2s1 U2901 ( .DIN1(n605), .DIN2(n702), .Q(n2666) );
  nnd2s1 U2902 ( .DIN1(n2668), .DIN2(n2669), .Q(\IDinst/n5567 ) );
  nnd2s1 U2903 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][10] ), .Q(n2669) );
  nnd2s1 U2904 ( .DIN1(n607), .DIN2(n2643), .Q(n2668) );
  nnd2s1 U2905 ( .DIN1(n2670), .DIN2(n2671), .Q(\IDinst/n5566 ) );
  nnd2s1 U2906 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][10] ), .Q(n2671) );
  nnd2s1 U2907 ( .DIN1(n609), .DIN2(n2643), .Q(n2670) );
  nnd2s1 U2908 ( .DIN1(n2672), .DIN2(n2673), .Q(\IDinst/n5565 ) );
  nnd2s1 U2909 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][10] ), .Q(n2673) );
  nnd2s1 U2910 ( .DIN1(n611), .DIN2(n2643), .Q(n2672) );
  nnd2s1 U2911 ( .DIN1(n2674), .DIN2(n2675), .Q(\IDinst/n5564 ) );
  nnd2s1 U2912 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][10] ), .Q(n2675) );
  nnd2s1 U2913 ( .DIN1(n581), .DIN2(n2643), .Q(n2674) );
  nnd2s1 U2914 ( .DIN1(n2676), .DIN2(n2677), .Q(\IDinst/n5563 ) );
  nnd2s1 U2915 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][10] ), .Q(n2677) );
  nnd2s1 U2916 ( .DIN1(n583), .DIN2(n2643), .Q(n2676) );
  nnd2s1 U2917 ( .DIN1(n2678), .DIN2(n2679), .Q(\IDinst/n5562 ) );
  nnd2s1 U2918 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][10] ), .Q(n2679) );
  nnd2s1 U2919 ( .DIN1(n585), .DIN2(n2643), .Q(n2678) );
  nnd2s1 U2920 ( .DIN1(n2680), .DIN2(n2681), .Q(\IDinst/n5561 ) );
  nnd2s1 U2921 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][10] ), .Q(n2681) );
  nnd2s1 U2922 ( .DIN1(n587), .DIN2(n2643), .Q(n2680) );
  nnd2s1 U2923 ( .DIN1(n2682), .DIN2(n2683), .Q(\IDinst/n5560 ) );
  nnd2s1 U2924 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][10] ), .Q(n2683) );
  nnd2s1 U2925 ( .DIN1(n573), .DIN2(n2643), .Q(n2682) );
  nnd2s1 U2926 ( .DIN1(n2684), .DIN2(n2685), .Q(\IDinst/n5559 ) );
  nnd2s1 U2927 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][10] ), .Q(n2685) );
  nnd2s1 U2928 ( .DIN1(n575), .DIN2(n2643), .Q(n2684) );
  nnd2s1 U2929 ( .DIN1(n2686), .DIN2(n2687), .Q(\IDinst/n5558 ) );
  nnd2s1 U2930 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][10] ), .Q(n2687) );
  nnd2s1 U2931 ( .DIN1(n577), .DIN2(n2643), .Q(n2686) );
  nnd2s1 U2932 ( .DIN1(n2688), .DIN2(n2689), .Q(\IDinst/n5557 ) );
  nnd2s1 U2933 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][10] ), .Q(n2689) );
  nnd2s1 U2934 ( .DIN1(n579), .DIN2(n2643), .Q(n2688) );
  nnd2s1 U2935 ( .DIN1(n2690), .DIN2(n2691), .Q(\IDinst/n5556 ) );
  nnd2s1 U2936 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][10] ), .Q(n2691) );
  nnd2s1 U2937 ( .DIN1(n565), .DIN2(n2643), .Q(n2690) );
  nnd2s1 U2938 ( .DIN1(n2692), .DIN2(n2693), .Q(\IDinst/n5555 ) );
  nnd2s1 U2939 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][10] ), .Q(n2693) );
  nnd2s1 U2940 ( .DIN1(n567), .DIN2(n2643), .Q(n2692) );
  nnd2s1 U2941 ( .DIN1(n2694), .DIN2(n2695), .Q(\IDinst/n5554 ) );
  nnd2s1 U2942 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][10] ), .Q(n2695) );
  nnd2s1 U2943 ( .DIN1(n569), .DIN2(n2643), .Q(n2694) );
  nnd2s1 U2944 ( .DIN1(n2696), .DIN2(n2697), .Q(\IDinst/n5553 ) );
  nnd2s1 U2945 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][10] ), .Q(n2697) );
  nnd2s1 U2946 ( .DIN1(n571), .DIN2(n2643), .Q(n2696) );
  nnd2s1 U2947 ( .DIN1(n2698), .DIN2(n2699), .Q(\IDinst/n5552 ) );
  nnd2s1 U2948 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][10] ), .Q(n2699) );
  nnd2s1 U2949 ( .DIN1(n557), .DIN2(n2643), .Q(n2698) );
  nnd2s1 U2950 ( .DIN1(n2700), .DIN2(n2701), .Q(\IDinst/n5551 ) );
  nnd2s1 U2951 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][10] ), .Q(n2701) );
  nnd2s1 U2952 ( .DIN1(n559), .DIN2(n2643), .Q(n2700) );
  nnd2s1 U2953 ( .DIN1(n2702), .DIN2(n2703), .Q(\IDinst/n5550 ) );
  nnd2s1 U2954 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][10] ), .Q(n2703) );
  nnd2s1 U2955 ( .DIN1(n561), .DIN2(n2643), .Q(n2702) );
  nnd2s1 U2956 ( .DIN1(n2704), .DIN2(n2705), .Q(\IDinst/n5549 ) );
  nnd2s1 U2957 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][10] ), .Q(n2705) );
  nnd2s1 U2958 ( .DIN1(n563), .DIN2(n2643), .Q(n2704) );
  nnd2s1 U2959 ( .DIN1(n2572), .DIN2(n2706), .Q(n2643) );
  nnd2s1 U2960 ( .DIN1(n2574), .DIN2(n196), .Q(n2706) );
  nnd2s1 U2961 ( .DIN1(n2707), .DIN2(n2708), .Q(\IDinst/n5548 ) );
  nnd2s1 U2962 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][11] ), .Q(n2708) );
  nnd2s1 U2963 ( .DIN1(n596), .DIN2(n708), .Q(n2707) );
  nnd2s1 U2964 ( .DIN1(n2710), .DIN2(n2711), .Q(\IDinst/n5547 ) );
  nnd2s1 U2965 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][11] ), .Q(n2711) );
  nnd2s1 U2966 ( .DIN1(n598), .DIN2(n2709), .Q(n2710) );
  nnd2s1 U2967 ( .DIN1(n2712), .DIN2(n2713), .Q(\IDinst/n5546 ) );
  nnd2s1 U2968 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][11] ), .Q(n2713) );
  nnd2s1 U2969 ( .DIN1(n600), .DIN2(n708), .Q(n2712) );
  nnd2s1 U2970 ( .DIN1(n2714), .DIN2(n2715), .Q(\IDinst/n5545 ) );
  nnd2s1 U2971 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][11] ), .Q(n2715) );
  nnd2s1 U2972 ( .DIN1(n602), .DIN2(n2709), .Q(n2714) );
  nnd2s1 U2973 ( .DIN1(n2716), .DIN2(n2717), .Q(\IDinst/n5544 ) );
  nnd2s1 U2974 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][11] ), .Q(n2717) );
  nnd2s1 U2975 ( .DIN1(n588), .DIN2(n708), .Q(n2716) );
  nnd2s1 U2976 ( .DIN1(n2718), .DIN2(n2719), .Q(\IDinst/n5543 ) );
  nnd2s1 U2977 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][11] ), .Q(n2719) );
  nnd2s1 U2978 ( .DIN1(n590), .DIN2(n2709), .Q(n2718) );
  nnd2s1 U2979 ( .DIN1(n2720), .DIN2(n2721), .Q(\IDinst/n5542 ) );
  nnd2s1 U2980 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][11] ), .Q(n2721) );
  nnd2s1 U2981 ( .DIN1(n592), .DIN2(n708), .Q(n2720) );
  nnd2s1 U2982 ( .DIN1(n2722), .DIN2(n2723), .Q(\IDinst/n5541 ) );
  nnd2s1 U2983 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][11] ), .Q(n2723) );
  nnd2s1 U2984 ( .DIN1(n594), .DIN2(n2709), .Q(n2722) );
  nnd2s1 U2985 ( .DIN1(n2724), .DIN2(n2725), .Q(\IDinst/n5540 ) );
  nnd2s1 U2986 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][11] ), .Q(n2725) );
  nnd2s1 U2987 ( .DIN1(n612), .DIN2(n708), .Q(n2724) );
  nnd2s1 U2988 ( .DIN1(n2726), .DIN2(n2727), .Q(\IDinst/n5539 ) );
  nnd2s1 U2989 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][11] ), .Q(n2727) );
  nnd2s1 U2990 ( .DIN1(n614), .DIN2(n2709), .Q(n2726) );
  nnd2s1 U2991 ( .DIN1(n2728), .DIN2(n2729), .Q(\IDinst/n5538 ) );
  nnd2s1 U2992 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][11] ), .Q(n2729) );
  nnd2s1 U2993 ( .DIN1(n616), .DIN2(n708), .Q(n2728) );
  nnd2s1 U2994 ( .DIN1(n2730), .DIN2(n2731), .Q(\IDinst/n5537 ) );
  nnd2s1 U2995 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][11] ), .Q(n2731) );
  nnd2s1 U2996 ( .DIN1(n618), .DIN2(n2709), .Q(n2730) );
  nnd2s1 U2997 ( .DIN1(n2732), .DIN2(n2733), .Q(\IDinst/n5536 ) );
  nnd2s1 U2998 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][11] ), .Q(n2733) );
  nnd2s1 U2999 ( .DIN1(n604), .DIN2(n708), .Q(n2732) );
  nnd2s1 U3000 ( .DIN1(n2734), .DIN2(n2735), .Q(\IDinst/n5535 ) );
  nnd2s1 U3001 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][11] ), .Q(n2735) );
  nnd2s1 U3002 ( .DIN1(n606), .DIN2(n2709), .Q(n2734) );
  nnd2s1 U3003 ( .DIN1(n2736), .DIN2(n2737), .Q(\IDinst/n5534 ) );
  nnd2s1 U3004 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][11] ), .Q(n2737) );
  nnd2s1 U3005 ( .DIN1(n608), .DIN2(n708), .Q(n2736) );
  nnd2s1 U3006 ( .DIN1(n2738), .DIN2(n2739), .Q(\IDinst/n5533 ) );
  nnd2s1 U3007 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][11] ), .Q(n2739) );
  nnd2s1 U3008 ( .DIN1(n610), .DIN2(n2709), .Q(n2738) );
  nnd2s1 U3009 ( .DIN1(n2740), .DIN2(n2741), .Q(\IDinst/n5532 ) );
  nnd2s1 U3010 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][11] ), .Q(n2741) );
  nnd2s1 U3011 ( .DIN1(n580), .DIN2(n708), .Q(n2740) );
  nnd2s1 U3012 ( .DIN1(n2742), .DIN2(n2743), .Q(\IDinst/n5531 ) );
  nnd2s1 U3013 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][11] ), .Q(n2743) );
  nnd2s1 U3014 ( .DIN1(n582), .DIN2(n2709), .Q(n2742) );
  nnd2s1 U3015 ( .DIN1(n2744), .DIN2(n2745), .Q(\IDinst/n5530 ) );
  nnd2s1 U3016 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][11] ), .Q(n2745) );
  nnd2s1 U3017 ( .DIN1(n584), .DIN2(n708), .Q(n2744) );
  nnd2s1 U3018 ( .DIN1(n2746), .DIN2(n2747), .Q(\IDinst/n5529 ) );
  nnd2s1 U3019 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][11] ), .Q(n2747) );
  nnd2s1 U3020 ( .DIN1(n586), .DIN2(n2709), .Q(n2746) );
  nnd2s1 U3021 ( .DIN1(n2748), .DIN2(n2749), .Q(\IDinst/n5528 ) );
  nnd2s1 U3022 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][11] ), .Q(n2749) );
  nnd2s1 U3023 ( .DIN1(n572), .DIN2(n708), .Q(n2748) );
  nnd2s1 U3024 ( .DIN1(n2750), .DIN2(n2751), .Q(\IDinst/n5527 ) );
  nnd2s1 U3025 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][11] ), .Q(n2751) );
  nnd2s1 U3026 ( .DIN1(n574), .DIN2(n2709), .Q(n2750) );
  nnd2s1 U3027 ( .DIN1(n2752), .DIN2(n2753), .Q(\IDinst/n5526 ) );
  nnd2s1 U3028 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][11] ), .Q(n2753) );
  nnd2s1 U3029 ( .DIN1(n576), .DIN2(n708), .Q(n2752) );
  nnd2s1 U3030 ( .DIN1(n2754), .DIN2(n2755), .Q(\IDinst/n5525 ) );
  nnd2s1 U3031 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][11] ), .Q(n2755) );
  nnd2s1 U3032 ( .DIN1(n578), .DIN2(n2709), .Q(n2754) );
  nnd2s1 U3033 ( .DIN1(n2756), .DIN2(n2757), .Q(\IDinst/n5524 ) );
  nnd2s1 U3034 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][11] ), .Q(n2757) );
  nnd2s1 U3035 ( .DIN1(n564), .DIN2(n708), .Q(n2756) );
  nnd2s1 U3036 ( .DIN1(n2758), .DIN2(n2759), .Q(\IDinst/n5523 ) );
  nnd2s1 U3037 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][11] ), .Q(n2759) );
  nnd2s1 U3038 ( .DIN1(n566), .DIN2(n2709), .Q(n2758) );
  nnd2s1 U3039 ( .DIN1(n2760), .DIN2(n2761), .Q(\IDinst/n5522 ) );
  nnd2s1 U3040 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][11] ), .Q(n2761) );
  nnd2s1 U3041 ( .DIN1(n568), .DIN2(n708), .Q(n2760) );
  nnd2s1 U3042 ( .DIN1(n2762), .DIN2(n2763), .Q(\IDinst/n5521 ) );
  nnd2s1 U3043 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][11] ), .Q(n2763) );
  nnd2s1 U3044 ( .DIN1(n570), .DIN2(n2709), .Q(n2762) );
  nnd2s1 U3045 ( .DIN1(n2764), .DIN2(n2765), .Q(\IDinst/n5520 ) );
  nnd2s1 U3046 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][11] ), .Q(n2765) );
  nnd2s1 U3047 ( .DIN1(n556), .DIN2(n708), .Q(n2764) );
  nnd2s1 U3048 ( .DIN1(n2766), .DIN2(n2767), .Q(\IDinst/n5519 ) );
  nnd2s1 U3049 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][11] ), .Q(n2767) );
  nnd2s1 U3050 ( .DIN1(n558), .DIN2(n2709), .Q(n2766) );
  nnd2s1 U3051 ( .DIN1(n2768), .DIN2(n2769), .Q(\IDinst/n5518 ) );
  nnd2s1 U3052 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][11] ), .Q(n2769) );
  nnd2s1 U3053 ( .DIN1(n560), .DIN2(n708), .Q(n2768) );
  nnd2s1 U3054 ( .DIN1(n2770), .DIN2(n2771), .Q(\IDinst/n5517 ) );
  nnd2s1 U3055 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][11] ), .Q(n2771) );
  nnd2s1 U3056 ( .DIN1(n562), .DIN2(n2709), .Q(n2770) );
  nnd2s1 U3057 ( .DIN1(n2572), .DIN2(n2772), .Q(n2709) );
  nnd2s1 U3058 ( .DIN1(n2574), .DIN2(n194), .Q(n2772) );
  nnd2s1 U3059 ( .DIN1(n2773), .DIN2(n2774), .Q(\IDinst/n5516 ) );
  nnd2s1 U3060 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][12] ), .Q(n2774) );
  nnd2s1 U3061 ( .DIN1(n597), .DIN2(n721), .Q(n2773) );
  nnd2s1 U3062 ( .DIN1(n2776), .DIN2(n2777), .Q(\IDinst/n5515 ) );
  nnd2s1 U3063 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][12] ), .Q(n2777) );
  nnd2s1 U3064 ( .DIN1(n599), .DIN2(n2775), .Q(n2776) );
  nnd2s1 U3065 ( .DIN1(n2778), .DIN2(n2779), .Q(\IDinst/n5514 ) );
  nnd2s1 U3066 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][12] ), .Q(n2779) );
  nnd2s1 U3067 ( .DIN1(n601), .DIN2(n721), .Q(n2778) );
  nnd2s1 U3068 ( .DIN1(n2780), .DIN2(n2781), .Q(\IDinst/n5513 ) );
  nnd2s1 U3069 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][12] ), .Q(n2781) );
  nnd2s1 U3070 ( .DIN1(n603), .DIN2(n2775), .Q(n2780) );
  nnd2s1 U3071 ( .DIN1(n2782), .DIN2(n2783), .Q(\IDinst/n5512 ) );
  nnd2s1 U3072 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][12] ), .Q(n2783) );
  nnd2s1 U3073 ( .DIN1(n589), .DIN2(n721), .Q(n2782) );
  nnd2s1 U3074 ( .DIN1(n2784), .DIN2(n2785), .Q(\IDinst/n5511 ) );
  nnd2s1 U3075 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][12] ), .Q(n2785) );
  nnd2s1 U3076 ( .DIN1(n591), .DIN2(n2775), .Q(n2784) );
  nnd2s1 U3077 ( .DIN1(n2786), .DIN2(n2787), .Q(\IDinst/n5510 ) );
  nnd2s1 U3078 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][12] ), .Q(n2787) );
  nnd2s1 U3079 ( .DIN1(n593), .DIN2(n721), .Q(n2786) );
  nnd2s1 U3080 ( .DIN1(n2788), .DIN2(n2789), .Q(\IDinst/n5509 ) );
  nnd2s1 U3081 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][12] ), .Q(n2789) );
  nnd2s1 U3082 ( .DIN1(n595), .DIN2(n2775), .Q(n2788) );
  nnd2s1 U3083 ( .DIN1(n2790), .DIN2(n2791), .Q(\IDinst/n5508 ) );
  nnd2s1 U3084 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][12] ), .Q(n2791) );
  nnd2s1 U3085 ( .DIN1(n613), .DIN2(n721), .Q(n2790) );
  nnd2s1 U3086 ( .DIN1(n2792), .DIN2(n2793), .Q(\IDinst/n5507 ) );
  nnd2s1 U3087 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][12] ), .Q(n2793) );
  nnd2s1 U3088 ( .DIN1(n615), .DIN2(n2775), .Q(n2792) );
  nnd2s1 U3089 ( .DIN1(n2794), .DIN2(n2795), .Q(\IDinst/n5506 ) );
  nnd2s1 U3090 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][12] ), .Q(n2795) );
  nnd2s1 U3091 ( .DIN1(n617), .DIN2(n721), .Q(n2794) );
  nnd2s1 U3092 ( .DIN1(n2796), .DIN2(n2797), .Q(\IDinst/n5505 ) );
  nnd2s1 U3093 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][12] ), .Q(n2797) );
  nnd2s1 U3094 ( .DIN1(n619), .DIN2(n2775), .Q(n2796) );
  nnd2s1 U3095 ( .DIN1(n2798), .DIN2(n2799), .Q(\IDinst/n5504 ) );
  nnd2s1 U3096 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][12] ), .Q(n2799) );
  nnd2s1 U3097 ( .DIN1(n605), .DIN2(n721), .Q(n2798) );
  nnd2s1 U3098 ( .DIN1(n2800), .DIN2(n2801), .Q(\IDinst/n5503 ) );
  nnd2s1 U3099 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][12] ), .Q(n2801) );
  nnd2s1 U3100 ( .DIN1(n607), .DIN2(n2775), .Q(n2800) );
  nnd2s1 U3101 ( .DIN1(n2802), .DIN2(n2803), .Q(\IDinst/n5502 ) );
  nnd2s1 U3102 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][12] ), .Q(n2803) );
  nnd2s1 U3103 ( .DIN1(n609), .DIN2(n721), .Q(n2802) );
  nnd2s1 U3104 ( .DIN1(n2804), .DIN2(n2805), .Q(\IDinst/n5501 ) );
  nnd2s1 U3105 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][12] ), .Q(n2805) );
  nnd2s1 U3106 ( .DIN1(n611), .DIN2(n2775), .Q(n2804) );
  nnd2s1 U3107 ( .DIN1(n2806), .DIN2(n2807), .Q(\IDinst/n5500 ) );
  nnd2s1 U3108 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][12] ), .Q(n2807) );
  nnd2s1 U3109 ( .DIN1(n581), .DIN2(n721), .Q(n2806) );
  nnd2s1 U3110 ( .DIN1(n2808), .DIN2(n2809), .Q(\IDinst/n5499 ) );
  nnd2s1 U3111 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][12] ), .Q(n2809) );
  nnd2s1 U3112 ( .DIN1(n583), .DIN2(n2775), .Q(n2808) );
  nnd2s1 U3113 ( .DIN1(n2810), .DIN2(n2811), .Q(\IDinst/n5498 ) );
  nnd2s1 U3114 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][12] ), .Q(n2811) );
  nnd2s1 U3115 ( .DIN1(n585), .DIN2(n721), .Q(n2810) );
  nnd2s1 U3116 ( .DIN1(n2812), .DIN2(n2813), .Q(\IDinst/n5497 ) );
  nnd2s1 U3117 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][12] ), .Q(n2813) );
  nnd2s1 U3118 ( .DIN1(n587), .DIN2(n2775), .Q(n2812) );
  nnd2s1 U3119 ( .DIN1(n2814), .DIN2(n2815), .Q(\IDinst/n5496 ) );
  nnd2s1 U3120 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][12] ), .Q(n2815) );
  nnd2s1 U3121 ( .DIN1(n573), .DIN2(n721), .Q(n2814) );
  nnd2s1 U3122 ( .DIN1(n2816), .DIN2(n2817), .Q(\IDinst/n5495 ) );
  nnd2s1 U3123 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][12] ), .Q(n2817) );
  nnd2s1 U3124 ( .DIN1(n575), .DIN2(n2775), .Q(n2816) );
  nnd2s1 U3125 ( .DIN1(n2818), .DIN2(n2819), .Q(\IDinst/n5494 ) );
  nnd2s1 U3126 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][12] ), .Q(n2819) );
  nnd2s1 U3127 ( .DIN1(n577), .DIN2(n721), .Q(n2818) );
  nnd2s1 U3128 ( .DIN1(n2820), .DIN2(n2821), .Q(\IDinst/n5493 ) );
  nnd2s1 U3129 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][12] ), .Q(n2821) );
  nnd2s1 U3130 ( .DIN1(n579), .DIN2(n2775), .Q(n2820) );
  nnd2s1 U3131 ( .DIN1(n2822), .DIN2(n2823), .Q(\IDinst/n5492 ) );
  nnd2s1 U3132 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][12] ), .Q(n2823) );
  nnd2s1 U3133 ( .DIN1(n565), .DIN2(n721), .Q(n2822) );
  nnd2s1 U3134 ( .DIN1(n2824), .DIN2(n2825), .Q(\IDinst/n5491 ) );
  nnd2s1 U3135 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][12] ), .Q(n2825) );
  nnd2s1 U3136 ( .DIN1(n567), .DIN2(n2775), .Q(n2824) );
  nnd2s1 U3137 ( .DIN1(n2826), .DIN2(n2827), .Q(\IDinst/n5490 ) );
  nnd2s1 U3138 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][12] ), .Q(n2827) );
  nnd2s1 U3139 ( .DIN1(n569), .DIN2(n721), .Q(n2826) );
  nnd2s1 U3140 ( .DIN1(n2828), .DIN2(n2829), .Q(\IDinst/n5489 ) );
  nnd2s1 U3141 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][12] ), .Q(n2829) );
  nnd2s1 U3142 ( .DIN1(n571), .DIN2(n2775), .Q(n2828) );
  nnd2s1 U3143 ( .DIN1(n2830), .DIN2(n2831), .Q(\IDinst/n5488 ) );
  nnd2s1 U3144 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][12] ), .Q(n2831) );
  nnd2s1 U3145 ( .DIN1(n557), .DIN2(n721), .Q(n2830) );
  nnd2s1 U3146 ( .DIN1(n2832), .DIN2(n2833), .Q(\IDinst/n5487 ) );
  nnd2s1 U3147 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][12] ), .Q(n2833) );
  nnd2s1 U3148 ( .DIN1(n559), .DIN2(n2775), .Q(n2832) );
  nnd2s1 U3149 ( .DIN1(n2834), .DIN2(n2835), .Q(\IDinst/n5486 ) );
  nnd2s1 U3150 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][12] ), .Q(n2835) );
  nnd2s1 U3151 ( .DIN1(n561), .DIN2(n721), .Q(n2834) );
  nnd2s1 U3152 ( .DIN1(n2836), .DIN2(n2837), .Q(\IDinst/n5485 ) );
  nnd2s1 U3153 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][12] ), .Q(n2837) );
  nnd2s1 U3154 ( .DIN1(n563), .DIN2(n2775), .Q(n2836) );
  nnd2s1 U3155 ( .DIN1(n2572), .DIN2(n2838), .Q(n2775) );
  nnd2s1 U3156 ( .DIN1(n2574), .DIN2(n192), .Q(n2838) );
  nnd2s1 U3157 ( .DIN1(n2839), .DIN2(n2840), .Q(\IDinst/n5484 ) );
  nnd2s1 U3158 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][13] ), .Q(n2840) );
  nnd2s1 U3159 ( .DIN1(n596), .DIN2(n737), .Q(n2839) );
  nnd2s1 U3160 ( .DIN1(n2842), .DIN2(n2843), .Q(\IDinst/n5483 ) );
  nnd2s1 U3161 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][13] ), .Q(n2843) );
  nnd2s1 U3162 ( .DIN1(n598), .DIN2(n2841), .Q(n2842) );
  nnd2s1 U3163 ( .DIN1(n2844), .DIN2(n2845), .Q(\IDinst/n5482 ) );
  nnd2s1 U3164 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][13] ), .Q(n2845) );
  nnd2s1 U3165 ( .DIN1(n600), .DIN2(n737), .Q(n2844) );
  nnd2s1 U3166 ( .DIN1(n2846), .DIN2(n2847), .Q(\IDinst/n5481 ) );
  nnd2s1 U3167 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][13] ), .Q(n2847) );
  nnd2s1 U3168 ( .DIN1(n602), .DIN2(n2841), .Q(n2846) );
  nnd2s1 U3169 ( .DIN1(n2848), .DIN2(n2849), .Q(\IDinst/n5480 ) );
  nnd2s1 U3170 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][13] ), .Q(n2849) );
  nnd2s1 U3171 ( .DIN1(n588), .DIN2(n737), .Q(n2848) );
  nnd2s1 U3172 ( .DIN1(n2850), .DIN2(n2851), .Q(\IDinst/n5479 ) );
  nnd2s1 U3173 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][13] ), .Q(n2851) );
  nnd2s1 U3174 ( .DIN1(n590), .DIN2(n2841), .Q(n2850) );
  nnd2s1 U3175 ( .DIN1(n2852), .DIN2(n2853), .Q(\IDinst/n5478 ) );
  nnd2s1 U3176 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][13] ), .Q(n2853) );
  nnd2s1 U3177 ( .DIN1(n592), .DIN2(n737), .Q(n2852) );
  nnd2s1 U3178 ( .DIN1(n2854), .DIN2(n2855), .Q(\IDinst/n5477 ) );
  nnd2s1 U3179 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][13] ), .Q(n2855) );
  nnd2s1 U3180 ( .DIN1(n594), .DIN2(n2841), .Q(n2854) );
  nnd2s1 U3181 ( .DIN1(n2856), .DIN2(n2857), .Q(\IDinst/n5476 ) );
  nnd2s1 U3182 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][13] ), .Q(n2857) );
  nnd2s1 U3183 ( .DIN1(n612), .DIN2(n737), .Q(n2856) );
  nnd2s1 U3184 ( .DIN1(n2858), .DIN2(n2859), .Q(\IDinst/n5475 ) );
  nnd2s1 U3185 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][13] ), .Q(n2859) );
  nnd2s1 U3186 ( .DIN1(n614), .DIN2(n2841), .Q(n2858) );
  nnd2s1 U3187 ( .DIN1(n2860), .DIN2(n2861), .Q(\IDinst/n5474 ) );
  nnd2s1 U3188 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][13] ), .Q(n2861) );
  nnd2s1 U3189 ( .DIN1(n616), .DIN2(n737), .Q(n2860) );
  nnd2s1 U3190 ( .DIN1(n2862), .DIN2(n2863), .Q(\IDinst/n5473 ) );
  nnd2s1 U3191 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][13] ), .Q(n2863) );
  nnd2s1 U3192 ( .DIN1(n618), .DIN2(n2841), .Q(n2862) );
  nnd2s1 U3193 ( .DIN1(n2864), .DIN2(n2865), .Q(\IDinst/n5472 ) );
  nnd2s1 U3194 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][13] ), .Q(n2865) );
  nnd2s1 U3195 ( .DIN1(n604), .DIN2(n737), .Q(n2864) );
  nnd2s1 U3196 ( .DIN1(n2866), .DIN2(n2867), .Q(\IDinst/n5471 ) );
  nnd2s1 U3197 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][13] ), .Q(n2867) );
  nnd2s1 U3198 ( .DIN1(n606), .DIN2(n2841), .Q(n2866) );
  nnd2s1 U3199 ( .DIN1(n2868), .DIN2(n2869), .Q(\IDinst/n5470 ) );
  nnd2s1 U3200 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][13] ), .Q(n2869) );
  nnd2s1 U3201 ( .DIN1(n608), .DIN2(n737), .Q(n2868) );
  nnd2s1 U3202 ( .DIN1(n2870), .DIN2(n2871), .Q(\IDinst/n5469 ) );
  nnd2s1 U3203 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][13] ), .Q(n2871) );
  nnd2s1 U3204 ( .DIN1(n610), .DIN2(n2841), .Q(n2870) );
  nnd2s1 U3205 ( .DIN1(n2872), .DIN2(n2873), .Q(\IDinst/n5468 ) );
  nnd2s1 U3206 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][13] ), .Q(n2873) );
  nnd2s1 U3207 ( .DIN1(n580), .DIN2(n737), .Q(n2872) );
  nnd2s1 U3208 ( .DIN1(n2874), .DIN2(n2875), .Q(\IDinst/n5467 ) );
  nnd2s1 U3209 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][13] ), .Q(n2875) );
  nnd2s1 U3210 ( .DIN1(n582), .DIN2(n2841), .Q(n2874) );
  nnd2s1 U3211 ( .DIN1(n2876), .DIN2(n2877), .Q(\IDinst/n5466 ) );
  nnd2s1 U3212 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][13] ), .Q(n2877) );
  nnd2s1 U3213 ( .DIN1(n584), .DIN2(n737), .Q(n2876) );
  nnd2s1 U3214 ( .DIN1(n2878), .DIN2(n2879), .Q(\IDinst/n5465 ) );
  nnd2s1 U3215 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][13] ), .Q(n2879) );
  nnd2s1 U3216 ( .DIN1(n586), .DIN2(n2841), .Q(n2878) );
  nnd2s1 U3217 ( .DIN1(n2880), .DIN2(n2881), .Q(\IDinst/n5464 ) );
  nnd2s1 U3218 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][13] ), .Q(n2881) );
  nnd2s1 U3219 ( .DIN1(n572), .DIN2(n737), .Q(n2880) );
  nnd2s1 U3220 ( .DIN1(n2882), .DIN2(n2883), .Q(\IDinst/n5463 ) );
  nnd2s1 U3221 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][13] ), .Q(n2883) );
  nnd2s1 U3222 ( .DIN1(n574), .DIN2(n2841), .Q(n2882) );
  nnd2s1 U3223 ( .DIN1(n2884), .DIN2(n2885), .Q(\IDinst/n5462 ) );
  nnd2s1 U3224 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][13] ), .Q(n2885) );
  nnd2s1 U3225 ( .DIN1(n576), .DIN2(n737), .Q(n2884) );
  nnd2s1 U3226 ( .DIN1(n2886), .DIN2(n2887), .Q(\IDinst/n5461 ) );
  nnd2s1 U3227 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][13] ), .Q(n2887) );
  nnd2s1 U3228 ( .DIN1(n578), .DIN2(n2841), .Q(n2886) );
  nnd2s1 U3229 ( .DIN1(n2888), .DIN2(n2889), .Q(\IDinst/n5460 ) );
  nnd2s1 U3230 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][13] ), .Q(n2889) );
  nnd2s1 U3231 ( .DIN1(n564), .DIN2(n737), .Q(n2888) );
  nnd2s1 U3232 ( .DIN1(n2890), .DIN2(n2891), .Q(\IDinst/n5459 ) );
  nnd2s1 U3233 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][13] ), .Q(n2891) );
  nnd2s1 U3234 ( .DIN1(n566), .DIN2(n2841), .Q(n2890) );
  nnd2s1 U3235 ( .DIN1(n2892), .DIN2(n2893), .Q(\IDinst/n5458 ) );
  nnd2s1 U3236 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][13] ), .Q(n2893) );
  nnd2s1 U3237 ( .DIN1(n568), .DIN2(n737), .Q(n2892) );
  nnd2s1 U3238 ( .DIN1(n2894), .DIN2(n2895), .Q(\IDinst/n5457 ) );
  nnd2s1 U3239 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][13] ), .Q(n2895) );
  nnd2s1 U3240 ( .DIN1(n570), .DIN2(n2841), .Q(n2894) );
  nnd2s1 U3241 ( .DIN1(n2896), .DIN2(n2897), .Q(\IDinst/n5456 ) );
  nnd2s1 U3242 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][13] ), .Q(n2897) );
  nnd2s1 U3243 ( .DIN1(n556), .DIN2(n737), .Q(n2896) );
  nnd2s1 U3244 ( .DIN1(n2898), .DIN2(n2899), .Q(\IDinst/n5455 ) );
  nnd2s1 U3245 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][13] ), .Q(n2899) );
  nnd2s1 U3246 ( .DIN1(n558), .DIN2(n2841), .Q(n2898) );
  nnd2s1 U3247 ( .DIN1(n2900), .DIN2(n2901), .Q(\IDinst/n5454 ) );
  nnd2s1 U3248 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][13] ), .Q(n2901) );
  nnd2s1 U3249 ( .DIN1(n560), .DIN2(n737), .Q(n2900) );
  nnd2s1 U3250 ( .DIN1(n2902), .DIN2(n2903), .Q(\IDinst/n5453 ) );
  nnd2s1 U3251 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][13] ), .Q(n2903) );
  nnd2s1 U3252 ( .DIN1(n562), .DIN2(n2841), .Q(n2902) );
  nnd2s1 U3253 ( .DIN1(n2572), .DIN2(n2904), .Q(n2841) );
  nnd2s1 U3254 ( .DIN1(n2574), .DIN2(n190), .Q(n2904) );
  nnd2s1 U3255 ( .DIN1(n2905), .DIN2(n2906), .Q(\IDinst/n5452 ) );
  nnd2s1 U3256 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][14] ), .Q(n2906) );
  nnd2s1 U3257 ( .DIN1(n597), .DIN2(n765), .Q(n2905) );
  nnd2s1 U3258 ( .DIN1(n2908), .DIN2(n2909), .Q(\IDinst/n5451 ) );
  nnd2s1 U3259 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][14] ), .Q(n2909) );
  nnd2s1 U3260 ( .DIN1(n599), .DIN2(n2907), .Q(n2908) );
  nnd2s1 U3261 ( .DIN1(n2910), .DIN2(n2911), .Q(\IDinst/n5450 ) );
  nnd2s1 U3262 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][14] ), .Q(n2911) );
  nnd2s1 U3263 ( .DIN1(n601), .DIN2(n765), .Q(n2910) );
  nnd2s1 U3264 ( .DIN1(n2912), .DIN2(n2913), .Q(\IDinst/n5449 ) );
  nnd2s1 U3265 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][14] ), .Q(n2913) );
  nnd2s1 U3266 ( .DIN1(n603), .DIN2(n2907), .Q(n2912) );
  nnd2s1 U3267 ( .DIN1(n2914), .DIN2(n2915), .Q(\IDinst/n5448 ) );
  nnd2s1 U3268 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][14] ), .Q(n2915) );
  nnd2s1 U3269 ( .DIN1(n589), .DIN2(n765), .Q(n2914) );
  nnd2s1 U3270 ( .DIN1(n2916), .DIN2(n2917), .Q(\IDinst/n5447 ) );
  nnd2s1 U3271 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][14] ), .Q(n2917) );
  nnd2s1 U3272 ( .DIN1(n591), .DIN2(n2907), .Q(n2916) );
  nnd2s1 U3273 ( .DIN1(n2918), .DIN2(n2919), .Q(\IDinst/n5446 ) );
  nnd2s1 U3274 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][14] ), .Q(n2919) );
  nnd2s1 U3275 ( .DIN1(n593), .DIN2(n765), .Q(n2918) );
  nnd2s1 U3276 ( .DIN1(n2920), .DIN2(n2921), .Q(\IDinst/n5445 ) );
  nnd2s1 U3277 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][14] ), .Q(n2921) );
  nnd2s1 U3278 ( .DIN1(n595), .DIN2(n2907), .Q(n2920) );
  nnd2s1 U3279 ( .DIN1(n2922), .DIN2(n2923), .Q(\IDinst/n5444 ) );
  nnd2s1 U3280 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][14] ), .Q(n2923) );
  nnd2s1 U3281 ( .DIN1(n613), .DIN2(n765), .Q(n2922) );
  nnd2s1 U3282 ( .DIN1(n2924), .DIN2(n2925), .Q(\IDinst/n5443 ) );
  nnd2s1 U3283 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][14] ), .Q(n2925) );
  nnd2s1 U3284 ( .DIN1(n615), .DIN2(n2907), .Q(n2924) );
  nnd2s1 U3285 ( .DIN1(n2926), .DIN2(n2927), .Q(\IDinst/n5442 ) );
  nnd2s1 U3286 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][14] ), .Q(n2927) );
  nnd2s1 U3287 ( .DIN1(n617), .DIN2(n765), .Q(n2926) );
  nnd2s1 U3288 ( .DIN1(n2928), .DIN2(n2929), .Q(\IDinst/n5441 ) );
  nnd2s1 U3289 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][14] ), .Q(n2929) );
  nnd2s1 U3290 ( .DIN1(n619), .DIN2(n2907), .Q(n2928) );
  nnd2s1 U3291 ( .DIN1(n2930), .DIN2(n2931), .Q(\IDinst/n5440 ) );
  nnd2s1 U3292 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][14] ), .Q(n2931) );
  nnd2s1 U3293 ( .DIN1(n605), .DIN2(n765), .Q(n2930) );
  nnd2s1 U3294 ( .DIN1(n2932), .DIN2(n2933), .Q(\IDinst/n5439 ) );
  nnd2s1 U3295 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][14] ), .Q(n2933) );
  nnd2s1 U3296 ( .DIN1(n607), .DIN2(n2907), .Q(n2932) );
  nnd2s1 U3297 ( .DIN1(n2934), .DIN2(n2935), .Q(\IDinst/n5438 ) );
  nnd2s1 U3298 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][14] ), .Q(n2935) );
  nnd2s1 U3299 ( .DIN1(n609), .DIN2(n765), .Q(n2934) );
  nnd2s1 U3300 ( .DIN1(n2936), .DIN2(n2937), .Q(\IDinst/n5437 ) );
  nnd2s1 U3301 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][14] ), .Q(n2937) );
  nnd2s1 U3302 ( .DIN1(n611), .DIN2(n2907), .Q(n2936) );
  nnd2s1 U3303 ( .DIN1(n2938), .DIN2(n2939), .Q(\IDinst/n5436 ) );
  nnd2s1 U3304 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][14] ), .Q(n2939) );
  nnd2s1 U3305 ( .DIN1(n581), .DIN2(n765), .Q(n2938) );
  nnd2s1 U3306 ( .DIN1(n2940), .DIN2(n2941), .Q(\IDinst/n5435 ) );
  nnd2s1 U3307 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][14] ), .Q(n2941) );
  nnd2s1 U3308 ( .DIN1(n583), .DIN2(n2907), .Q(n2940) );
  nnd2s1 U3309 ( .DIN1(n2942), .DIN2(n2943), .Q(\IDinst/n5434 ) );
  nnd2s1 U3310 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][14] ), .Q(n2943) );
  nnd2s1 U3311 ( .DIN1(n585), .DIN2(n765), .Q(n2942) );
  nnd2s1 U3312 ( .DIN1(n2944), .DIN2(n2945), .Q(\IDinst/n5433 ) );
  nnd2s1 U3313 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][14] ), .Q(n2945) );
  nnd2s1 U3314 ( .DIN1(n587), .DIN2(n2907), .Q(n2944) );
  nnd2s1 U3315 ( .DIN1(n2946), .DIN2(n2947), .Q(\IDinst/n5432 ) );
  nnd2s1 U3316 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][14] ), .Q(n2947) );
  nnd2s1 U3317 ( .DIN1(n573), .DIN2(n765), .Q(n2946) );
  nnd2s1 U3318 ( .DIN1(n2948), .DIN2(n2949), .Q(\IDinst/n5431 ) );
  nnd2s1 U3319 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][14] ), .Q(n2949) );
  nnd2s1 U3320 ( .DIN1(n575), .DIN2(n2907), .Q(n2948) );
  nnd2s1 U3321 ( .DIN1(n2950), .DIN2(n2951), .Q(\IDinst/n5430 ) );
  nnd2s1 U3322 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][14] ), .Q(n2951) );
  nnd2s1 U3323 ( .DIN1(n577), .DIN2(n765), .Q(n2950) );
  nnd2s1 U3324 ( .DIN1(n2952), .DIN2(n2953), .Q(\IDinst/n5429 ) );
  nnd2s1 U3325 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][14] ), .Q(n2953) );
  nnd2s1 U3326 ( .DIN1(n579), .DIN2(n2907), .Q(n2952) );
  nnd2s1 U3327 ( .DIN1(n2954), .DIN2(n2955), .Q(\IDinst/n5428 ) );
  nnd2s1 U3328 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][14] ), .Q(n2955) );
  nnd2s1 U3329 ( .DIN1(n565), .DIN2(n765), .Q(n2954) );
  nnd2s1 U3330 ( .DIN1(n2956), .DIN2(n2957), .Q(\IDinst/n5427 ) );
  nnd2s1 U3331 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][14] ), .Q(n2957) );
  nnd2s1 U3332 ( .DIN1(n567), .DIN2(n2907), .Q(n2956) );
  nnd2s1 U3333 ( .DIN1(n2958), .DIN2(n2959), .Q(\IDinst/n5426 ) );
  nnd2s1 U3334 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][14] ), .Q(n2959) );
  nnd2s1 U3335 ( .DIN1(n569), .DIN2(n765), .Q(n2958) );
  nnd2s1 U3336 ( .DIN1(n2960), .DIN2(n2961), .Q(\IDinst/n5425 ) );
  nnd2s1 U3337 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][14] ), .Q(n2961) );
  nnd2s1 U3338 ( .DIN1(n571), .DIN2(n2907), .Q(n2960) );
  nnd2s1 U3339 ( .DIN1(n2962), .DIN2(n2963), .Q(\IDinst/n5424 ) );
  nnd2s1 U3340 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][14] ), .Q(n2963) );
  nnd2s1 U3341 ( .DIN1(n557), .DIN2(n765), .Q(n2962) );
  nnd2s1 U3342 ( .DIN1(n2964), .DIN2(n2965), .Q(\IDinst/n5423 ) );
  nnd2s1 U3343 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][14] ), .Q(n2965) );
  nnd2s1 U3344 ( .DIN1(n559), .DIN2(n2907), .Q(n2964) );
  nnd2s1 U3345 ( .DIN1(n2966), .DIN2(n2967), .Q(\IDinst/n5422 ) );
  nnd2s1 U3346 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][14] ), .Q(n2967) );
  nnd2s1 U3347 ( .DIN1(n561), .DIN2(n765), .Q(n2966) );
  nnd2s1 U3348 ( .DIN1(n2968), .DIN2(n2969), .Q(\IDinst/n5421 ) );
  nnd2s1 U3349 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][14] ), .Q(n2969) );
  nnd2s1 U3350 ( .DIN1(n563), .DIN2(n2907), .Q(n2968) );
  nnd2s1 U3351 ( .DIN1(n2572), .DIN2(n2970), .Q(n2907) );
  nnd2s1 U3352 ( .DIN1(n2574), .DIN2(n188), .Q(n2970) );
  or3s1 U3353 ( .DIN1(\IDinst/opcode_of_WB[2] ), .DIN2(n9404), .DIN3(n2574), 
        .Q(n2572) );
  nnd2s1 U3354 ( .DIN1(n2971), .DIN2(n2972), .Q(\IDinst/n5420 ) );
  nnd2s1 U3355 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][15] ), .Q(n2972) );
  nnd2s1 U3356 ( .DIN1(n596), .DIN2(n445), .Q(n2971) );
  nnd2s1 U3357 ( .DIN1(n2973), .DIN2(n2974), .Q(\IDinst/n5419 ) );
  nnd2s1 U3358 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][15] ), .Q(n2974) );
  nnd2s1 U3359 ( .DIN1(n598), .DIN2(n444), .Q(n2973) );
  nnd2s1 U3360 ( .DIN1(n2975), .DIN2(n2976), .Q(\IDinst/n5418 ) );
  nnd2s1 U3361 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][15] ), .Q(n2976) );
  nnd2s1 U3362 ( .DIN1(n600), .DIN2(n445), .Q(n2975) );
  nnd2s1 U3363 ( .DIN1(n2977), .DIN2(n2978), .Q(\IDinst/n5417 ) );
  nnd2s1 U3364 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][15] ), .Q(n2978) );
  nnd2s1 U3365 ( .DIN1(n602), .DIN2(n444), .Q(n2977) );
  nnd2s1 U3366 ( .DIN1(n2979), .DIN2(n2980), .Q(\IDinst/n5416 ) );
  nnd2s1 U3367 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][15] ), .Q(n2980) );
  nnd2s1 U3368 ( .DIN1(n588), .DIN2(n445), .Q(n2979) );
  nnd2s1 U3369 ( .DIN1(n2981), .DIN2(n2982), .Q(\IDinst/n5415 ) );
  nnd2s1 U3370 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][15] ), .Q(n2982) );
  nnd2s1 U3371 ( .DIN1(n590), .DIN2(n444), .Q(n2981) );
  nnd2s1 U3372 ( .DIN1(n2983), .DIN2(n2984), .Q(\IDinst/n5414 ) );
  nnd2s1 U3373 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][15] ), .Q(n2984) );
  nnd2s1 U3374 ( .DIN1(n592), .DIN2(n445), .Q(n2983) );
  nnd2s1 U3375 ( .DIN1(n2985), .DIN2(n2986), .Q(\IDinst/n5413 ) );
  nnd2s1 U3376 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][15] ), .Q(n2986) );
  nnd2s1 U3377 ( .DIN1(n594), .DIN2(n444), .Q(n2985) );
  nnd2s1 U3378 ( .DIN1(n2987), .DIN2(n2988), .Q(\IDinst/n5412 ) );
  nnd2s1 U3379 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][15] ), .Q(n2988) );
  nnd2s1 U3380 ( .DIN1(n612), .DIN2(n445), .Q(n2987) );
  nnd2s1 U3381 ( .DIN1(n2989), .DIN2(n2990), .Q(\IDinst/n5411 ) );
  nnd2s1 U3382 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][15] ), .Q(n2990) );
  nnd2s1 U3383 ( .DIN1(n614), .DIN2(n444), .Q(n2989) );
  nnd2s1 U3384 ( .DIN1(n2991), .DIN2(n2992), .Q(\IDinst/n5410 ) );
  nnd2s1 U3385 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][15] ), .Q(n2992) );
  nnd2s1 U3386 ( .DIN1(n616), .DIN2(n445), .Q(n2991) );
  nnd2s1 U3387 ( .DIN1(n2993), .DIN2(n2994), .Q(\IDinst/n5409 ) );
  nnd2s1 U3388 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][15] ), .Q(n2994) );
  nnd2s1 U3389 ( .DIN1(n618), .DIN2(n444), .Q(n2993) );
  nnd2s1 U3390 ( .DIN1(n2995), .DIN2(n2996), .Q(\IDinst/n5408 ) );
  nnd2s1 U3391 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][15] ), .Q(n2996) );
  nnd2s1 U3392 ( .DIN1(n604), .DIN2(n445), .Q(n2995) );
  nnd2s1 U3393 ( .DIN1(n2997), .DIN2(n2998), .Q(\IDinst/n5407 ) );
  nnd2s1 U3394 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][15] ), .Q(n2998) );
  nnd2s1 U3395 ( .DIN1(n606), .DIN2(n444), .Q(n2997) );
  nnd2s1 U3396 ( .DIN1(n2999), .DIN2(n3000), .Q(\IDinst/n5406 ) );
  nnd2s1 U3397 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][15] ), .Q(n3000) );
  nnd2s1 U3398 ( .DIN1(n608), .DIN2(n445), .Q(n2999) );
  nnd2s1 U3399 ( .DIN1(n3001), .DIN2(n3002), .Q(\IDinst/n5405 ) );
  nnd2s1 U3400 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][15] ), .Q(n3002) );
  nnd2s1 U3401 ( .DIN1(n610), .DIN2(n444), .Q(n3001) );
  nnd2s1 U3402 ( .DIN1(n3003), .DIN2(n3004), .Q(\IDinst/n5404 ) );
  nnd2s1 U3403 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][15] ), .Q(n3004) );
  nnd2s1 U3404 ( .DIN1(n580), .DIN2(n445), .Q(n3003) );
  nnd2s1 U3405 ( .DIN1(n3005), .DIN2(n3006), .Q(\IDinst/n5403 ) );
  nnd2s1 U3406 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][15] ), .Q(n3006) );
  nnd2s1 U3407 ( .DIN1(n582), .DIN2(n444), .Q(n3005) );
  nnd2s1 U3408 ( .DIN1(n3007), .DIN2(n3008), .Q(\IDinst/n5402 ) );
  nnd2s1 U3409 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][15] ), .Q(n3008) );
  nnd2s1 U3410 ( .DIN1(n584), .DIN2(n445), .Q(n3007) );
  nnd2s1 U3411 ( .DIN1(n3009), .DIN2(n3010), .Q(\IDinst/n5401 ) );
  nnd2s1 U3412 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][15] ), .Q(n3010) );
  nnd2s1 U3413 ( .DIN1(n586), .DIN2(n444), .Q(n3009) );
  nnd2s1 U3414 ( .DIN1(n3011), .DIN2(n3012), .Q(\IDinst/n5400 ) );
  nnd2s1 U3415 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][15] ), .Q(n3012) );
  nnd2s1 U3416 ( .DIN1(n572), .DIN2(n445), .Q(n3011) );
  nnd2s1 U3417 ( .DIN1(n3013), .DIN2(n3014), .Q(\IDinst/n5399 ) );
  nnd2s1 U3418 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][15] ), .Q(n3014) );
  nnd2s1 U3419 ( .DIN1(n574), .DIN2(n444), .Q(n3013) );
  nnd2s1 U3420 ( .DIN1(n3015), .DIN2(n3016), .Q(\IDinst/n5398 ) );
  nnd2s1 U3421 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][15] ), .Q(n3016) );
  nnd2s1 U3422 ( .DIN1(n576), .DIN2(n445), .Q(n3015) );
  nnd2s1 U3423 ( .DIN1(n3017), .DIN2(n3018), .Q(\IDinst/n5397 ) );
  nnd2s1 U3424 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][15] ), .Q(n3018) );
  nnd2s1 U3425 ( .DIN1(n578), .DIN2(n444), .Q(n3017) );
  nnd2s1 U3426 ( .DIN1(n3019), .DIN2(n3020), .Q(\IDinst/n5396 ) );
  nnd2s1 U3427 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][15] ), .Q(n3020) );
  nnd2s1 U3428 ( .DIN1(n564), .DIN2(n445), .Q(n3019) );
  nnd2s1 U3429 ( .DIN1(n3021), .DIN2(n3022), .Q(\IDinst/n5395 ) );
  nnd2s1 U3430 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][15] ), .Q(n3022) );
  nnd2s1 U3431 ( .DIN1(n566), .DIN2(n444), .Q(n3021) );
  nnd2s1 U3432 ( .DIN1(n3023), .DIN2(n3024), .Q(\IDinst/n5394 ) );
  nnd2s1 U3433 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][15] ), .Q(n3024) );
  nnd2s1 U3434 ( .DIN1(n568), .DIN2(n445), .Q(n3023) );
  nnd2s1 U3435 ( .DIN1(n3025), .DIN2(n3026), .Q(\IDinst/n5393 ) );
  nnd2s1 U3436 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][15] ), .Q(n3026) );
  nnd2s1 U3437 ( .DIN1(n570), .DIN2(n444), .Q(n3025) );
  nnd2s1 U3438 ( .DIN1(n3027), .DIN2(n3028), .Q(\IDinst/n5392 ) );
  nnd2s1 U3439 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][15] ), .Q(n3028) );
  nnd2s1 U3440 ( .DIN1(n556), .DIN2(n445), .Q(n3027) );
  nnd2s1 U3441 ( .DIN1(n3029), .DIN2(n3030), .Q(\IDinst/n5391 ) );
  nnd2s1 U3442 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][15] ), .Q(n3030) );
  nnd2s1 U3443 ( .DIN1(n558), .DIN2(n444), .Q(n3029) );
  nnd2s1 U3444 ( .DIN1(n3031), .DIN2(n3032), .Q(\IDinst/n5390 ) );
  nnd2s1 U3445 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][15] ), .Q(n3032) );
  nnd2s1 U3446 ( .DIN1(n560), .DIN2(n445), .Q(n3031) );
  nnd2s1 U3447 ( .DIN1(n3033), .DIN2(n3034), .Q(\IDinst/n5389 ) );
  nnd2s1 U3448 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][15] ), .Q(n3034) );
  nnd2s1 U3449 ( .DIN1(n562), .DIN2(n444), .Q(n3033) );
  nnd2s1 U3450 ( .DIN1(n2574), .DIN2(n129), .Q(n3036) );
  nnd2s1 U3451 ( .DIN1(n9405), .DIN2(n3037), .Q(n2574) );
  nnd2s1 U3452 ( .DIN1(n3038), .DIN2(n3039), .Q(\IDinst/n5388 ) );
  nnd2s1 U3453 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][16] ), .Q(n3039) );
  nnd2s1 U3454 ( .DIN1(n597), .DIN2(n447), .Q(n3038) );
  nnd2s1 U3455 ( .DIN1(n3040), .DIN2(n3041), .Q(\IDinst/n5387 ) );
  nnd2s1 U3456 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][16] ), .Q(n3041) );
  nnd2s1 U3457 ( .DIN1(n599), .DIN2(n446), .Q(n3040) );
  nnd2s1 U3458 ( .DIN1(n3042), .DIN2(n3043), .Q(\IDinst/n5386 ) );
  nnd2s1 U3459 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][16] ), .Q(n3043) );
  nnd2s1 U3460 ( .DIN1(n601), .DIN2(n447), .Q(n3042) );
  nnd2s1 U3461 ( .DIN1(n3044), .DIN2(n3045), .Q(\IDinst/n5385 ) );
  nnd2s1 U3462 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][16] ), .Q(n3045) );
  nnd2s1 U3463 ( .DIN1(n603), .DIN2(n446), .Q(n3044) );
  nnd2s1 U3464 ( .DIN1(n3046), .DIN2(n3047), .Q(\IDinst/n5384 ) );
  nnd2s1 U3465 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][16] ), .Q(n3047) );
  nnd2s1 U3466 ( .DIN1(n589), .DIN2(n447), .Q(n3046) );
  nnd2s1 U3467 ( .DIN1(n3048), .DIN2(n3049), .Q(\IDinst/n5383 ) );
  nnd2s1 U3468 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][16] ), .Q(n3049) );
  nnd2s1 U3469 ( .DIN1(n591), .DIN2(n446), .Q(n3048) );
  nnd2s1 U3470 ( .DIN1(n3050), .DIN2(n3051), .Q(\IDinst/n5382 ) );
  nnd2s1 U3471 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][16] ), .Q(n3051) );
  nnd2s1 U3472 ( .DIN1(n593), .DIN2(n447), .Q(n3050) );
  nnd2s1 U3473 ( .DIN1(n3052), .DIN2(n3053), .Q(\IDinst/n5381 ) );
  nnd2s1 U3474 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][16] ), .Q(n3053) );
  nnd2s1 U3475 ( .DIN1(n595), .DIN2(n446), .Q(n3052) );
  nnd2s1 U3476 ( .DIN1(n3054), .DIN2(n3055), .Q(\IDinst/n5380 ) );
  nnd2s1 U3477 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][16] ), .Q(n3055) );
  nnd2s1 U3478 ( .DIN1(n613), .DIN2(n447), .Q(n3054) );
  nnd2s1 U3479 ( .DIN1(n3056), .DIN2(n3057), .Q(\IDinst/n5379 ) );
  nnd2s1 U3480 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][16] ), .Q(n3057) );
  nnd2s1 U3481 ( .DIN1(n615), .DIN2(n446), .Q(n3056) );
  nnd2s1 U3482 ( .DIN1(n3058), .DIN2(n3059), .Q(\IDinst/n5378 ) );
  nnd2s1 U3483 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][16] ), .Q(n3059) );
  nnd2s1 U3484 ( .DIN1(n617), .DIN2(n447), .Q(n3058) );
  nnd2s1 U3485 ( .DIN1(n3060), .DIN2(n3061), .Q(\IDinst/n5377 ) );
  nnd2s1 U3486 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][16] ), .Q(n3061) );
  nnd2s1 U3487 ( .DIN1(n619), .DIN2(n446), .Q(n3060) );
  nnd2s1 U3488 ( .DIN1(n3062), .DIN2(n3063), .Q(\IDinst/n5376 ) );
  nnd2s1 U3489 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][16] ), .Q(n3063) );
  nnd2s1 U3490 ( .DIN1(n605), .DIN2(n447), .Q(n3062) );
  nnd2s1 U3491 ( .DIN1(n3064), .DIN2(n3065), .Q(\IDinst/n5375 ) );
  nnd2s1 U3492 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][16] ), .Q(n3065) );
  nnd2s1 U3493 ( .DIN1(n607), .DIN2(n446), .Q(n3064) );
  nnd2s1 U3494 ( .DIN1(n3066), .DIN2(n3067), .Q(\IDinst/n5374 ) );
  nnd2s1 U3495 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][16] ), .Q(n3067) );
  nnd2s1 U3496 ( .DIN1(n609), .DIN2(n447), .Q(n3066) );
  nnd2s1 U3497 ( .DIN1(n3068), .DIN2(n3069), .Q(\IDinst/n5373 ) );
  nnd2s1 U3498 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][16] ), .Q(n3069) );
  nnd2s1 U3499 ( .DIN1(n611), .DIN2(n446), .Q(n3068) );
  nnd2s1 U3500 ( .DIN1(n3070), .DIN2(n3071), .Q(\IDinst/n5372 ) );
  nnd2s1 U3501 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][16] ), .Q(n3071) );
  nnd2s1 U3502 ( .DIN1(n581), .DIN2(n447), .Q(n3070) );
  nnd2s1 U3503 ( .DIN1(n3072), .DIN2(n3073), .Q(\IDinst/n5371 ) );
  nnd2s1 U3504 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][16] ), .Q(n3073) );
  nnd2s1 U3505 ( .DIN1(n583), .DIN2(n446), .Q(n3072) );
  nnd2s1 U3506 ( .DIN1(n3074), .DIN2(n3075), .Q(\IDinst/n5370 ) );
  nnd2s1 U3507 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][16] ), .Q(n3075) );
  nnd2s1 U3508 ( .DIN1(n585), .DIN2(n447), .Q(n3074) );
  nnd2s1 U3509 ( .DIN1(n3076), .DIN2(n3077), .Q(\IDinst/n5369 ) );
  nnd2s1 U3510 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][16] ), .Q(n3077) );
  nnd2s1 U3511 ( .DIN1(n587), .DIN2(n446), .Q(n3076) );
  nnd2s1 U3512 ( .DIN1(n3078), .DIN2(n3079), .Q(\IDinst/n5368 ) );
  nnd2s1 U3513 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][16] ), .Q(n3079) );
  nnd2s1 U3514 ( .DIN1(n573), .DIN2(n447), .Q(n3078) );
  nnd2s1 U3515 ( .DIN1(n3080), .DIN2(n3081), .Q(\IDinst/n5367 ) );
  nnd2s1 U3516 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][16] ), .Q(n3081) );
  nnd2s1 U3517 ( .DIN1(n575), .DIN2(n446), .Q(n3080) );
  nnd2s1 U3518 ( .DIN1(n3082), .DIN2(n3083), .Q(\IDinst/n5366 ) );
  nnd2s1 U3519 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][16] ), .Q(n3083) );
  nnd2s1 U3520 ( .DIN1(n577), .DIN2(n447), .Q(n3082) );
  nnd2s1 U3521 ( .DIN1(n3084), .DIN2(n3085), .Q(\IDinst/n5365 ) );
  nnd2s1 U3522 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][16] ), .Q(n3085) );
  nnd2s1 U3523 ( .DIN1(n579), .DIN2(n446), .Q(n3084) );
  nnd2s1 U3524 ( .DIN1(n3086), .DIN2(n3087), .Q(\IDinst/n5364 ) );
  nnd2s1 U3525 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][16] ), .Q(n3087) );
  nnd2s1 U3526 ( .DIN1(n565), .DIN2(n447), .Q(n3086) );
  nnd2s1 U3527 ( .DIN1(n3088), .DIN2(n3089), .Q(\IDinst/n5363 ) );
  nnd2s1 U3528 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][16] ), .Q(n3089) );
  nnd2s1 U3529 ( .DIN1(n567), .DIN2(n446), .Q(n3088) );
  nnd2s1 U3530 ( .DIN1(n3090), .DIN2(n3091), .Q(\IDinst/n5362 ) );
  nnd2s1 U3531 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][16] ), .Q(n3091) );
  nnd2s1 U3532 ( .DIN1(n569), .DIN2(n447), .Q(n3090) );
  nnd2s1 U3533 ( .DIN1(n3092), .DIN2(n3093), .Q(\IDinst/n5361 ) );
  nnd2s1 U3534 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][16] ), .Q(n3093) );
  nnd2s1 U3535 ( .DIN1(n571), .DIN2(n446), .Q(n3092) );
  nnd2s1 U3536 ( .DIN1(n3094), .DIN2(n3095), .Q(\IDinst/n5360 ) );
  nnd2s1 U3537 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][16] ), .Q(n3095) );
  nnd2s1 U3538 ( .DIN1(n557), .DIN2(n447), .Q(n3094) );
  nnd2s1 U3539 ( .DIN1(n3096), .DIN2(n3097), .Q(\IDinst/n5359 ) );
  nnd2s1 U3540 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][16] ), .Q(n3097) );
  nnd2s1 U3541 ( .DIN1(n559), .DIN2(n446), .Q(n3096) );
  nnd2s1 U3542 ( .DIN1(n3098), .DIN2(n3099), .Q(\IDinst/n5358 ) );
  nnd2s1 U3543 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][16] ), .Q(n3099) );
  nnd2s1 U3544 ( .DIN1(n561), .DIN2(n447), .Q(n3098) );
  nnd2s1 U3545 ( .DIN1(n3100), .DIN2(n3101), .Q(\IDinst/n5357 ) );
  nnd2s1 U3546 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][16] ), .Q(n3101) );
  nnd2s1 U3547 ( .DIN1(n563), .DIN2(n446), .Q(n3100) );
  nnd2s1 U3548 ( .DIN1(n3103), .DIN2(n185), .Q(n3102) );
  nnd2s1 U3549 ( .DIN1(n3104), .DIN2(n3105), .Q(\IDinst/n5356 ) );
  nnd2s1 U3550 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][17] ), .Q(n3105) );
  nnd2s1 U3551 ( .DIN1(n596), .DIN2(n449), .Q(n3104) );
  nnd2s1 U3552 ( .DIN1(n3106), .DIN2(n3107), .Q(\IDinst/n5355 ) );
  nnd2s1 U3553 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][17] ), .Q(n3107) );
  nnd2s1 U3554 ( .DIN1(n598), .DIN2(n448), .Q(n3106) );
  nnd2s1 U3555 ( .DIN1(n3108), .DIN2(n3109), .Q(\IDinst/n5354 ) );
  nnd2s1 U3556 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][17] ), .Q(n3109) );
  nnd2s1 U3557 ( .DIN1(n600), .DIN2(n449), .Q(n3108) );
  nnd2s1 U3558 ( .DIN1(n3110), .DIN2(n3111), .Q(\IDinst/n5353 ) );
  nnd2s1 U3559 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][17] ), .Q(n3111) );
  nnd2s1 U3560 ( .DIN1(n602), .DIN2(n448), .Q(n3110) );
  nnd2s1 U3561 ( .DIN1(n3112), .DIN2(n3113), .Q(\IDinst/n5352 ) );
  nnd2s1 U3562 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][17] ), .Q(n3113) );
  nnd2s1 U3563 ( .DIN1(n588), .DIN2(n449), .Q(n3112) );
  nnd2s1 U3564 ( .DIN1(n3114), .DIN2(n3115), .Q(\IDinst/n5351 ) );
  nnd2s1 U3565 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][17] ), .Q(n3115) );
  nnd2s1 U3566 ( .DIN1(n590), .DIN2(n448), .Q(n3114) );
  nnd2s1 U3567 ( .DIN1(n3116), .DIN2(n3117), .Q(\IDinst/n5350 ) );
  nnd2s1 U3568 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][17] ), .Q(n3117) );
  nnd2s1 U3569 ( .DIN1(n592), .DIN2(n449), .Q(n3116) );
  nnd2s1 U3570 ( .DIN1(n3118), .DIN2(n3119), .Q(\IDinst/n5349 ) );
  nnd2s1 U3571 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][17] ), .Q(n3119) );
  nnd2s1 U3572 ( .DIN1(n594), .DIN2(n448), .Q(n3118) );
  nnd2s1 U3573 ( .DIN1(n3120), .DIN2(n3121), .Q(\IDinst/n5348 ) );
  nnd2s1 U3574 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][17] ), .Q(n3121) );
  nnd2s1 U3575 ( .DIN1(n612), .DIN2(n449), .Q(n3120) );
  nnd2s1 U3576 ( .DIN1(n3122), .DIN2(n3123), .Q(\IDinst/n5347 ) );
  nnd2s1 U3577 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][17] ), .Q(n3123) );
  nnd2s1 U3578 ( .DIN1(n614), .DIN2(n448), .Q(n3122) );
  nnd2s1 U3579 ( .DIN1(n3124), .DIN2(n3125), .Q(\IDinst/n5346 ) );
  nnd2s1 U3580 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][17] ), .Q(n3125) );
  nnd2s1 U3581 ( .DIN1(n616), .DIN2(n449), .Q(n3124) );
  nnd2s1 U3582 ( .DIN1(n3126), .DIN2(n3127), .Q(\IDinst/n5345 ) );
  nnd2s1 U3583 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][17] ), .Q(n3127) );
  nnd2s1 U3584 ( .DIN1(n618), .DIN2(n448), .Q(n3126) );
  nnd2s1 U3585 ( .DIN1(n3128), .DIN2(n3129), .Q(\IDinst/n5344 ) );
  nnd2s1 U3586 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][17] ), .Q(n3129) );
  nnd2s1 U3587 ( .DIN1(n604), .DIN2(n449), .Q(n3128) );
  nnd2s1 U3588 ( .DIN1(n3130), .DIN2(n3131), .Q(\IDinst/n5343 ) );
  nnd2s1 U3589 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][17] ), .Q(n3131) );
  nnd2s1 U3590 ( .DIN1(n606), .DIN2(n448), .Q(n3130) );
  nnd2s1 U3591 ( .DIN1(n3132), .DIN2(n3133), .Q(\IDinst/n5342 ) );
  nnd2s1 U3592 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][17] ), .Q(n3133) );
  nnd2s1 U3593 ( .DIN1(n608), .DIN2(n449), .Q(n3132) );
  nnd2s1 U3594 ( .DIN1(n3134), .DIN2(n3135), .Q(\IDinst/n5341 ) );
  nnd2s1 U3595 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][17] ), .Q(n3135) );
  nnd2s1 U3596 ( .DIN1(n610), .DIN2(n448), .Q(n3134) );
  nnd2s1 U3597 ( .DIN1(n3136), .DIN2(n3137), .Q(\IDinst/n5340 ) );
  nnd2s1 U3598 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][17] ), .Q(n3137) );
  nnd2s1 U3599 ( .DIN1(n580), .DIN2(n449), .Q(n3136) );
  nnd2s1 U3600 ( .DIN1(n3138), .DIN2(n3139), .Q(\IDinst/n5339 ) );
  nnd2s1 U3601 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][17] ), .Q(n3139) );
  nnd2s1 U3602 ( .DIN1(n582), .DIN2(n448), .Q(n3138) );
  nnd2s1 U3603 ( .DIN1(n3140), .DIN2(n3141), .Q(\IDinst/n5338 ) );
  nnd2s1 U3604 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][17] ), .Q(n3141) );
  nnd2s1 U3605 ( .DIN1(n584), .DIN2(n449), .Q(n3140) );
  nnd2s1 U3606 ( .DIN1(n3142), .DIN2(n3143), .Q(\IDinst/n5337 ) );
  nnd2s1 U3607 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][17] ), .Q(n3143) );
  nnd2s1 U3608 ( .DIN1(n586), .DIN2(n448), .Q(n3142) );
  nnd2s1 U3609 ( .DIN1(n3144), .DIN2(n3145), .Q(\IDinst/n5336 ) );
  nnd2s1 U3610 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][17] ), .Q(n3145) );
  nnd2s1 U3611 ( .DIN1(n572), .DIN2(n449), .Q(n3144) );
  nnd2s1 U3612 ( .DIN1(n3146), .DIN2(n3147), .Q(\IDinst/n5335 ) );
  nnd2s1 U3613 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][17] ), .Q(n3147) );
  nnd2s1 U3614 ( .DIN1(n574), .DIN2(n448), .Q(n3146) );
  nnd2s1 U3615 ( .DIN1(n3148), .DIN2(n3149), .Q(\IDinst/n5334 ) );
  nnd2s1 U3616 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][17] ), .Q(n3149) );
  nnd2s1 U3617 ( .DIN1(n576), .DIN2(n449), .Q(n3148) );
  nnd2s1 U3618 ( .DIN1(n3150), .DIN2(n3151), .Q(\IDinst/n5333 ) );
  nnd2s1 U3619 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][17] ), .Q(n3151) );
  nnd2s1 U3620 ( .DIN1(n578), .DIN2(n448), .Q(n3150) );
  nnd2s1 U3621 ( .DIN1(n3152), .DIN2(n3153), .Q(\IDinst/n5332 ) );
  nnd2s1 U3622 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][17] ), .Q(n3153) );
  nnd2s1 U3623 ( .DIN1(n564), .DIN2(n449), .Q(n3152) );
  nnd2s1 U3624 ( .DIN1(n3154), .DIN2(n3155), .Q(\IDinst/n5331 ) );
  nnd2s1 U3625 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][17] ), .Q(n3155) );
  nnd2s1 U3626 ( .DIN1(n566), .DIN2(n448), .Q(n3154) );
  nnd2s1 U3627 ( .DIN1(n3156), .DIN2(n3157), .Q(\IDinst/n5330 ) );
  nnd2s1 U3628 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][17] ), .Q(n3157) );
  nnd2s1 U3629 ( .DIN1(n568), .DIN2(n449), .Q(n3156) );
  nnd2s1 U3630 ( .DIN1(n3158), .DIN2(n3159), .Q(\IDinst/n5329 ) );
  nnd2s1 U3631 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][17] ), .Q(n3159) );
  nnd2s1 U3632 ( .DIN1(n570), .DIN2(n448), .Q(n3158) );
  nnd2s1 U3633 ( .DIN1(n3160), .DIN2(n3161), .Q(\IDinst/n5328 ) );
  nnd2s1 U3634 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][17] ), .Q(n3161) );
  nnd2s1 U3635 ( .DIN1(n556), .DIN2(n449), .Q(n3160) );
  nnd2s1 U3636 ( .DIN1(n3162), .DIN2(n3163), .Q(\IDinst/n5327 ) );
  nnd2s1 U3637 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][17] ), .Q(n3163) );
  nnd2s1 U3638 ( .DIN1(n558), .DIN2(n448), .Q(n3162) );
  nnd2s1 U3639 ( .DIN1(n3164), .DIN2(n3165), .Q(\IDinst/n5326 ) );
  nnd2s1 U3640 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][17] ), .Q(n3165) );
  nnd2s1 U3641 ( .DIN1(n560), .DIN2(n449), .Q(n3164) );
  nnd2s1 U3642 ( .DIN1(n3166), .DIN2(n3167), .Q(\IDinst/n5325 ) );
  nnd2s1 U3643 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][17] ), .Q(n3167) );
  nnd2s1 U3644 ( .DIN1(n562), .DIN2(n448), .Q(n3166) );
  nnd2s1 U3645 ( .DIN1(n3103), .DIN2(n183), .Q(n3168) );
  nnd2s1 U3646 ( .DIN1(n3169), .DIN2(n3170), .Q(\IDinst/n5324 ) );
  nnd2s1 U3647 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][18] ), .Q(n3170) );
  nnd2s1 U3648 ( .DIN1(n597), .DIN2(n451), .Q(n3169) );
  nnd2s1 U3649 ( .DIN1(n3171), .DIN2(n3172), .Q(\IDinst/n5323 ) );
  nnd2s1 U3650 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][18] ), .Q(n3172) );
  nnd2s1 U3651 ( .DIN1(n599), .DIN2(n450), .Q(n3171) );
  nnd2s1 U3652 ( .DIN1(n3173), .DIN2(n3174), .Q(\IDinst/n5322 ) );
  nnd2s1 U3653 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][18] ), .Q(n3174) );
  nnd2s1 U3654 ( .DIN1(n601), .DIN2(n451), .Q(n3173) );
  nnd2s1 U3655 ( .DIN1(n3175), .DIN2(n3176), .Q(\IDinst/n5321 ) );
  nnd2s1 U3656 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][18] ), .Q(n3176) );
  nnd2s1 U3657 ( .DIN1(n603), .DIN2(n450), .Q(n3175) );
  nnd2s1 U3658 ( .DIN1(n3177), .DIN2(n3178), .Q(\IDinst/n5320 ) );
  nnd2s1 U3659 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][18] ), .Q(n3178) );
  nnd2s1 U3660 ( .DIN1(n589), .DIN2(n451), .Q(n3177) );
  nnd2s1 U3661 ( .DIN1(n3179), .DIN2(n3180), .Q(\IDinst/n5319 ) );
  nnd2s1 U3662 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][18] ), .Q(n3180) );
  nnd2s1 U3663 ( .DIN1(n591), .DIN2(n450), .Q(n3179) );
  nnd2s1 U3664 ( .DIN1(n3181), .DIN2(n3182), .Q(\IDinst/n5318 ) );
  nnd2s1 U3665 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][18] ), .Q(n3182) );
  nnd2s1 U3666 ( .DIN1(n593), .DIN2(n451), .Q(n3181) );
  nnd2s1 U3667 ( .DIN1(n3183), .DIN2(n3184), .Q(\IDinst/n5317 ) );
  nnd2s1 U3668 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][18] ), .Q(n3184) );
  nnd2s1 U3669 ( .DIN1(n595), .DIN2(n450), .Q(n3183) );
  nnd2s1 U3670 ( .DIN1(n3185), .DIN2(n3186), .Q(\IDinst/n5316 ) );
  nnd2s1 U3671 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][18] ), .Q(n3186) );
  nnd2s1 U3672 ( .DIN1(n613), .DIN2(n451), .Q(n3185) );
  nnd2s1 U3673 ( .DIN1(n3187), .DIN2(n3188), .Q(\IDinst/n5315 ) );
  nnd2s1 U3674 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][18] ), .Q(n3188) );
  nnd2s1 U3675 ( .DIN1(n615), .DIN2(n450), .Q(n3187) );
  nnd2s1 U3676 ( .DIN1(n3189), .DIN2(n3190), .Q(\IDinst/n5314 ) );
  nnd2s1 U3677 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][18] ), .Q(n3190) );
  nnd2s1 U3678 ( .DIN1(n617), .DIN2(n451), .Q(n3189) );
  nnd2s1 U3679 ( .DIN1(n3191), .DIN2(n3192), .Q(\IDinst/n5313 ) );
  nnd2s1 U3680 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][18] ), .Q(n3192) );
  nnd2s1 U3681 ( .DIN1(n619), .DIN2(n450), .Q(n3191) );
  nnd2s1 U3682 ( .DIN1(n3193), .DIN2(n3194), .Q(\IDinst/n5312 ) );
  nnd2s1 U3683 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][18] ), .Q(n3194) );
  nnd2s1 U3684 ( .DIN1(n605), .DIN2(n451), .Q(n3193) );
  nnd2s1 U3685 ( .DIN1(n3195), .DIN2(n3196), .Q(\IDinst/n5311 ) );
  nnd2s1 U3686 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][18] ), .Q(n3196) );
  nnd2s1 U3687 ( .DIN1(n607), .DIN2(n450), .Q(n3195) );
  nnd2s1 U3688 ( .DIN1(n3197), .DIN2(n3198), .Q(\IDinst/n5310 ) );
  nnd2s1 U3689 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][18] ), .Q(n3198) );
  nnd2s1 U3690 ( .DIN1(n609), .DIN2(n451), .Q(n3197) );
  nnd2s1 U3691 ( .DIN1(n3199), .DIN2(n3200), .Q(\IDinst/n5309 ) );
  nnd2s1 U3692 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][18] ), .Q(n3200) );
  nnd2s1 U3693 ( .DIN1(n611), .DIN2(n450), .Q(n3199) );
  nnd2s1 U3694 ( .DIN1(n3201), .DIN2(n3202), .Q(\IDinst/n5308 ) );
  nnd2s1 U3695 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][18] ), .Q(n3202) );
  nnd2s1 U3696 ( .DIN1(n581), .DIN2(n451), .Q(n3201) );
  nnd2s1 U3697 ( .DIN1(n3203), .DIN2(n3204), .Q(\IDinst/n5307 ) );
  nnd2s1 U3698 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][18] ), .Q(n3204) );
  nnd2s1 U3699 ( .DIN1(n583), .DIN2(n450), .Q(n3203) );
  nnd2s1 U3700 ( .DIN1(n3205), .DIN2(n3206), .Q(\IDinst/n5306 ) );
  nnd2s1 U3701 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][18] ), .Q(n3206) );
  nnd2s1 U3702 ( .DIN1(n585), .DIN2(n451), .Q(n3205) );
  nnd2s1 U3703 ( .DIN1(n3207), .DIN2(n3208), .Q(\IDinst/n5305 ) );
  nnd2s1 U3704 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][18] ), .Q(n3208) );
  nnd2s1 U3705 ( .DIN1(n587), .DIN2(n450), .Q(n3207) );
  nnd2s1 U3706 ( .DIN1(n3209), .DIN2(n3210), .Q(\IDinst/n5304 ) );
  nnd2s1 U3707 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][18] ), .Q(n3210) );
  nnd2s1 U3708 ( .DIN1(n573), .DIN2(n451), .Q(n3209) );
  nnd2s1 U3709 ( .DIN1(n3211), .DIN2(n3212), .Q(\IDinst/n5303 ) );
  nnd2s1 U3710 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][18] ), .Q(n3212) );
  nnd2s1 U3711 ( .DIN1(n575), .DIN2(n450), .Q(n3211) );
  nnd2s1 U3712 ( .DIN1(n3213), .DIN2(n3214), .Q(\IDinst/n5302 ) );
  nnd2s1 U3713 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][18] ), .Q(n3214) );
  nnd2s1 U3714 ( .DIN1(n577), .DIN2(n451), .Q(n3213) );
  nnd2s1 U3715 ( .DIN1(n3215), .DIN2(n3216), .Q(\IDinst/n5301 ) );
  nnd2s1 U3716 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][18] ), .Q(n3216) );
  nnd2s1 U3717 ( .DIN1(n579), .DIN2(n450), .Q(n3215) );
  nnd2s1 U3718 ( .DIN1(n3217), .DIN2(n3218), .Q(\IDinst/n5300 ) );
  nnd2s1 U3719 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][18] ), .Q(n3218) );
  nnd2s1 U3720 ( .DIN1(n565), .DIN2(n451), .Q(n3217) );
  nnd2s1 U3721 ( .DIN1(n3219), .DIN2(n3220), .Q(\IDinst/n5299 ) );
  nnd2s1 U3722 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][18] ), .Q(n3220) );
  nnd2s1 U3723 ( .DIN1(n567), .DIN2(n450), .Q(n3219) );
  nnd2s1 U3724 ( .DIN1(n3221), .DIN2(n3222), .Q(\IDinst/n5298 ) );
  nnd2s1 U3725 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][18] ), .Q(n3222) );
  nnd2s1 U3726 ( .DIN1(n569), .DIN2(n451), .Q(n3221) );
  nnd2s1 U3727 ( .DIN1(n3223), .DIN2(n3224), .Q(\IDinst/n5297 ) );
  nnd2s1 U3728 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][18] ), .Q(n3224) );
  nnd2s1 U3729 ( .DIN1(n571), .DIN2(n450), .Q(n3223) );
  nnd2s1 U3730 ( .DIN1(n3225), .DIN2(n3226), .Q(\IDinst/n5296 ) );
  nnd2s1 U3731 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][18] ), .Q(n3226) );
  nnd2s1 U3732 ( .DIN1(n557), .DIN2(n451), .Q(n3225) );
  nnd2s1 U3733 ( .DIN1(n3227), .DIN2(n3228), .Q(\IDinst/n5295 ) );
  nnd2s1 U3734 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][18] ), .Q(n3228) );
  nnd2s1 U3735 ( .DIN1(n559), .DIN2(n450), .Q(n3227) );
  nnd2s1 U3736 ( .DIN1(n3229), .DIN2(n3230), .Q(\IDinst/n5294 ) );
  nnd2s1 U3737 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][18] ), .Q(n3230) );
  nnd2s1 U3738 ( .DIN1(n561), .DIN2(n451), .Q(n3229) );
  nnd2s1 U3739 ( .DIN1(n3231), .DIN2(n3232), .Q(\IDinst/n5293 ) );
  nnd2s1 U3740 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][18] ), .Q(n3232) );
  nnd2s1 U3741 ( .DIN1(n563), .DIN2(n450), .Q(n3231) );
  nnd2s1 U3742 ( .DIN1(n3103), .DIN2(n181), .Q(n3233) );
  nnd2s1 U3743 ( .DIN1(n3234), .DIN2(n3235), .Q(\IDinst/n5292 ) );
  nnd2s1 U3744 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][19] ), .Q(n3235) );
  nnd2s1 U3745 ( .DIN1(n596), .DIN2(n453), .Q(n3234) );
  nnd2s1 U3746 ( .DIN1(n3236), .DIN2(n3237), .Q(\IDinst/n5291 ) );
  nnd2s1 U3747 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][19] ), .Q(n3237) );
  nnd2s1 U3748 ( .DIN1(n598), .DIN2(n452), .Q(n3236) );
  nnd2s1 U3749 ( .DIN1(n3238), .DIN2(n3239), .Q(\IDinst/n5290 ) );
  nnd2s1 U3750 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][19] ), .Q(n3239) );
  nnd2s1 U3751 ( .DIN1(n600), .DIN2(n453), .Q(n3238) );
  nnd2s1 U3752 ( .DIN1(n3240), .DIN2(n3241), .Q(\IDinst/n5289 ) );
  nnd2s1 U3753 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][19] ), .Q(n3241) );
  nnd2s1 U3754 ( .DIN1(n602), .DIN2(n452), .Q(n3240) );
  nnd2s1 U3755 ( .DIN1(n3242), .DIN2(n3243), .Q(\IDinst/n5288 ) );
  nnd2s1 U3756 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][19] ), .Q(n3243) );
  nnd2s1 U3757 ( .DIN1(n588), .DIN2(n453), .Q(n3242) );
  nnd2s1 U3758 ( .DIN1(n3244), .DIN2(n3245), .Q(\IDinst/n5287 ) );
  nnd2s1 U3759 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][19] ), .Q(n3245) );
  nnd2s1 U3760 ( .DIN1(n590), .DIN2(n452), .Q(n3244) );
  nnd2s1 U3761 ( .DIN1(n3246), .DIN2(n3247), .Q(\IDinst/n5286 ) );
  nnd2s1 U3762 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][19] ), .Q(n3247) );
  nnd2s1 U3763 ( .DIN1(n592), .DIN2(n453), .Q(n3246) );
  nnd2s1 U3764 ( .DIN1(n3248), .DIN2(n3249), .Q(\IDinst/n5285 ) );
  nnd2s1 U3765 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][19] ), .Q(n3249) );
  nnd2s1 U3766 ( .DIN1(n594), .DIN2(n452), .Q(n3248) );
  nnd2s1 U3767 ( .DIN1(n3250), .DIN2(n3251), .Q(\IDinst/n5284 ) );
  nnd2s1 U3768 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][19] ), .Q(n3251) );
  nnd2s1 U3769 ( .DIN1(n612), .DIN2(n453), .Q(n3250) );
  nnd2s1 U3770 ( .DIN1(n3252), .DIN2(n3253), .Q(\IDinst/n5283 ) );
  nnd2s1 U3771 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][19] ), .Q(n3253) );
  nnd2s1 U3772 ( .DIN1(n614), .DIN2(n452), .Q(n3252) );
  nnd2s1 U3773 ( .DIN1(n3254), .DIN2(n3255), .Q(\IDinst/n5282 ) );
  nnd2s1 U3774 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][19] ), .Q(n3255) );
  nnd2s1 U3775 ( .DIN1(n616), .DIN2(n453), .Q(n3254) );
  nnd2s1 U3776 ( .DIN1(n3256), .DIN2(n3257), .Q(\IDinst/n5281 ) );
  nnd2s1 U3777 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][19] ), .Q(n3257) );
  nnd2s1 U3778 ( .DIN1(n618), .DIN2(n452), .Q(n3256) );
  nnd2s1 U3779 ( .DIN1(n3258), .DIN2(n3259), .Q(\IDinst/n5280 ) );
  nnd2s1 U3780 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][19] ), .Q(n3259) );
  nnd2s1 U3781 ( .DIN1(n604), .DIN2(n453), .Q(n3258) );
  nnd2s1 U3782 ( .DIN1(n3260), .DIN2(n3261), .Q(\IDinst/n5279 ) );
  nnd2s1 U3783 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][19] ), .Q(n3261) );
  nnd2s1 U3784 ( .DIN1(n606), .DIN2(n452), .Q(n3260) );
  nnd2s1 U3785 ( .DIN1(n3262), .DIN2(n3263), .Q(\IDinst/n5278 ) );
  nnd2s1 U3786 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][19] ), .Q(n3263) );
  nnd2s1 U3787 ( .DIN1(n608), .DIN2(n453), .Q(n3262) );
  nnd2s1 U3788 ( .DIN1(n3264), .DIN2(n3265), .Q(\IDinst/n5277 ) );
  nnd2s1 U3789 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][19] ), .Q(n3265) );
  nnd2s1 U3790 ( .DIN1(n610), .DIN2(n452), .Q(n3264) );
  nnd2s1 U3791 ( .DIN1(n3266), .DIN2(n3267), .Q(\IDinst/n5276 ) );
  nnd2s1 U3792 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][19] ), .Q(n3267) );
  nnd2s1 U3793 ( .DIN1(n580), .DIN2(n453), .Q(n3266) );
  nnd2s1 U3794 ( .DIN1(n3268), .DIN2(n3269), .Q(\IDinst/n5275 ) );
  nnd2s1 U3795 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][19] ), .Q(n3269) );
  nnd2s1 U3796 ( .DIN1(n582), .DIN2(n452), .Q(n3268) );
  nnd2s1 U3797 ( .DIN1(n3270), .DIN2(n3271), .Q(\IDinst/n5274 ) );
  nnd2s1 U3798 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][19] ), .Q(n3271) );
  nnd2s1 U3799 ( .DIN1(n584), .DIN2(n453), .Q(n3270) );
  nnd2s1 U3800 ( .DIN1(n3272), .DIN2(n3273), .Q(\IDinst/n5273 ) );
  nnd2s1 U3801 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][19] ), .Q(n3273) );
  nnd2s1 U3802 ( .DIN1(n586), .DIN2(n452), .Q(n3272) );
  nnd2s1 U3803 ( .DIN1(n3274), .DIN2(n3275), .Q(\IDinst/n5272 ) );
  nnd2s1 U3804 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][19] ), .Q(n3275) );
  nnd2s1 U3805 ( .DIN1(n572), .DIN2(n453), .Q(n3274) );
  nnd2s1 U3806 ( .DIN1(n3276), .DIN2(n3277), .Q(\IDinst/n5271 ) );
  nnd2s1 U3807 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][19] ), .Q(n3277) );
  nnd2s1 U3808 ( .DIN1(n574), .DIN2(n452), .Q(n3276) );
  nnd2s1 U3809 ( .DIN1(n3278), .DIN2(n3279), .Q(\IDinst/n5270 ) );
  nnd2s1 U3810 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][19] ), .Q(n3279) );
  nnd2s1 U3811 ( .DIN1(n576), .DIN2(n453), .Q(n3278) );
  nnd2s1 U3812 ( .DIN1(n3280), .DIN2(n3281), .Q(\IDinst/n5269 ) );
  nnd2s1 U3813 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][19] ), .Q(n3281) );
  nnd2s1 U3814 ( .DIN1(n578), .DIN2(n452), .Q(n3280) );
  nnd2s1 U3815 ( .DIN1(n3282), .DIN2(n3283), .Q(\IDinst/n5268 ) );
  nnd2s1 U3816 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][19] ), .Q(n3283) );
  nnd2s1 U3817 ( .DIN1(n564), .DIN2(n453), .Q(n3282) );
  nnd2s1 U3818 ( .DIN1(n3284), .DIN2(n3285), .Q(\IDinst/n5267 ) );
  nnd2s1 U3819 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][19] ), .Q(n3285) );
  nnd2s1 U3820 ( .DIN1(n566), .DIN2(n452), .Q(n3284) );
  nnd2s1 U3821 ( .DIN1(n3286), .DIN2(n3287), .Q(\IDinst/n5266 ) );
  nnd2s1 U3822 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][19] ), .Q(n3287) );
  nnd2s1 U3823 ( .DIN1(n568), .DIN2(n453), .Q(n3286) );
  nnd2s1 U3824 ( .DIN1(n3288), .DIN2(n3289), .Q(\IDinst/n5265 ) );
  nnd2s1 U3825 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][19] ), .Q(n3289) );
  nnd2s1 U3826 ( .DIN1(n570), .DIN2(n452), .Q(n3288) );
  nnd2s1 U3827 ( .DIN1(n3290), .DIN2(n3291), .Q(\IDinst/n5264 ) );
  nnd2s1 U3828 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][19] ), .Q(n3291) );
  nnd2s1 U3829 ( .DIN1(n556), .DIN2(n453), .Q(n3290) );
  nnd2s1 U3830 ( .DIN1(n3292), .DIN2(n3293), .Q(\IDinst/n5263 ) );
  nnd2s1 U3831 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][19] ), .Q(n3293) );
  nnd2s1 U3832 ( .DIN1(n558), .DIN2(n452), .Q(n3292) );
  nnd2s1 U3833 ( .DIN1(n3294), .DIN2(n3295), .Q(\IDinst/n5262 ) );
  nnd2s1 U3834 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][19] ), .Q(n3295) );
  nnd2s1 U3835 ( .DIN1(n560), .DIN2(n453), .Q(n3294) );
  nnd2s1 U3836 ( .DIN1(n3296), .DIN2(n3297), .Q(\IDinst/n5261 ) );
  nnd2s1 U3837 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][19] ), .Q(n3297) );
  nnd2s1 U3838 ( .DIN1(n562), .DIN2(n452), .Q(n3296) );
  nnd2s1 U3839 ( .DIN1(n3103), .DIN2(n179), .Q(n3298) );
  nnd2s1 U3840 ( .DIN1(n3299), .DIN2(n3300), .Q(\IDinst/n5260 ) );
  nnd2s1 U3841 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][20] ), .Q(n3300) );
  nnd2s1 U3842 ( .DIN1(n597), .DIN2(n455), .Q(n3299) );
  nnd2s1 U3843 ( .DIN1(n3301), .DIN2(n3302), .Q(\IDinst/n5259 ) );
  nnd2s1 U3844 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][20] ), .Q(n3302) );
  nnd2s1 U3845 ( .DIN1(n599), .DIN2(n454), .Q(n3301) );
  nnd2s1 U3846 ( .DIN1(n3303), .DIN2(n3304), .Q(\IDinst/n5258 ) );
  nnd2s1 U3847 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][20] ), .Q(n3304) );
  nnd2s1 U3848 ( .DIN1(n601), .DIN2(n455), .Q(n3303) );
  nnd2s1 U3849 ( .DIN1(n3305), .DIN2(n3306), .Q(\IDinst/n5257 ) );
  nnd2s1 U3850 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][20] ), .Q(n3306) );
  nnd2s1 U3851 ( .DIN1(n603), .DIN2(n454), .Q(n3305) );
  nnd2s1 U3852 ( .DIN1(n3307), .DIN2(n3308), .Q(\IDinst/n5256 ) );
  nnd2s1 U3853 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][20] ), .Q(n3308) );
  nnd2s1 U3854 ( .DIN1(n589), .DIN2(n455), .Q(n3307) );
  nnd2s1 U3855 ( .DIN1(n3309), .DIN2(n3310), .Q(\IDinst/n5255 ) );
  nnd2s1 U3856 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][20] ), .Q(n3310) );
  nnd2s1 U3857 ( .DIN1(n591), .DIN2(n454), .Q(n3309) );
  nnd2s1 U3858 ( .DIN1(n3311), .DIN2(n3312), .Q(\IDinst/n5254 ) );
  nnd2s1 U3859 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][20] ), .Q(n3312) );
  nnd2s1 U3860 ( .DIN1(n593), .DIN2(n455), .Q(n3311) );
  nnd2s1 U3861 ( .DIN1(n3313), .DIN2(n3314), .Q(\IDinst/n5253 ) );
  nnd2s1 U3862 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][20] ), .Q(n3314) );
  nnd2s1 U3863 ( .DIN1(n595), .DIN2(n454), .Q(n3313) );
  nnd2s1 U3864 ( .DIN1(n3315), .DIN2(n3316), .Q(\IDinst/n5252 ) );
  nnd2s1 U3865 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][20] ), .Q(n3316) );
  nnd2s1 U3866 ( .DIN1(n613), .DIN2(n455), .Q(n3315) );
  nnd2s1 U3867 ( .DIN1(n3317), .DIN2(n3318), .Q(\IDinst/n5251 ) );
  nnd2s1 U3868 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][20] ), .Q(n3318) );
  nnd2s1 U3869 ( .DIN1(n615), .DIN2(n454), .Q(n3317) );
  nnd2s1 U3870 ( .DIN1(n3319), .DIN2(n3320), .Q(\IDinst/n5250 ) );
  nnd2s1 U3871 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][20] ), .Q(n3320) );
  nnd2s1 U3872 ( .DIN1(n617), .DIN2(n455), .Q(n3319) );
  nnd2s1 U3873 ( .DIN1(n3321), .DIN2(n3322), .Q(\IDinst/n5249 ) );
  nnd2s1 U3874 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][20] ), .Q(n3322) );
  nnd2s1 U3875 ( .DIN1(n619), .DIN2(n454), .Q(n3321) );
  nnd2s1 U3876 ( .DIN1(n3323), .DIN2(n3324), .Q(\IDinst/n5248 ) );
  nnd2s1 U3877 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][20] ), .Q(n3324) );
  nnd2s1 U3878 ( .DIN1(n605), .DIN2(n455), .Q(n3323) );
  nnd2s1 U3879 ( .DIN1(n3325), .DIN2(n3326), .Q(\IDinst/n5247 ) );
  nnd2s1 U3880 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][20] ), .Q(n3326) );
  nnd2s1 U3881 ( .DIN1(n607), .DIN2(n454), .Q(n3325) );
  nnd2s1 U3882 ( .DIN1(n3327), .DIN2(n3328), .Q(\IDinst/n5246 ) );
  nnd2s1 U3883 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][20] ), .Q(n3328) );
  nnd2s1 U3884 ( .DIN1(n609), .DIN2(n455), .Q(n3327) );
  nnd2s1 U3885 ( .DIN1(n3329), .DIN2(n3330), .Q(\IDinst/n5245 ) );
  nnd2s1 U3886 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][20] ), .Q(n3330) );
  nnd2s1 U3887 ( .DIN1(n611), .DIN2(n454), .Q(n3329) );
  nnd2s1 U3888 ( .DIN1(n3331), .DIN2(n3332), .Q(\IDinst/n5244 ) );
  nnd2s1 U3889 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][20] ), .Q(n3332) );
  nnd2s1 U3890 ( .DIN1(n581), .DIN2(n455), .Q(n3331) );
  nnd2s1 U3891 ( .DIN1(n3333), .DIN2(n3334), .Q(\IDinst/n5243 ) );
  nnd2s1 U3892 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][20] ), .Q(n3334) );
  nnd2s1 U3893 ( .DIN1(n583), .DIN2(n454), .Q(n3333) );
  nnd2s1 U3894 ( .DIN1(n3335), .DIN2(n3336), .Q(\IDinst/n5242 ) );
  nnd2s1 U3895 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][20] ), .Q(n3336) );
  nnd2s1 U3896 ( .DIN1(n585), .DIN2(n455), .Q(n3335) );
  nnd2s1 U3897 ( .DIN1(n3337), .DIN2(n3338), .Q(\IDinst/n5241 ) );
  nnd2s1 U3898 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][20] ), .Q(n3338) );
  nnd2s1 U3899 ( .DIN1(n587), .DIN2(n454), .Q(n3337) );
  nnd2s1 U3900 ( .DIN1(n3339), .DIN2(n3340), .Q(\IDinst/n5240 ) );
  nnd2s1 U3901 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][20] ), .Q(n3340) );
  nnd2s1 U3902 ( .DIN1(n573), .DIN2(n455), .Q(n3339) );
  nnd2s1 U3903 ( .DIN1(n3341), .DIN2(n3342), .Q(\IDinst/n5239 ) );
  nnd2s1 U3904 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][20] ), .Q(n3342) );
  nnd2s1 U3905 ( .DIN1(n575), .DIN2(n454), .Q(n3341) );
  nnd2s1 U3906 ( .DIN1(n3343), .DIN2(n3344), .Q(\IDinst/n5238 ) );
  nnd2s1 U3907 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][20] ), .Q(n3344) );
  nnd2s1 U3908 ( .DIN1(n577), .DIN2(n455), .Q(n3343) );
  nnd2s1 U3909 ( .DIN1(n3345), .DIN2(n3346), .Q(\IDinst/n5237 ) );
  nnd2s1 U3910 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][20] ), .Q(n3346) );
  nnd2s1 U3911 ( .DIN1(n579), .DIN2(n454), .Q(n3345) );
  nnd2s1 U3912 ( .DIN1(n3347), .DIN2(n3348), .Q(\IDinst/n5236 ) );
  nnd2s1 U3913 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][20] ), .Q(n3348) );
  nnd2s1 U3914 ( .DIN1(n565), .DIN2(n455), .Q(n3347) );
  nnd2s1 U3915 ( .DIN1(n3349), .DIN2(n3350), .Q(\IDinst/n5235 ) );
  nnd2s1 U3916 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][20] ), .Q(n3350) );
  nnd2s1 U3917 ( .DIN1(n567), .DIN2(n454), .Q(n3349) );
  nnd2s1 U3918 ( .DIN1(n3351), .DIN2(n3352), .Q(\IDinst/n5234 ) );
  nnd2s1 U3919 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][20] ), .Q(n3352) );
  nnd2s1 U3920 ( .DIN1(n569), .DIN2(n455), .Q(n3351) );
  nnd2s1 U3921 ( .DIN1(n3353), .DIN2(n3354), .Q(\IDinst/n5233 ) );
  nnd2s1 U3922 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][20] ), .Q(n3354) );
  nnd2s1 U3923 ( .DIN1(n571), .DIN2(n454), .Q(n3353) );
  nnd2s1 U3924 ( .DIN1(n3355), .DIN2(n3356), .Q(\IDinst/n5232 ) );
  nnd2s1 U3925 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][20] ), .Q(n3356) );
  nnd2s1 U3926 ( .DIN1(n557), .DIN2(n455), .Q(n3355) );
  nnd2s1 U3927 ( .DIN1(n3357), .DIN2(n3358), .Q(\IDinst/n5231 ) );
  nnd2s1 U3928 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][20] ), .Q(n3358) );
  nnd2s1 U3929 ( .DIN1(n559), .DIN2(n454), .Q(n3357) );
  nnd2s1 U3930 ( .DIN1(n3359), .DIN2(n3360), .Q(\IDinst/n5230 ) );
  nnd2s1 U3931 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][20] ), .Q(n3360) );
  nnd2s1 U3932 ( .DIN1(n561), .DIN2(n455), .Q(n3359) );
  nnd2s1 U3933 ( .DIN1(n3361), .DIN2(n3362), .Q(\IDinst/n5229 ) );
  nnd2s1 U3934 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][20] ), .Q(n3362) );
  nnd2s1 U3935 ( .DIN1(n563), .DIN2(n454), .Q(n3361) );
  nnd2s1 U3936 ( .DIN1(n3103), .DIN2(n177), .Q(n3363) );
  nnd2s1 U3937 ( .DIN1(n3364), .DIN2(n3365), .Q(\IDinst/n5228 ) );
  nnd2s1 U3938 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][21] ), .Q(n3365) );
  nnd2s1 U3939 ( .DIN1(n596), .DIN2(n457), .Q(n3364) );
  nnd2s1 U3940 ( .DIN1(n3366), .DIN2(n3367), .Q(\IDinst/n5227 ) );
  nnd2s1 U3941 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][21] ), .Q(n3367) );
  nnd2s1 U3942 ( .DIN1(n598), .DIN2(n456), .Q(n3366) );
  nnd2s1 U3943 ( .DIN1(n3368), .DIN2(n3369), .Q(\IDinst/n5226 ) );
  nnd2s1 U3944 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][21] ), .Q(n3369) );
  nnd2s1 U3945 ( .DIN1(n600), .DIN2(n457), .Q(n3368) );
  nnd2s1 U3946 ( .DIN1(n3370), .DIN2(n3371), .Q(\IDinst/n5225 ) );
  nnd2s1 U3947 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][21] ), .Q(n3371) );
  nnd2s1 U3948 ( .DIN1(n602), .DIN2(n456), .Q(n3370) );
  nnd2s1 U3949 ( .DIN1(n3372), .DIN2(n3373), .Q(\IDinst/n5224 ) );
  nnd2s1 U3950 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][21] ), .Q(n3373) );
  nnd2s1 U3951 ( .DIN1(n588), .DIN2(n457), .Q(n3372) );
  nnd2s1 U3952 ( .DIN1(n3374), .DIN2(n3375), .Q(\IDinst/n5223 ) );
  nnd2s1 U3953 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][21] ), .Q(n3375) );
  nnd2s1 U3954 ( .DIN1(n590), .DIN2(n456), .Q(n3374) );
  nnd2s1 U3955 ( .DIN1(n3376), .DIN2(n3377), .Q(\IDinst/n5222 ) );
  nnd2s1 U3956 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][21] ), .Q(n3377) );
  nnd2s1 U3957 ( .DIN1(n592), .DIN2(n457), .Q(n3376) );
  nnd2s1 U3958 ( .DIN1(n3378), .DIN2(n3379), .Q(\IDinst/n5221 ) );
  nnd2s1 U3959 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][21] ), .Q(n3379) );
  nnd2s1 U3960 ( .DIN1(n594), .DIN2(n456), .Q(n3378) );
  nnd2s1 U3961 ( .DIN1(n3380), .DIN2(n3381), .Q(\IDinst/n5220 ) );
  nnd2s1 U3962 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][21] ), .Q(n3381) );
  nnd2s1 U3963 ( .DIN1(n612), .DIN2(n457), .Q(n3380) );
  nnd2s1 U3964 ( .DIN1(n3382), .DIN2(n3383), .Q(\IDinst/n5219 ) );
  nnd2s1 U3965 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][21] ), .Q(n3383) );
  nnd2s1 U3966 ( .DIN1(n614), .DIN2(n456), .Q(n3382) );
  nnd2s1 U3967 ( .DIN1(n3384), .DIN2(n3385), .Q(\IDinst/n5218 ) );
  nnd2s1 U3968 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][21] ), .Q(n3385) );
  nnd2s1 U3969 ( .DIN1(n616), .DIN2(n457), .Q(n3384) );
  nnd2s1 U3970 ( .DIN1(n3386), .DIN2(n3387), .Q(\IDinst/n5217 ) );
  nnd2s1 U3971 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][21] ), .Q(n3387) );
  nnd2s1 U3972 ( .DIN1(n618), .DIN2(n456), .Q(n3386) );
  nnd2s1 U3973 ( .DIN1(n3388), .DIN2(n3389), .Q(\IDinst/n5216 ) );
  nnd2s1 U3974 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][21] ), .Q(n3389) );
  nnd2s1 U3975 ( .DIN1(n604), .DIN2(n457), .Q(n3388) );
  nnd2s1 U3976 ( .DIN1(n3390), .DIN2(n3391), .Q(\IDinst/n5215 ) );
  nnd2s1 U3977 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][21] ), .Q(n3391) );
  nnd2s1 U3978 ( .DIN1(n606), .DIN2(n456), .Q(n3390) );
  nnd2s1 U3979 ( .DIN1(n3392), .DIN2(n3393), .Q(\IDinst/n5214 ) );
  nnd2s1 U3980 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][21] ), .Q(n3393) );
  nnd2s1 U3981 ( .DIN1(n608), .DIN2(n457), .Q(n3392) );
  nnd2s1 U3982 ( .DIN1(n3394), .DIN2(n3395), .Q(\IDinst/n5213 ) );
  nnd2s1 U3983 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][21] ), .Q(n3395) );
  nnd2s1 U3984 ( .DIN1(n610), .DIN2(n456), .Q(n3394) );
  nnd2s1 U3985 ( .DIN1(n3396), .DIN2(n3397), .Q(\IDinst/n5212 ) );
  nnd2s1 U3986 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][21] ), .Q(n3397) );
  nnd2s1 U3987 ( .DIN1(n580), .DIN2(n457), .Q(n3396) );
  nnd2s1 U3988 ( .DIN1(n3398), .DIN2(n3399), .Q(\IDinst/n5211 ) );
  nnd2s1 U3989 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][21] ), .Q(n3399) );
  nnd2s1 U3990 ( .DIN1(n582), .DIN2(n456), .Q(n3398) );
  nnd2s1 U3991 ( .DIN1(n3400), .DIN2(n3401), .Q(\IDinst/n5210 ) );
  nnd2s1 U3992 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][21] ), .Q(n3401) );
  nnd2s1 U3993 ( .DIN1(n584), .DIN2(n457), .Q(n3400) );
  nnd2s1 U3994 ( .DIN1(n3402), .DIN2(n3403), .Q(\IDinst/n5209 ) );
  nnd2s1 U3995 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][21] ), .Q(n3403) );
  nnd2s1 U3996 ( .DIN1(n586), .DIN2(n456), .Q(n3402) );
  nnd2s1 U3997 ( .DIN1(n3404), .DIN2(n3405), .Q(\IDinst/n5208 ) );
  nnd2s1 U3998 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][21] ), .Q(n3405) );
  nnd2s1 U3999 ( .DIN1(n572), .DIN2(n457), .Q(n3404) );
  nnd2s1 U4000 ( .DIN1(n3406), .DIN2(n3407), .Q(\IDinst/n5207 ) );
  nnd2s1 U4001 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][21] ), .Q(n3407) );
  nnd2s1 U4002 ( .DIN1(n574), .DIN2(n456), .Q(n3406) );
  nnd2s1 U4003 ( .DIN1(n3408), .DIN2(n3409), .Q(\IDinst/n5206 ) );
  nnd2s1 U4004 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][21] ), .Q(n3409) );
  nnd2s1 U4005 ( .DIN1(n576), .DIN2(n457), .Q(n3408) );
  nnd2s1 U4006 ( .DIN1(n3410), .DIN2(n3411), .Q(\IDinst/n5205 ) );
  nnd2s1 U4007 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][21] ), .Q(n3411) );
  nnd2s1 U4008 ( .DIN1(n578), .DIN2(n456), .Q(n3410) );
  nnd2s1 U4009 ( .DIN1(n3412), .DIN2(n3413), .Q(\IDinst/n5204 ) );
  nnd2s1 U4010 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][21] ), .Q(n3413) );
  nnd2s1 U4011 ( .DIN1(n564), .DIN2(n457), .Q(n3412) );
  nnd2s1 U4012 ( .DIN1(n3414), .DIN2(n3415), .Q(\IDinst/n5203 ) );
  nnd2s1 U4013 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][21] ), .Q(n3415) );
  nnd2s1 U4014 ( .DIN1(n566), .DIN2(n456), .Q(n3414) );
  nnd2s1 U4015 ( .DIN1(n3416), .DIN2(n3417), .Q(\IDinst/n5202 ) );
  nnd2s1 U4016 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][21] ), .Q(n3417) );
  nnd2s1 U4017 ( .DIN1(n568), .DIN2(n457), .Q(n3416) );
  nnd2s1 U4018 ( .DIN1(n3418), .DIN2(n3419), .Q(\IDinst/n5201 ) );
  nnd2s1 U4019 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][21] ), .Q(n3419) );
  nnd2s1 U4020 ( .DIN1(n570), .DIN2(n456), .Q(n3418) );
  nnd2s1 U4021 ( .DIN1(n3420), .DIN2(n3421), .Q(\IDinst/n5200 ) );
  nnd2s1 U4022 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][21] ), .Q(n3421) );
  nnd2s1 U4023 ( .DIN1(n556), .DIN2(n457), .Q(n3420) );
  nnd2s1 U4024 ( .DIN1(n3422), .DIN2(n3423), .Q(\IDinst/n5199 ) );
  nnd2s1 U4025 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][21] ), .Q(n3423) );
  nnd2s1 U4026 ( .DIN1(n558), .DIN2(n456), .Q(n3422) );
  nnd2s1 U4027 ( .DIN1(n3424), .DIN2(n3425), .Q(\IDinst/n5198 ) );
  nnd2s1 U4028 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][21] ), .Q(n3425) );
  nnd2s1 U4029 ( .DIN1(n560), .DIN2(n457), .Q(n3424) );
  nnd2s1 U4030 ( .DIN1(n3426), .DIN2(n3427), .Q(\IDinst/n5197 ) );
  nnd2s1 U4031 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][21] ), .Q(n3427) );
  nnd2s1 U4032 ( .DIN1(n562), .DIN2(n456), .Q(n3426) );
  nnd2s1 U4033 ( .DIN1(n3103), .DIN2(n175), .Q(n3428) );
  nnd2s1 U4034 ( .DIN1(n3429), .DIN2(n3430), .Q(\IDinst/n5196 ) );
  nnd2s1 U4035 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][22] ), .Q(n3430) );
  nnd2s1 U4036 ( .DIN1(n597), .DIN2(n459), .Q(n3429) );
  nnd2s1 U4037 ( .DIN1(n3431), .DIN2(n3432), .Q(\IDinst/n5195 ) );
  nnd2s1 U4038 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][22] ), .Q(n3432) );
  nnd2s1 U4039 ( .DIN1(n599), .DIN2(n458), .Q(n3431) );
  nnd2s1 U4040 ( .DIN1(n3433), .DIN2(n3434), .Q(\IDinst/n5194 ) );
  nnd2s1 U4041 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][22] ), .Q(n3434) );
  nnd2s1 U4042 ( .DIN1(n601), .DIN2(n459), .Q(n3433) );
  nnd2s1 U4043 ( .DIN1(n3435), .DIN2(n3436), .Q(\IDinst/n5193 ) );
  nnd2s1 U4044 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][22] ), .Q(n3436) );
  nnd2s1 U4045 ( .DIN1(n603), .DIN2(n458), .Q(n3435) );
  nnd2s1 U4046 ( .DIN1(n3437), .DIN2(n3438), .Q(\IDinst/n5192 ) );
  nnd2s1 U4047 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][22] ), .Q(n3438) );
  nnd2s1 U4048 ( .DIN1(n589), .DIN2(n459), .Q(n3437) );
  nnd2s1 U4049 ( .DIN1(n3439), .DIN2(n3440), .Q(\IDinst/n5191 ) );
  nnd2s1 U4050 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][22] ), .Q(n3440) );
  nnd2s1 U4051 ( .DIN1(n591), .DIN2(n458), .Q(n3439) );
  nnd2s1 U4052 ( .DIN1(n3441), .DIN2(n3442), .Q(\IDinst/n5190 ) );
  nnd2s1 U4053 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][22] ), .Q(n3442) );
  nnd2s1 U4054 ( .DIN1(n593), .DIN2(n459), .Q(n3441) );
  nnd2s1 U4055 ( .DIN1(n3443), .DIN2(n3444), .Q(\IDinst/n5189 ) );
  nnd2s1 U4056 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][22] ), .Q(n3444) );
  nnd2s1 U4057 ( .DIN1(n595), .DIN2(n458), .Q(n3443) );
  nnd2s1 U4058 ( .DIN1(n3445), .DIN2(n3446), .Q(\IDinst/n5188 ) );
  nnd2s1 U4059 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][22] ), .Q(n3446) );
  nnd2s1 U4060 ( .DIN1(n613), .DIN2(n459), .Q(n3445) );
  nnd2s1 U4061 ( .DIN1(n3447), .DIN2(n3448), .Q(\IDinst/n5187 ) );
  nnd2s1 U4062 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][22] ), .Q(n3448) );
  nnd2s1 U4063 ( .DIN1(n615), .DIN2(n458), .Q(n3447) );
  nnd2s1 U4064 ( .DIN1(n3449), .DIN2(n3450), .Q(\IDinst/n5186 ) );
  nnd2s1 U4065 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][22] ), .Q(n3450) );
  nnd2s1 U4066 ( .DIN1(n617), .DIN2(n459), .Q(n3449) );
  nnd2s1 U4067 ( .DIN1(n3451), .DIN2(n3452), .Q(\IDinst/n5185 ) );
  nnd2s1 U4068 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][22] ), .Q(n3452) );
  nnd2s1 U4069 ( .DIN1(n619), .DIN2(n458), .Q(n3451) );
  nnd2s1 U4070 ( .DIN1(n3453), .DIN2(n3454), .Q(\IDinst/n5184 ) );
  nnd2s1 U4071 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][22] ), .Q(n3454) );
  nnd2s1 U4072 ( .DIN1(n605), .DIN2(n459), .Q(n3453) );
  nnd2s1 U4073 ( .DIN1(n3455), .DIN2(n3456), .Q(\IDinst/n5183 ) );
  nnd2s1 U4074 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][22] ), .Q(n3456) );
  nnd2s1 U4075 ( .DIN1(n607), .DIN2(n458), .Q(n3455) );
  nnd2s1 U4076 ( .DIN1(n3457), .DIN2(n3458), .Q(\IDinst/n5182 ) );
  nnd2s1 U4077 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][22] ), .Q(n3458) );
  nnd2s1 U4078 ( .DIN1(n609), .DIN2(n459), .Q(n3457) );
  nnd2s1 U4079 ( .DIN1(n3459), .DIN2(n3460), .Q(\IDinst/n5181 ) );
  nnd2s1 U4080 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][22] ), .Q(n3460) );
  nnd2s1 U4081 ( .DIN1(n611), .DIN2(n458), .Q(n3459) );
  nnd2s1 U4082 ( .DIN1(n3461), .DIN2(n3462), .Q(\IDinst/n5180 ) );
  nnd2s1 U4083 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][22] ), .Q(n3462) );
  nnd2s1 U4084 ( .DIN1(n581), .DIN2(n459), .Q(n3461) );
  nnd2s1 U4085 ( .DIN1(n3463), .DIN2(n3464), .Q(\IDinst/n5179 ) );
  nnd2s1 U4086 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][22] ), .Q(n3464) );
  nnd2s1 U4087 ( .DIN1(n583), .DIN2(n458), .Q(n3463) );
  nnd2s1 U4088 ( .DIN1(n3465), .DIN2(n3466), .Q(\IDinst/n5178 ) );
  nnd2s1 U4089 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][22] ), .Q(n3466) );
  nnd2s1 U4090 ( .DIN1(n585), .DIN2(n459), .Q(n3465) );
  nnd2s1 U4091 ( .DIN1(n3467), .DIN2(n3468), .Q(\IDinst/n5177 ) );
  nnd2s1 U4092 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][22] ), .Q(n3468) );
  nnd2s1 U4093 ( .DIN1(n587), .DIN2(n458), .Q(n3467) );
  nnd2s1 U4094 ( .DIN1(n3469), .DIN2(n3470), .Q(\IDinst/n5176 ) );
  nnd2s1 U4095 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][22] ), .Q(n3470) );
  nnd2s1 U4096 ( .DIN1(n573), .DIN2(n459), .Q(n3469) );
  nnd2s1 U4097 ( .DIN1(n3471), .DIN2(n3472), .Q(\IDinst/n5175 ) );
  nnd2s1 U4098 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][22] ), .Q(n3472) );
  nnd2s1 U4099 ( .DIN1(n575), .DIN2(n458), .Q(n3471) );
  nnd2s1 U4100 ( .DIN1(n3473), .DIN2(n3474), .Q(\IDinst/n5174 ) );
  nnd2s1 U4101 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][22] ), .Q(n3474) );
  nnd2s1 U4102 ( .DIN1(n577), .DIN2(n459), .Q(n3473) );
  nnd2s1 U4103 ( .DIN1(n3475), .DIN2(n3476), .Q(\IDinst/n5173 ) );
  nnd2s1 U4104 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][22] ), .Q(n3476) );
  nnd2s1 U4105 ( .DIN1(n579), .DIN2(n458), .Q(n3475) );
  nnd2s1 U4106 ( .DIN1(n3477), .DIN2(n3478), .Q(\IDinst/n5172 ) );
  nnd2s1 U4107 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][22] ), .Q(n3478) );
  nnd2s1 U4108 ( .DIN1(n565), .DIN2(n459), .Q(n3477) );
  nnd2s1 U4109 ( .DIN1(n3479), .DIN2(n3480), .Q(\IDinst/n5171 ) );
  nnd2s1 U4110 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][22] ), .Q(n3480) );
  nnd2s1 U4111 ( .DIN1(n567), .DIN2(n458), .Q(n3479) );
  nnd2s1 U4112 ( .DIN1(n3481), .DIN2(n3482), .Q(\IDinst/n5170 ) );
  nnd2s1 U4113 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][22] ), .Q(n3482) );
  nnd2s1 U4114 ( .DIN1(n569), .DIN2(n459), .Q(n3481) );
  nnd2s1 U4115 ( .DIN1(n3483), .DIN2(n3484), .Q(\IDinst/n5169 ) );
  nnd2s1 U4116 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][22] ), .Q(n3484) );
  nnd2s1 U4117 ( .DIN1(n571), .DIN2(n458), .Q(n3483) );
  nnd2s1 U4118 ( .DIN1(n3485), .DIN2(n3486), .Q(\IDinst/n5168 ) );
  nnd2s1 U4119 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][22] ), .Q(n3486) );
  nnd2s1 U4120 ( .DIN1(n557), .DIN2(n459), .Q(n3485) );
  nnd2s1 U4121 ( .DIN1(n3487), .DIN2(n3488), .Q(\IDinst/n5167 ) );
  nnd2s1 U4122 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][22] ), .Q(n3488) );
  nnd2s1 U4123 ( .DIN1(n559), .DIN2(n458), .Q(n3487) );
  nnd2s1 U4124 ( .DIN1(n3489), .DIN2(n3490), .Q(\IDinst/n5166 ) );
  nnd2s1 U4125 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][22] ), .Q(n3490) );
  nnd2s1 U4126 ( .DIN1(n561), .DIN2(n459), .Q(n3489) );
  nnd2s1 U4127 ( .DIN1(n3491), .DIN2(n3492), .Q(\IDinst/n5165 ) );
  nnd2s1 U4128 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][22] ), .Q(n3492) );
  nnd2s1 U4129 ( .DIN1(n563), .DIN2(n458), .Q(n3491) );
  nnd2s1 U4130 ( .DIN1(n3103), .DIN2(n173), .Q(n3493) );
  nnd2s1 U4131 ( .DIN1(n3494), .DIN2(n3495), .Q(\IDinst/n5164 ) );
  nnd2s1 U4132 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][23] ), .Q(n3495) );
  nnd2s1 U4133 ( .DIN1(n596), .DIN2(n689), .Q(n3494) );
  nnd2s1 U4134 ( .DIN1(n3497), .DIN2(n3498), .Q(\IDinst/n5163 ) );
  nnd2s1 U4135 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][23] ), .Q(n3498) );
  nnd2s1 U4136 ( .DIN1(n598), .DIN2(n689), .Q(n3497) );
  nnd2s1 U4137 ( .DIN1(n3499), .DIN2(n3500), .Q(\IDinst/n5162 ) );
  nnd2s1 U4138 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][23] ), .Q(n3500) );
  nnd2s1 U4139 ( .DIN1(n600), .DIN2(n689), .Q(n3499) );
  nnd2s1 U4140 ( .DIN1(n3501), .DIN2(n3502), .Q(\IDinst/n5161 ) );
  nnd2s1 U4141 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][23] ), .Q(n3502) );
  nnd2s1 U4142 ( .DIN1(n602), .DIN2(n689), .Q(n3501) );
  nnd2s1 U4143 ( .DIN1(n3503), .DIN2(n3504), .Q(\IDinst/n5160 ) );
  nnd2s1 U4144 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][23] ), .Q(n3504) );
  nnd2s1 U4145 ( .DIN1(n588), .DIN2(n689), .Q(n3503) );
  nnd2s1 U4146 ( .DIN1(n3505), .DIN2(n3506), .Q(\IDinst/n5159 ) );
  nnd2s1 U4147 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][23] ), .Q(n3506) );
  nnd2s1 U4148 ( .DIN1(n590), .DIN2(n689), .Q(n3505) );
  nnd2s1 U4149 ( .DIN1(n3507), .DIN2(n3508), .Q(\IDinst/n5158 ) );
  nnd2s1 U4150 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][23] ), .Q(n3508) );
  nnd2s1 U4151 ( .DIN1(n592), .DIN2(n689), .Q(n3507) );
  nnd2s1 U4152 ( .DIN1(n3509), .DIN2(n3510), .Q(\IDinst/n5157 ) );
  nnd2s1 U4153 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][23] ), .Q(n3510) );
  nnd2s1 U4154 ( .DIN1(n594), .DIN2(n689), .Q(n3509) );
  nnd2s1 U4155 ( .DIN1(n3511), .DIN2(n3512), .Q(\IDinst/n5156 ) );
  nnd2s1 U4156 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][23] ), .Q(n3512) );
  nnd2s1 U4157 ( .DIN1(n612), .DIN2(n689), .Q(n3511) );
  nnd2s1 U4158 ( .DIN1(n3513), .DIN2(n3514), .Q(\IDinst/n5155 ) );
  nnd2s1 U4159 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][23] ), .Q(n3514) );
  nnd2s1 U4160 ( .DIN1(n614), .DIN2(n689), .Q(n3513) );
  nnd2s1 U4161 ( .DIN1(n3515), .DIN2(n3516), .Q(\IDinst/n5154 ) );
  nnd2s1 U4162 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][23] ), .Q(n3516) );
  nnd2s1 U4163 ( .DIN1(n616), .DIN2(n689), .Q(n3515) );
  nnd2s1 U4164 ( .DIN1(n3517), .DIN2(n3518), .Q(\IDinst/n5153 ) );
  nnd2s1 U4165 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][23] ), .Q(n3518) );
  nnd2s1 U4166 ( .DIN1(n618), .DIN2(n689), .Q(n3517) );
  nnd2s1 U4167 ( .DIN1(n3519), .DIN2(n3520), .Q(\IDinst/n5152 ) );
  nnd2s1 U4168 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][23] ), .Q(n3520) );
  nnd2s1 U4169 ( .DIN1(n604), .DIN2(n689), .Q(n3519) );
  nnd2s1 U4170 ( .DIN1(n3521), .DIN2(n3522), .Q(\IDinst/n5151 ) );
  nnd2s1 U4171 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][23] ), .Q(n3522) );
  nnd2s1 U4172 ( .DIN1(n606), .DIN2(n3496), .Q(n3521) );
  nnd2s1 U4173 ( .DIN1(n3523), .DIN2(n3524), .Q(\IDinst/n5150 ) );
  nnd2s1 U4174 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][23] ), .Q(n3524) );
  nnd2s1 U4175 ( .DIN1(n608), .DIN2(n3496), .Q(n3523) );
  nnd2s1 U4176 ( .DIN1(n3525), .DIN2(n3526), .Q(\IDinst/n5149 ) );
  nnd2s1 U4177 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][23] ), .Q(n3526) );
  nnd2s1 U4178 ( .DIN1(n610), .DIN2(n3496), .Q(n3525) );
  nnd2s1 U4179 ( .DIN1(n3527), .DIN2(n3528), .Q(\IDinst/n5148 ) );
  nnd2s1 U4180 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][23] ), .Q(n3528) );
  nnd2s1 U4181 ( .DIN1(n580), .DIN2(n3496), .Q(n3527) );
  nnd2s1 U4182 ( .DIN1(n3529), .DIN2(n3530), .Q(\IDinst/n5147 ) );
  nnd2s1 U4183 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][23] ), .Q(n3530) );
  nnd2s1 U4184 ( .DIN1(n582), .DIN2(n3496), .Q(n3529) );
  nnd2s1 U4185 ( .DIN1(n3531), .DIN2(n3532), .Q(\IDinst/n5146 ) );
  nnd2s1 U4186 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][23] ), .Q(n3532) );
  nnd2s1 U4187 ( .DIN1(n584), .DIN2(n3496), .Q(n3531) );
  nnd2s1 U4188 ( .DIN1(n3533), .DIN2(n3534), .Q(\IDinst/n5145 ) );
  nnd2s1 U4189 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][23] ), .Q(n3534) );
  nnd2s1 U4190 ( .DIN1(n586), .DIN2(n3496), .Q(n3533) );
  nnd2s1 U4191 ( .DIN1(n3535), .DIN2(n3536), .Q(\IDinst/n5144 ) );
  nnd2s1 U4192 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][23] ), .Q(n3536) );
  nnd2s1 U4193 ( .DIN1(n572), .DIN2(n3496), .Q(n3535) );
  nnd2s1 U4194 ( .DIN1(n3537), .DIN2(n3538), .Q(\IDinst/n5143 ) );
  nnd2s1 U4195 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][23] ), .Q(n3538) );
  nnd2s1 U4196 ( .DIN1(n574), .DIN2(n3496), .Q(n3537) );
  nnd2s1 U4197 ( .DIN1(n3539), .DIN2(n3540), .Q(\IDinst/n5142 ) );
  nnd2s1 U4198 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][23] ), .Q(n3540) );
  nnd2s1 U4199 ( .DIN1(n576), .DIN2(n3496), .Q(n3539) );
  nnd2s1 U4200 ( .DIN1(n3541), .DIN2(n3542), .Q(\IDinst/n5141 ) );
  nnd2s1 U4201 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][23] ), .Q(n3542) );
  nnd2s1 U4202 ( .DIN1(n578), .DIN2(n3496), .Q(n3541) );
  nnd2s1 U4203 ( .DIN1(n3543), .DIN2(n3544), .Q(\IDinst/n5140 ) );
  nnd2s1 U4204 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][23] ), .Q(n3544) );
  nnd2s1 U4205 ( .DIN1(n564), .DIN2(n3496), .Q(n3543) );
  nnd2s1 U4206 ( .DIN1(n3545), .DIN2(n3546), .Q(\IDinst/n5139 ) );
  nnd2s1 U4207 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][23] ), .Q(n3546) );
  nnd2s1 U4208 ( .DIN1(n566), .DIN2(n3496), .Q(n3545) );
  nnd2s1 U4209 ( .DIN1(n3547), .DIN2(n3548), .Q(\IDinst/n5138 ) );
  nnd2s1 U4210 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][23] ), .Q(n3548) );
  nnd2s1 U4211 ( .DIN1(n568), .DIN2(n3496), .Q(n3547) );
  nnd2s1 U4212 ( .DIN1(n3549), .DIN2(n3550), .Q(\IDinst/n5137 ) );
  nnd2s1 U4213 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][23] ), .Q(n3550) );
  nnd2s1 U4214 ( .DIN1(n570), .DIN2(n3496), .Q(n3549) );
  nnd2s1 U4215 ( .DIN1(n3551), .DIN2(n3552), .Q(\IDinst/n5136 ) );
  nnd2s1 U4216 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][23] ), .Q(n3552) );
  nnd2s1 U4217 ( .DIN1(n556), .DIN2(n3496), .Q(n3551) );
  nnd2s1 U4218 ( .DIN1(n3553), .DIN2(n3554), .Q(\IDinst/n5135 ) );
  nnd2s1 U4219 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][23] ), .Q(n3554) );
  nnd2s1 U4220 ( .DIN1(n558), .DIN2(n3496), .Q(n3553) );
  nnd2s1 U4221 ( .DIN1(n3555), .DIN2(n3556), .Q(\IDinst/n5134 ) );
  nnd2s1 U4222 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][23] ), .Q(n3556) );
  nnd2s1 U4223 ( .DIN1(n560), .DIN2(n3496), .Q(n3555) );
  nnd2s1 U4224 ( .DIN1(n3557), .DIN2(n3558), .Q(\IDinst/n5133 ) );
  nnd2s1 U4225 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][23] ), .Q(n3558) );
  nnd2s1 U4226 ( .DIN1(n562), .DIN2(n3496), .Q(n3557) );
  nnd2s1 U4227 ( .DIN1(n3035), .DIN2(n3559), .Q(n3496) );
  nnd2s1 U4228 ( .DIN1(n3103), .DIN2(n171), .Q(n3559) );
  nnd2s1 U4229 ( .DIN1(n3560), .DIN2(n3561), .Q(\IDinst/n5132 ) );
  nnd2s1 U4230 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][24] ), .Q(n3561) );
  nnd2s1 U4231 ( .DIN1(n597), .DIN2(n691), .Q(n3560) );
  nnd2s1 U4232 ( .DIN1(n3563), .DIN2(n3564), .Q(\IDinst/n5131 ) );
  nnd2s1 U4233 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][24] ), .Q(n3564) );
  nnd2s1 U4234 ( .DIN1(n599), .DIN2(n691), .Q(n3563) );
  nnd2s1 U4235 ( .DIN1(n3565), .DIN2(n3566), .Q(\IDinst/n5130 ) );
  nnd2s1 U4236 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][24] ), .Q(n3566) );
  nnd2s1 U4237 ( .DIN1(n601), .DIN2(n691), .Q(n3565) );
  nnd2s1 U4238 ( .DIN1(n3567), .DIN2(n3568), .Q(\IDinst/n5129 ) );
  nnd2s1 U4239 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][24] ), .Q(n3568) );
  nnd2s1 U4240 ( .DIN1(n603), .DIN2(n691), .Q(n3567) );
  nnd2s1 U4241 ( .DIN1(n3569), .DIN2(n3570), .Q(\IDinst/n5128 ) );
  nnd2s1 U4242 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][24] ), .Q(n3570) );
  nnd2s1 U4243 ( .DIN1(n589), .DIN2(n691), .Q(n3569) );
  nnd2s1 U4244 ( .DIN1(n3571), .DIN2(n3572), .Q(\IDinst/n5127 ) );
  nnd2s1 U4245 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][24] ), .Q(n3572) );
  nnd2s1 U4246 ( .DIN1(n591), .DIN2(n691), .Q(n3571) );
  nnd2s1 U4247 ( .DIN1(n3573), .DIN2(n3574), .Q(\IDinst/n5126 ) );
  nnd2s1 U4248 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][24] ), .Q(n3574) );
  nnd2s1 U4249 ( .DIN1(n593), .DIN2(n691), .Q(n3573) );
  nnd2s1 U4250 ( .DIN1(n3575), .DIN2(n3576), .Q(\IDinst/n5125 ) );
  nnd2s1 U4251 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][24] ), .Q(n3576) );
  nnd2s1 U4252 ( .DIN1(n595), .DIN2(n691), .Q(n3575) );
  nnd2s1 U4253 ( .DIN1(n3577), .DIN2(n3578), .Q(\IDinst/n5124 ) );
  nnd2s1 U4254 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][24] ), .Q(n3578) );
  nnd2s1 U4255 ( .DIN1(n613), .DIN2(n691), .Q(n3577) );
  nnd2s1 U4256 ( .DIN1(n3579), .DIN2(n3580), .Q(\IDinst/n5123 ) );
  nnd2s1 U4257 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][24] ), .Q(n3580) );
  nnd2s1 U4258 ( .DIN1(n615), .DIN2(n691), .Q(n3579) );
  nnd2s1 U4259 ( .DIN1(n3581), .DIN2(n3582), .Q(\IDinst/n5122 ) );
  nnd2s1 U4260 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][24] ), .Q(n3582) );
  nnd2s1 U4261 ( .DIN1(n617), .DIN2(n691), .Q(n3581) );
  nnd2s1 U4262 ( .DIN1(n3583), .DIN2(n3584), .Q(\IDinst/n5121 ) );
  nnd2s1 U4263 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][24] ), .Q(n3584) );
  nnd2s1 U4264 ( .DIN1(n619), .DIN2(n691), .Q(n3583) );
  nnd2s1 U4265 ( .DIN1(n3585), .DIN2(n3586), .Q(\IDinst/n5120 ) );
  nnd2s1 U4266 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][24] ), .Q(n3586) );
  nnd2s1 U4267 ( .DIN1(n605), .DIN2(n691), .Q(n3585) );
  nnd2s1 U4268 ( .DIN1(n3587), .DIN2(n3588), .Q(\IDinst/n5119 ) );
  nnd2s1 U4269 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][24] ), .Q(n3588) );
  nnd2s1 U4270 ( .DIN1(n607), .DIN2(n3562), .Q(n3587) );
  nnd2s1 U4271 ( .DIN1(n3589), .DIN2(n3590), .Q(\IDinst/n5118 ) );
  nnd2s1 U4272 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][24] ), .Q(n3590) );
  nnd2s1 U4273 ( .DIN1(n609), .DIN2(n3562), .Q(n3589) );
  nnd2s1 U4274 ( .DIN1(n3591), .DIN2(n3592), .Q(\IDinst/n5117 ) );
  nnd2s1 U4275 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][24] ), .Q(n3592) );
  nnd2s1 U4276 ( .DIN1(n611), .DIN2(n3562), .Q(n3591) );
  nnd2s1 U4277 ( .DIN1(n3593), .DIN2(n3594), .Q(\IDinst/n5116 ) );
  nnd2s1 U4278 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][24] ), .Q(n3594) );
  nnd2s1 U4279 ( .DIN1(n581), .DIN2(n3562), .Q(n3593) );
  nnd2s1 U4280 ( .DIN1(n3595), .DIN2(n3596), .Q(\IDinst/n5115 ) );
  nnd2s1 U4281 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][24] ), .Q(n3596) );
  nnd2s1 U4282 ( .DIN1(n583), .DIN2(n3562), .Q(n3595) );
  nnd2s1 U4283 ( .DIN1(n3597), .DIN2(n3598), .Q(\IDinst/n5114 ) );
  nnd2s1 U4284 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][24] ), .Q(n3598) );
  nnd2s1 U4285 ( .DIN1(n585), .DIN2(n3562), .Q(n3597) );
  nnd2s1 U4286 ( .DIN1(n3599), .DIN2(n3600), .Q(\IDinst/n5113 ) );
  nnd2s1 U4287 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][24] ), .Q(n3600) );
  nnd2s1 U4288 ( .DIN1(n587), .DIN2(n3562), .Q(n3599) );
  nnd2s1 U4289 ( .DIN1(n3601), .DIN2(n3602), .Q(\IDinst/n5112 ) );
  nnd2s1 U4290 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][24] ), .Q(n3602) );
  nnd2s1 U4291 ( .DIN1(n573), .DIN2(n3562), .Q(n3601) );
  nnd2s1 U4292 ( .DIN1(n3603), .DIN2(n3604), .Q(\IDinst/n5111 ) );
  nnd2s1 U4293 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][24] ), .Q(n3604) );
  nnd2s1 U4294 ( .DIN1(n575), .DIN2(n3562), .Q(n3603) );
  nnd2s1 U4295 ( .DIN1(n3605), .DIN2(n3606), .Q(\IDinst/n5110 ) );
  nnd2s1 U4296 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][24] ), .Q(n3606) );
  nnd2s1 U4297 ( .DIN1(n577), .DIN2(n3562), .Q(n3605) );
  nnd2s1 U4298 ( .DIN1(n3607), .DIN2(n3608), .Q(\IDinst/n5109 ) );
  nnd2s1 U4299 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][24] ), .Q(n3608) );
  nnd2s1 U4300 ( .DIN1(n579), .DIN2(n3562), .Q(n3607) );
  nnd2s1 U4301 ( .DIN1(n3609), .DIN2(n3610), .Q(\IDinst/n5108 ) );
  nnd2s1 U4302 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][24] ), .Q(n3610) );
  nnd2s1 U4303 ( .DIN1(n565), .DIN2(n3562), .Q(n3609) );
  nnd2s1 U4304 ( .DIN1(n3611), .DIN2(n3612), .Q(\IDinst/n5107 ) );
  nnd2s1 U4305 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][24] ), .Q(n3612) );
  nnd2s1 U4306 ( .DIN1(n567), .DIN2(n3562), .Q(n3611) );
  nnd2s1 U4307 ( .DIN1(n3613), .DIN2(n3614), .Q(\IDinst/n5106 ) );
  nnd2s1 U4308 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][24] ), .Q(n3614) );
  nnd2s1 U4309 ( .DIN1(n569), .DIN2(n3562), .Q(n3613) );
  nnd2s1 U4310 ( .DIN1(n3615), .DIN2(n3616), .Q(\IDinst/n5105 ) );
  nnd2s1 U4311 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][24] ), .Q(n3616) );
  nnd2s1 U4312 ( .DIN1(n571), .DIN2(n3562), .Q(n3615) );
  nnd2s1 U4313 ( .DIN1(n3617), .DIN2(n3618), .Q(\IDinst/n5104 ) );
  nnd2s1 U4314 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][24] ), .Q(n3618) );
  nnd2s1 U4315 ( .DIN1(n557), .DIN2(n3562), .Q(n3617) );
  nnd2s1 U4316 ( .DIN1(n3619), .DIN2(n3620), .Q(\IDinst/n5103 ) );
  nnd2s1 U4317 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][24] ), .Q(n3620) );
  nnd2s1 U4318 ( .DIN1(n559), .DIN2(n3562), .Q(n3619) );
  nnd2s1 U4319 ( .DIN1(n3621), .DIN2(n3622), .Q(\IDinst/n5102 ) );
  nnd2s1 U4320 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][24] ), .Q(n3622) );
  nnd2s1 U4321 ( .DIN1(n561), .DIN2(n3562), .Q(n3621) );
  nnd2s1 U4322 ( .DIN1(n3623), .DIN2(n3624), .Q(\IDinst/n5101 ) );
  nnd2s1 U4323 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][24] ), .Q(n3624) );
  nnd2s1 U4324 ( .DIN1(n563), .DIN2(n3562), .Q(n3623) );
  nnd2s1 U4325 ( .DIN1(n3035), .DIN2(n3625), .Q(n3562) );
  nnd2s1 U4326 ( .DIN1(n3103), .DIN2(n169), .Q(n3625) );
  nnd2s1 U4327 ( .DIN1(n3626), .DIN2(n3627), .Q(\IDinst/n5100 ) );
  nnd2s1 U4328 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][25] ), .Q(n3627) );
  nnd2s1 U4329 ( .DIN1(n596), .DIN2(n695), .Q(n3626) );
  nnd2s1 U4330 ( .DIN1(n3629), .DIN2(n3630), .Q(\IDinst/n5099 ) );
  nnd2s1 U4331 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][25] ), .Q(n3630) );
  nnd2s1 U4332 ( .DIN1(n598), .DIN2(n695), .Q(n3629) );
  nnd2s1 U4333 ( .DIN1(n3631), .DIN2(n3632), .Q(\IDinst/n5098 ) );
  nnd2s1 U4334 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][25] ), .Q(n3632) );
  nnd2s1 U4335 ( .DIN1(n600), .DIN2(n695), .Q(n3631) );
  nnd2s1 U4336 ( .DIN1(n3633), .DIN2(n3634), .Q(\IDinst/n5097 ) );
  nnd2s1 U4337 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][25] ), .Q(n3634) );
  nnd2s1 U4338 ( .DIN1(n602), .DIN2(n695), .Q(n3633) );
  nnd2s1 U4339 ( .DIN1(n3635), .DIN2(n3636), .Q(\IDinst/n5096 ) );
  nnd2s1 U4340 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][25] ), .Q(n3636) );
  nnd2s1 U4341 ( .DIN1(n588), .DIN2(n695), .Q(n3635) );
  nnd2s1 U4342 ( .DIN1(n3637), .DIN2(n3638), .Q(\IDinst/n5095 ) );
  nnd2s1 U4343 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][25] ), .Q(n3638) );
  nnd2s1 U4344 ( .DIN1(n590), .DIN2(n695), .Q(n3637) );
  nnd2s1 U4345 ( .DIN1(n3639), .DIN2(n3640), .Q(\IDinst/n5094 ) );
  nnd2s1 U4346 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][25] ), .Q(n3640) );
  nnd2s1 U4347 ( .DIN1(n592), .DIN2(n695), .Q(n3639) );
  nnd2s1 U4348 ( .DIN1(n3641), .DIN2(n3642), .Q(\IDinst/n5093 ) );
  nnd2s1 U4349 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][25] ), .Q(n3642) );
  nnd2s1 U4350 ( .DIN1(n594), .DIN2(n695), .Q(n3641) );
  nnd2s1 U4351 ( .DIN1(n3643), .DIN2(n3644), .Q(\IDinst/n5092 ) );
  nnd2s1 U4352 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][25] ), .Q(n3644) );
  nnd2s1 U4353 ( .DIN1(n612), .DIN2(n695), .Q(n3643) );
  nnd2s1 U4354 ( .DIN1(n3645), .DIN2(n3646), .Q(\IDinst/n5091 ) );
  nnd2s1 U4355 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][25] ), .Q(n3646) );
  nnd2s1 U4356 ( .DIN1(n614), .DIN2(n695), .Q(n3645) );
  nnd2s1 U4357 ( .DIN1(n3647), .DIN2(n3648), .Q(\IDinst/n5090 ) );
  nnd2s1 U4358 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][25] ), .Q(n3648) );
  nnd2s1 U4359 ( .DIN1(n616), .DIN2(n695), .Q(n3647) );
  nnd2s1 U4360 ( .DIN1(n3649), .DIN2(n3650), .Q(\IDinst/n5089 ) );
  nnd2s1 U4361 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][25] ), .Q(n3650) );
  nnd2s1 U4362 ( .DIN1(n618), .DIN2(n695), .Q(n3649) );
  nnd2s1 U4363 ( .DIN1(n3651), .DIN2(n3652), .Q(\IDinst/n5088 ) );
  nnd2s1 U4364 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][25] ), .Q(n3652) );
  nnd2s1 U4365 ( .DIN1(n604), .DIN2(n695), .Q(n3651) );
  nnd2s1 U4366 ( .DIN1(n3653), .DIN2(n3654), .Q(\IDinst/n5087 ) );
  nnd2s1 U4367 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][25] ), .Q(n3654) );
  nnd2s1 U4368 ( .DIN1(n606), .DIN2(n3628), .Q(n3653) );
  nnd2s1 U4369 ( .DIN1(n3655), .DIN2(n3656), .Q(\IDinst/n5086 ) );
  nnd2s1 U4370 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][25] ), .Q(n3656) );
  nnd2s1 U4371 ( .DIN1(n608), .DIN2(n3628), .Q(n3655) );
  nnd2s1 U4372 ( .DIN1(n3657), .DIN2(n3658), .Q(\IDinst/n5085 ) );
  nnd2s1 U4373 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][25] ), .Q(n3658) );
  nnd2s1 U4374 ( .DIN1(n610), .DIN2(n3628), .Q(n3657) );
  nnd2s1 U4375 ( .DIN1(n3659), .DIN2(n3660), .Q(\IDinst/n5084 ) );
  nnd2s1 U4376 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][25] ), .Q(n3660) );
  nnd2s1 U4377 ( .DIN1(n580), .DIN2(n3628), .Q(n3659) );
  nnd2s1 U4378 ( .DIN1(n3661), .DIN2(n3662), .Q(\IDinst/n5083 ) );
  nnd2s1 U4379 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][25] ), .Q(n3662) );
  nnd2s1 U4380 ( .DIN1(n582), .DIN2(n3628), .Q(n3661) );
  nnd2s1 U4381 ( .DIN1(n3663), .DIN2(n3664), .Q(\IDinst/n5082 ) );
  nnd2s1 U4382 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][25] ), .Q(n3664) );
  nnd2s1 U4383 ( .DIN1(n584), .DIN2(n3628), .Q(n3663) );
  nnd2s1 U4384 ( .DIN1(n3665), .DIN2(n3666), .Q(\IDinst/n5081 ) );
  nnd2s1 U4385 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][25] ), .Q(n3666) );
  nnd2s1 U4386 ( .DIN1(n586), .DIN2(n3628), .Q(n3665) );
  nnd2s1 U4387 ( .DIN1(n3667), .DIN2(n3668), .Q(\IDinst/n5080 ) );
  nnd2s1 U4388 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][25] ), .Q(n3668) );
  nnd2s1 U4389 ( .DIN1(n572), .DIN2(n3628), .Q(n3667) );
  nnd2s1 U4390 ( .DIN1(n3669), .DIN2(n3670), .Q(\IDinst/n5079 ) );
  nnd2s1 U4391 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][25] ), .Q(n3670) );
  nnd2s1 U4392 ( .DIN1(n574), .DIN2(n3628), .Q(n3669) );
  nnd2s1 U4393 ( .DIN1(n3671), .DIN2(n3672), .Q(\IDinst/n5078 ) );
  nnd2s1 U4394 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][25] ), .Q(n3672) );
  nnd2s1 U4395 ( .DIN1(n576), .DIN2(n3628), .Q(n3671) );
  nnd2s1 U4396 ( .DIN1(n3673), .DIN2(n3674), .Q(\IDinst/n5077 ) );
  nnd2s1 U4397 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][25] ), .Q(n3674) );
  nnd2s1 U4398 ( .DIN1(n578), .DIN2(n3628), .Q(n3673) );
  nnd2s1 U4399 ( .DIN1(n3675), .DIN2(n3676), .Q(\IDinst/n5076 ) );
  nnd2s1 U4400 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][25] ), .Q(n3676) );
  nnd2s1 U4401 ( .DIN1(n564), .DIN2(n3628), .Q(n3675) );
  nnd2s1 U4402 ( .DIN1(n3677), .DIN2(n3678), .Q(\IDinst/n5075 ) );
  nnd2s1 U4403 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][25] ), .Q(n3678) );
  nnd2s1 U4404 ( .DIN1(n566), .DIN2(n3628), .Q(n3677) );
  nnd2s1 U4405 ( .DIN1(n3679), .DIN2(n3680), .Q(\IDinst/n5074 ) );
  nnd2s1 U4406 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][25] ), .Q(n3680) );
  nnd2s1 U4407 ( .DIN1(n568), .DIN2(n3628), .Q(n3679) );
  nnd2s1 U4408 ( .DIN1(n3681), .DIN2(n3682), .Q(\IDinst/n5073 ) );
  nnd2s1 U4409 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][25] ), .Q(n3682) );
  nnd2s1 U4410 ( .DIN1(n570), .DIN2(n3628), .Q(n3681) );
  nnd2s1 U4411 ( .DIN1(n3683), .DIN2(n3684), .Q(\IDinst/n5072 ) );
  nnd2s1 U4412 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][25] ), .Q(n3684) );
  nnd2s1 U4413 ( .DIN1(n556), .DIN2(n3628), .Q(n3683) );
  nnd2s1 U4414 ( .DIN1(n3685), .DIN2(n3686), .Q(\IDinst/n5071 ) );
  nnd2s1 U4415 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][25] ), .Q(n3686) );
  nnd2s1 U4416 ( .DIN1(n558), .DIN2(n3628), .Q(n3685) );
  nnd2s1 U4417 ( .DIN1(n3687), .DIN2(n3688), .Q(\IDinst/n5070 ) );
  nnd2s1 U4418 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][25] ), .Q(n3688) );
  nnd2s1 U4419 ( .DIN1(n560), .DIN2(n3628), .Q(n3687) );
  nnd2s1 U4420 ( .DIN1(n3689), .DIN2(n3690), .Q(\IDinst/n5069 ) );
  nnd2s1 U4421 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][25] ), .Q(n3690) );
  nnd2s1 U4422 ( .DIN1(n562), .DIN2(n3628), .Q(n3689) );
  nnd2s1 U4423 ( .DIN1(n3035), .DIN2(n3691), .Q(n3628) );
  nnd2s1 U4424 ( .DIN1(n3103), .DIN2(n167), .Q(n3691) );
  nnd2s1 U4425 ( .DIN1(n3692), .DIN2(n3693), .Q(\IDinst/n5068 ) );
  nnd2s1 U4426 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][26] ), .Q(n3693) );
  nnd2s1 U4427 ( .DIN1(n597), .DIN2(n699), .Q(n3692) );
  nnd2s1 U4428 ( .DIN1(n3695), .DIN2(n3696), .Q(\IDinst/n5067 ) );
  nnd2s1 U4429 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][26] ), .Q(n3696) );
  nnd2s1 U4430 ( .DIN1(n599), .DIN2(n699), .Q(n3695) );
  nnd2s1 U4431 ( .DIN1(n3697), .DIN2(n3698), .Q(\IDinst/n5066 ) );
  nnd2s1 U4432 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][26] ), .Q(n3698) );
  nnd2s1 U4433 ( .DIN1(n601), .DIN2(n699), .Q(n3697) );
  nnd2s1 U4434 ( .DIN1(n3699), .DIN2(n3700), .Q(\IDinst/n5065 ) );
  nnd2s1 U4435 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][26] ), .Q(n3700) );
  nnd2s1 U4436 ( .DIN1(n603), .DIN2(n699), .Q(n3699) );
  nnd2s1 U4437 ( .DIN1(n3701), .DIN2(n3702), .Q(\IDinst/n5064 ) );
  nnd2s1 U4438 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][26] ), .Q(n3702) );
  nnd2s1 U4439 ( .DIN1(n589), .DIN2(n699), .Q(n3701) );
  nnd2s1 U4440 ( .DIN1(n3703), .DIN2(n3704), .Q(\IDinst/n5063 ) );
  nnd2s1 U4441 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][26] ), .Q(n3704) );
  nnd2s1 U4442 ( .DIN1(n591), .DIN2(n699), .Q(n3703) );
  nnd2s1 U4443 ( .DIN1(n3705), .DIN2(n3706), .Q(\IDinst/n5062 ) );
  nnd2s1 U4444 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][26] ), .Q(n3706) );
  nnd2s1 U4445 ( .DIN1(n593), .DIN2(n699), .Q(n3705) );
  nnd2s1 U4446 ( .DIN1(n3707), .DIN2(n3708), .Q(\IDinst/n5061 ) );
  nnd2s1 U4447 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][26] ), .Q(n3708) );
  nnd2s1 U4448 ( .DIN1(n595), .DIN2(n699), .Q(n3707) );
  nnd2s1 U4449 ( .DIN1(n3709), .DIN2(n3710), .Q(\IDinst/n5060 ) );
  nnd2s1 U4450 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][26] ), .Q(n3710) );
  nnd2s1 U4451 ( .DIN1(n613), .DIN2(n699), .Q(n3709) );
  nnd2s1 U4452 ( .DIN1(n3711), .DIN2(n3712), .Q(\IDinst/n5059 ) );
  nnd2s1 U4453 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][26] ), .Q(n3712) );
  nnd2s1 U4454 ( .DIN1(n615), .DIN2(n699), .Q(n3711) );
  nnd2s1 U4455 ( .DIN1(n3713), .DIN2(n3714), .Q(\IDinst/n5058 ) );
  nnd2s1 U4456 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][26] ), .Q(n3714) );
  nnd2s1 U4457 ( .DIN1(n617), .DIN2(n699), .Q(n3713) );
  nnd2s1 U4458 ( .DIN1(n3715), .DIN2(n3716), .Q(\IDinst/n5057 ) );
  nnd2s1 U4459 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][26] ), .Q(n3716) );
  nnd2s1 U4460 ( .DIN1(n619), .DIN2(n699), .Q(n3715) );
  nnd2s1 U4461 ( .DIN1(n3717), .DIN2(n3718), .Q(\IDinst/n5056 ) );
  nnd2s1 U4462 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][26] ), .Q(n3718) );
  nnd2s1 U4463 ( .DIN1(n605), .DIN2(n699), .Q(n3717) );
  nnd2s1 U4464 ( .DIN1(n3719), .DIN2(n3720), .Q(\IDinst/n5055 ) );
  nnd2s1 U4465 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][26] ), .Q(n3720) );
  nnd2s1 U4466 ( .DIN1(n607), .DIN2(n3694), .Q(n3719) );
  nnd2s1 U4467 ( .DIN1(n3721), .DIN2(n3722), .Q(\IDinst/n5054 ) );
  nnd2s1 U4468 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][26] ), .Q(n3722) );
  nnd2s1 U4469 ( .DIN1(n609), .DIN2(n3694), .Q(n3721) );
  nnd2s1 U4470 ( .DIN1(n3723), .DIN2(n3724), .Q(\IDinst/n5053 ) );
  nnd2s1 U4471 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][26] ), .Q(n3724) );
  nnd2s1 U4472 ( .DIN1(n611), .DIN2(n3694), .Q(n3723) );
  nnd2s1 U4473 ( .DIN1(n3725), .DIN2(n3726), .Q(\IDinst/n5052 ) );
  nnd2s1 U4474 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][26] ), .Q(n3726) );
  nnd2s1 U4475 ( .DIN1(n581), .DIN2(n3694), .Q(n3725) );
  nnd2s1 U4476 ( .DIN1(n3727), .DIN2(n3728), .Q(\IDinst/n5051 ) );
  nnd2s1 U4477 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][26] ), .Q(n3728) );
  nnd2s1 U4478 ( .DIN1(n583), .DIN2(n3694), .Q(n3727) );
  nnd2s1 U4479 ( .DIN1(n3729), .DIN2(n3730), .Q(\IDinst/n5050 ) );
  nnd2s1 U4480 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][26] ), .Q(n3730) );
  nnd2s1 U4481 ( .DIN1(n585), .DIN2(n3694), .Q(n3729) );
  nnd2s1 U4482 ( .DIN1(n3731), .DIN2(n3732), .Q(\IDinst/n5049 ) );
  nnd2s1 U4483 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][26] ), .Q(n3732) );
  nnd2s1 U4484 ( .DIN1(n587), .DIN2(n3694), .Q(n3731) );
  nnd2s1 U4485 ( .DIN1(n3733), .DIN2(n3734), .Q(\IDinst/n5048 ) );
  nnd2s1 U4486 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][26] ), .Q(n3734) );
  nnd2s1 U4487 ( .DIN1(n573), .DIN2(n3694), .Q(n3733) );
  nnd2s1 U4488 ( .DIN1(n3735), .DIN2(n3736), .Q(\IDinst/n5047 ) );
  nnd2s1 U4489 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][26] ), .Q(n3736) );
  nnd2s1 U4490 ( .DIN1(n575), .DIN2(n3694), .Q(n3735) );
  nnd2s1 U4491 ( .DIN1(n3737), .DIN2(n3738), .Q(\IDinst/n5046 ) );
  nnd2s1 U4492 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][26] ), .Q(n3738) );
  nnd2s1 U4493 ( .DIN1(n577), .DIN2(n3694), .Q(n3737) );
  nnd2s1 U4494 ( .DIN1(n3739), .DIN2(n3740), .Q(\IDinst/n5045 ) );
  nnd2s1 U4495 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][26] ), .Q(n3740) );
  nnd2s1 U4496 ( .DIN1(n579), .DIN2(n3694), .Q(n3739) );
  nnd2s1 U4497 ( .DIN1(n3741), .DIN2(n3742), .Q(\IDinst/n5044 ) );
  nnd2s1 U4498 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][26] ), .Q(n3742) );
  nnd2s1 U4499 ( .DIN1(n565), .DIN2(n3694), .Q(n3741) );
  nnd2s1 U4500 ( .DIN1(n3743), .DIN2(n3744), .Q(\IDinst/n5043 ) );
  nnd2s1 U4501 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][26] ), .Q(n3744) );
  nnd2s1 U4502 ( .DIN1(n567), .DIN2(n3694), .Q(n3743) );
  nnd2s1 U4503 ( .DIN1(n3745), .DIN2(n3746), .Q(\IDinst/n5042 ) );
  nnd2s1 U4504 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][26] ), .Q(n3746) );
  nnd2s1 U4505 ( .DIN1(n569), .DIN2(n3694), .Q(n3745) );
  nnd2s1 U4506 ( .DIN1(n3747), .DIN2(n3748), .Q(\IDinst/n5041 ) );
  nnd2s1 U4507 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][26] ), .Q(n3748) );
  nnd2s1 U4508 ( .DIN1(n571), .DIN2(n3694), .Q(n3747) );
  nnd2s1 U4509 ( .DIN1(n3749), .DIN2(n3750), .Q(\IDinst/n5040 ) );
  nnd2s1 U4510 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][26] ), .Q(n3750) );
  nnd2s1 U4511 ( .DIN1(n557), .DIN2(n3694), .Q(n3749) );
  nnd2s1 U4512 ( .DIN1(n3751), .DIN2(n3752), .Q(\IDinst/n5039 ) );
  nnd2s1 U4513 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][26] ), .Q(n3752) );
  nnd2s1 U4514 ( .DIN1(n559), .DIN2(n3694), .Q(n3751) );
  nnd2s1 U4515 ( .DIN1(n3753), .DIN2(n3754), .Q(\IDinst/n5038 ) );
  nnd2s1 U4516 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][26] ), .Q(n3754) );
  nnd2s1 U4517 ( .DIN1(n561), .DIN2(n3694), .Q(n3753) );
  nnd2s1 U4518 ( .DIN1(n3755), .DIN2(n3756), .Q(\IDinst/n5037 ) );
  nnd2s1 U4519 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][26] ), .Q(n3756) );
  nnd2s1 U4520 ( .DIN1(n563), .DIN2(n3694), .Q(n3755) );
  nnd2s1 U4521 ( .DIN1(n3035), .DIN2(n3757), .Q(n3694) );
  nnd2s1 U4522 ( .DIN1(n3103), .DIN2(n165), .Q(n3757) );
  nnd2s1 U4523 ( .DIN1(n3758), .DIN2(n3759), .Q(\IDinst/n5036 ) );
  nnd2s1 U4524 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][27] ), .Q(n3759) );
  nnd2s1 U4525 ( .DIN1(n596), .DIN2(n704), .Q(n3758) );
  nnd2s1 U4526 ( .DIN1(n3761), .DIN2(n3762), .Q(\IDinst/n5035 ) );
  nnd2s1 U4527 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][27] ), .Q(n3762) );
  nnd2s1 U4528 ( .DIN1(n598), .DIN2(n704), .Q(n3761) );
  nnd2s1 U4529 ( .DIN1(n3763), .DIN2(n3764), .Q(\IDinst/n5034 ) );
  nnd2s1 U4530 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][27] ), .Q(n3764) );
  nnd2s1 U4531 ( .DIN1(n600), .DIN2(n704), .Q(n3763) );
  nnd2s1 U4532 ( .DIN1(n3765), .DIN2(n3766), .Q(\IDinst/n5033 ) );
  nnd2s1 U4533 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][27] ), .Q(n3766) );
  nnd2s1 U4534 ( .DIN1(n602), .DIN2(n704), .Q(n3765) );
  nnd2s1 U4535 ( .DIN1(n3767), .DIN2(n3768), .Q(\IDinst/n5032 ) );
  nnd2s1 U4536 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][27] ), .Q(n3768) );
  nnd2s1 U4537 ( .DIN1(n588), .DIN2(n704), .Q(n3767) );
  nnd2s1 U4538 ( .DIN1(n3769), .DIN2(n3770), .Q(\IDinst/n5031 ) );
  nnd2s1 U4539 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][27] ), .Q(n3770) );
  nnd2s1 U4540 ( .DIN1(n590), .DIN2(n704), .Q(n3769) );
  nnd2s1 U4541 ( .DIN1(n3771), .DIN2(n3772), .Q(\IDinst/n5030 ) );
  nnd2s1 U4542 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][27] ), .Q(n3772) );
  nnd2s1 U4543 ( .DIN1(n592), .DIN2(n704), .Q(n3771) );
  nnd2s1 U4544 ( .DIN1(n3773), .DIN2(n3774), .Q(\IDinst/n5029 ) );
  nnd2s1 U4545 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][27] ), .Q(n3774) );
  nnd2s1 U4546 ( .DIN1(n594), .DIN2(n704), .Q(n3773) );
  nnd2s1 U4547 ( .DIN1(n3775), .DIN2(n3776), .Q(\IDinst/n5028 ) );
  nnd2s1 U4548 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][27] ), .Q(n3776) );
  nnd2s1 U4549 ( .DIN1(n612), .DIN2(n704), .Q(n3775) );
  nnd2s1 U4550 ( .DIN1(n3777), .DIN2(n3778), .Q(\IDinst/n5027 ) );
  nnd2s1 U4551 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][27] ), .Q(n3778) );
  nnd2s1 U4552 ( .DIN1(n614), .DIN2(n704), .Q(n3777) );
  nnd2s1 U4553 ( .DIN1(n3779), .DIN2(n3780), .Q(\IDinst/n5026 ) );
  nnd2s1 U4554 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][27] ), .Q(n3780) );
  nnd2s1 U4555 ( .DIN1(n616), .DIN2(n704), .Q(n3779) );
  nnd2s1 U4556 ( .DIN1(n3781), .DIN2(n3782), .Q(\IDinst/n5025 ) );
  nnd2s1 U4557 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][27] ), .Q(n3782) );
  nnd2s1 U4558 ( .DIN1(n618), .DIN2(n704), .Q(n3781) );
  nnd2s1 U4559 ( .DIN1(n3783), .DIN2(n3784), .Q(\IDinst/n5024 ) );
  nnd2s1 U4560 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][27] ), .Q(n3784) );
  nnd2s1 U4561 ( .DIN1(n604), .DIN2(n704), .Q(n3783) );
  nnd2s1 U4562 ( .DIN1(n3785), .DIN2(n3786), .Q(\IDinst/n5023 ) );
  nnd2s1 U4563 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][27] ), .Q(n3786) );
  nnd2s1 U4564 ( .DIN1(n606), .DIN2(n3760), .Q(n3785) );
  nnd2s1 U4565 ( .DIN1(n3787), .DIN2(n3788), .Q(\IDinst/n5022 ) );
  nnd2s1 U4566 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][27] ), .Q(n3788) );
  nnd2s1 U4567 ( .DIN1(n608), .DIN2(n3760), .Q(n3787) );
  nnd2s1 U4568 ( .DIN1(n3789), .DIN2(n3790), .Q(\IDinst/n5021 ) );
  nnd2s1 U4569 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][27] ), .Q(n3790) );
  nnd2s1 U4570 ( .DIN1(n610), .DIN2(n3760), .Q(n3789) );
  nnd2s1 U4571 ( .DIN1(n3791), .DIN2(n3792), .Q(\IDinst/n5020 ) );
  nnd2s1 U4572 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][27] ), .Q(n3792) );
  nnd2s1 U4573 ( .DIN1(n580), .DIN2(n3760), .Q(n3791) );
  nnd2s1 U4574 ( .DIN1(n3793), .DIN2(n3794), .Q(\IDinst/n5019 ) );
  nnd2s1 U4575 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][27] ), .Q(n3794) );
  nnd2s1 U4576 ( .DIN1(n582), .DIN2(n3760), .Q(n3793) );
  nnd2s1 U4577 ( .DIN1(n3795), .DIN2(n3796), .Q(\IDinst/n5018 ) );
  nnd2s1 U4578 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][27] ), .Q(n3796) );
  nnd2s1 U4579 ( .DIN1(n584), .DIN2(n3760), .Q(n3795) );
  nnd2s1 U4580 ( .DIN1(n3797), .DIN2(n3798), .Q(\IDinst/n5017 ) );
  nnd2s1 U4581 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][27] ), .Q(n3798) );
  nnd2s1 U4582 ( .DIN1(n586), .DIN2(n3760), .Q(n3797) );
  nnd2s1 U4583 ( .DIN1(n3799), .DIN2(n3800), .Q(\IDinst/n5016 ) );
  nnd2s1 U4584 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][27] ), .Q(n3800) );
  nnd2s1 U4585 ( .DIN1(n572), .DIN2(n3760), .Q(n3799) );
  nnd2s1 U4586 ( .DIN1(n3801), .DIN2(n3802), .Q(\IDinst/n5015 ) );
  nnd2s1 U4587 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][27] ), .Q(n3802) );
  nnd2s1 U4588 ( .DIN1(n574), .DIN2(n3760), .Q(n3801) );
  nnd2s1 U4589 ( .DIN1(n3803), .DIN2(n3804), .Q(\IDinst/n5014 ) );
  nnd2s1 U4590 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][27] ), .Q(n3804) );
  nnd2s1 U4591 ( .DIN1(n576), .DIN2(n3760), .Q(n3803) );
  nnd2s1 U4592 ( .DIN1(n3805), .DIN2(n3806), .Q(\IDinst/n5013 ) );
  nnd2s1 U4593 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][27] ), .Q(n3806) );
  nnd2s1 U4594 ( .DIN1(n578), .DIN2(n3760), .Q(n3805) );
  nnd2s1 U4595 ( .DIN1(n3807), .DIN2(n3808), .Q(\IDinst/n5012 ) );
  nnd2s1 U4596 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][27] ), .Q(n3808) );
  nnd2s1 U4597 ( .DIN1(n564), .DIN2(n3760), .Q(n3807) );
  nnd2s1 U4598 ( .DIN1(n3809), .DIN2(n3810), .Q(\IDinst/n5011 ) );
  nnd2s1 U4599 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][27] ), .Q(n3810) );
  nnd2s1 U4600 ( .DIN1(n566), .DIN2(n3760), .Q(n3809) );
  nnd2s1 U4601 ( .DIN1(n3811), .DIN2(n3812), .Q(\IDinst/n5010 ) );
  nnd2s1 U4602 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][27] ), .Q(n3812) );
  nnd2s1 U4603 ( .DIN1(n568), .DIN2(n3760), .Q(n3811) );
  nnd2s1 U4604 ( .DIN1(n3813), .DIN2(n3814), .Q(\IDinst/n5009 ) );
  nnd2s1 U4605 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][27] ), .Q(n3814) );
  nnd2s1 U4606 ( .DIN1(n570), .DIN2(n3760), .Q(n3813) );
  nnd2s1 U4607 ( .DIN1(n3815), .DIN2(n3816), .Q(\IDinst/n5008 ) );
  nnd2s1 U4608 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][27] ), .Q(n3816) );
  nnd2s1 U4609 ( .DIN1(n556), .DIN2(n3760), .Q(n3815) );
  nnd2s1 U4610 ( .DIN1(n3817), .DIN2(n3818), .Q(\IDinst/n5007 ) );
  nnd2s1 U4611 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][27] ), .Q(n3818) );
  nnd2s1 U4612 ( .DIN1(n558), .DIN2(n3760), .Q(n3817) );
  nnd2s1 U4613 ( .DIN1(n3819), .DIN2(n3820), .Q(\IDinst/n5006 ) );
  nnd2s1 U4614 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][27] ), .Q(n3820) );
  nnd2s1 U4615 ( .DIN1(n560), .DIN2(n3760), .Q(n3819) );
  nnd2s1 U4616 ( .DIN1(n3821), .DIN2(n3822), .Q(\IDinst/n5005 ) );
  nnd2s1 U4617 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][27] ), .Q(n3822) );
  nnd2s1 U4618 ( .DIN1(n562), .DIN2(n3760), .Q(n3821) );
  nnd2s1 U4619 ( .DIN1(n3035), .DIN2(n3823), .Q(n3760) );
  nnd2s1 U4620 ( .DIN1(n3103), .DIN2(n163), .Q(n3823) );
  nnd2s1 U4621 ( .DIN1(n3824), .DIN2(n3825), .Q(\IDinst/n5004 ) );
  nnd2s1 U4622 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][28] ), .Q(n3825) );
  nnd2s1 U4623 ( .DIN1(n597), .DIN2(n710), .Q(n3824) );
  nnd2s1 U4624 ( .DIN1(n3827), .DIN2(n3828), .Q(\IDinst/n5003 ) );
  nnd2s1 U4625 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][28] ), .Q(n3828) );
  nnd2s1 U4626 ( .DIN1(n599), .DIN2(n710), .Q(n3827) );
  nnd2s1 U4627 ( .DIN1(n3829), .DIN2(n3830), .Q(\IDinst/n5002 ) );
  nnd2s1 U4628 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][28] ), .Q(n3830) );
  nnd2s1 U4629 ( .DIN1(n601), .DIN2(n710), .Q(n3829) );
  nnd2s1 U4630 ( .DIN1(n3831), .DIN2(n3832), .Q(\IDinst/n5001 ) );
  nnd2s1 U4631 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][28] ), .Q(n3832) );
  nnd2s1 U4632 ( .DIN1(n603), .DIN2(n710), .Q(n3831) );
  nnd2s1 U4633 ( .DIN1(n3833), .DIN2(n3834), .Q(\IDinst/n5000 ) );
  nnd2s1 U4634 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][28] ), .Q(n3834) );
  nnd2s1 U4635 ( .DIN1(n589), .DIN2(n710), .Q(n3833) );
  nnd2s1 U4636 ( .DIN1(n3835), .DIN2(n3836), .Q(\IDinst/n4999 ) );
  nnd2s1 U4637 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][28] ), .Q(n3836) );
  nnd2s1 U4638 ( .DIN1(n591), .DIN2(n710), .Q(n3835) );
  nnd2s1 U4639 ( .DIN1(n3837), .DIN2(n3838), .Q(\IDinst/n4998 ) );
  nnd2s1 U4640 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][28] ), .Q(n3838) );
  nnd2s1 U4641 ( .DIN1(n593), .DIN2(n710), .Q(n3837) );
  nnd2s1 U4642 ( .DIN1(n3839), .DIN2(n3840), .Q(\IDinst/n4997 ) );
  nnd2s1 U4643 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][28] ), .Q(n3840) );
  nnd2s1 U4644 ( .DIN1(n595), .DIN2(n710), .Q(n3839) );
  nnd2s1 U4645 ( .DIN1(n3841), .DIN2(n3842), .Q(\IDinst/n4996 ) );
  nnd2s1 U4646 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][28] ), .Q(n3842) );
  nnd2s1 U4647 ( .DIN1(n613), .DIN2(n710), .Q(n3841) );
  nnd2s1 U4648 ( .DIN1(n3843), .DIN2(n3844), .Q(\IDinst/n4995 ) );
  nnd2s1 U4649 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][28] ), .Q(n3844) );
  nnd2s1 U4650 ( .DIN1(n615), .DIN2(n710), .Q(n3843) );
  nnd2s1 U4651 ( .DIN1(n3845), .DIN2(n3846), .Q(\IDinst/n4994 ) );
  nnd2s1 U4652 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][28] ), .Q(n3846) );
  nnd2s1 U4653 ( .DIN1(n617), .DIN2(n710), .Q(n3845) );
  nnd2s1 U4654 ( .DIN1(n3847), .DIN2(n3848), .Q(\IDinst/n4993 ) );
  nnd2s1 U4655 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][28] ), .Q(n3848) );
  nnd2s1 U4656 ( .DIN1(n619), .DIN2(n710), .Q(n3847) );
  nnd2s1 U4657 ( .DIN1(n3849), .DIN2(n3850), .Q(\IDinst/n4992 ) );
  nnd2s1 U4658 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][28] ), .Q(n3850) );
  nnd2s1 U4659 ( .DIN1(n605), .DIN2(n710), .Q(n3849) );
  nnd2s1 U4660 ( .DIN1(n3851), .DIN2(n3852), .Q(\IDinst/n4991 ) );
  nnd2s1 U4661 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][28] ), .Q(n3852) );
  nnd2s1 U4662 ( .DIN1(n607), .DIN2(n3826), .Q(n3851) );
  nnd2s1 U4663 ( .DIN1(n3853), .DIN2(n3854), .Q(\IDinst/n4990 ) );
  nnd2s1 U4664 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][28] ), .Q(n3854) );
  nnd2s1 U4665 ( .DIN1(n609), .DIN2(n3826), .Q(n3853) );
  nnd2s1 U4666 ( .DIN1(n3855), .DIN2(n3856), .Q(\IDinst/n4989 ) );
  nnd2s1 U4667 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][28] ), .Q(n3856) );
  nnd2s1 U4668 ( .DIN1(n611), .DIN2(n3826), .Q(n3855) );
  nnd2s1 U4669 ( .DIN1(n3857), .DIN2(n3858), .Q(\IDinst/n4988 ) );
  nnd2s1 U4670 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][28] ), .Q(n3858) );
  nnd2s1 U4671 ( .DIN1(n581), .DIN2(n3826), .Q(n3857) );
  nnd2s1 U4672 ( .DIN1(n3859), .DIN2(n3860), .Q(\IDinst/n4987 ) );
  nnd2s1 U4673 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][28] ), .Q(n3860) );
  nnd2s1 U4674 ( .DIN1(n583), .DIN2(n3826), .Q(n3859) );
  nnd2s1 U4675 ( .DIN1(n3861), .DIN2(n3862), .Q(\IDinst/n4986 ) );
  nnd2s1 U4676 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][28] ), .Q(n3862) );
  nnd2s1 U4677 ( .DIN1(n585), .DIN2(n3826), .Q(n3861) );
  nnd2s1 U4678 ( .DIN1(n3863), .DIN2(n3864), .Q(\IDinst/n4985 ) );
  nnd2s1 U4679 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][28] ), .Q(n3864) );
  nnd2s1 U4680 ( .DIN1(n587), .DIN2(n3826), .Q(n3863) );
  nnd2s1 U4681 ( .DIN1(n3865), .DIN2(n3866), .Q(\IDinst/n4984 ) );
  nnd2s1 U4682 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][28] ), .Q(n3866) );
  nnd2s1 U4683 ( .DIN1(n573), .DIN2(n3826), .Q(n3865) );
  nnd2s1 U4684 ( .DIN1(n3867), .DIN2(n3868), .Q(\IDinst/n4983 ) );
  nnd2s1 U4685 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][28] ), .Q(n3868) );
  nnd2s1 U4686 ( .DIN1(n575), .DIN2(n3826), .Q(n3867) );
  nnd2s1 U4687 ( .DIN1(n3869), .DIN2(n3870), .Q(\IDinst/n4982 ) );
  nnd2s1 U4688 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][28] ), .Q(n3870) );
  nnd2s1 U4689 ( .DIN1(n577), .DIN2(n3826), .Q(n3869) );
  nnd2s1 U4690 ( .DIN1(n3871), .DIN2(n3872), .Q(\IDinst/n4981 ) );
  nnd2s1 U4691 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][28] ), .Q(n3872) );
  nnd2s1 U4692 ( .DIN1(n579), .DIN2(n3826), .Q(n3871) );
  nnd2s1 U4693 ( .DIN1(n3873), .DIN2(n3874), .Q(\IDinst/n4980 ) );
  nnd2s1 U4694 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][28] ), .Q(n3874) );
  nnd2s1 U4695 ( .DIN1(n565), .DIN2(n3826), .Q(n3873) );
  nnd2s1 U4696 ( .DIN1(n3875), .DIN2(n3876), .Q(\IDinst/n4979 ) );
  nnd2s1 U4697 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][28] ), .Q(n3876) );
  nnd2s1 U4698 ( .DIN1(n567), .DIN2(n3826), .Q(n3875) );
  nnd2s1 U4699 ( .DIN1(n3877), .DIN2(n3878), .Q(\IDinst/n4978 ) );
  nnd2s1 U4700 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][28] ), .Q(n3878) );
  nnd2s1 U4701 ( .DIN1(n569), .DIN2(n3826), .Q(n3877) );
  nnd2s1 U4702 ( .DIN1(n3879), .DIN2(n3880), .Q(\IDinst/n4977 ) );
  nnd2s1 U4703 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][28] ), .Q(n3880) );
  nnd2s1 U4704 ( .DIN1(n571), .DIN2(n3826), .Q(n3879) );
  nnd2s1 U4705 ( .DIN1(n3881), .DIN2(n3882), .Q(\IDinst/n4976 ) );
  nnd2s1 U4706 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][28] ), .Q(n3882) );
  nnd2s1 U4707 ( .DIN1(n557), .DIN2(n3826), .Q(n3881) );
  nnd2s1 U4708 ( .DIN1(n3883), .DIN2(n3884), .Q(\IDinst/n4975 ) );
  nnd2s1 U4709 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][28] ), .Q(n3884) );
  nnd2s1 U4710 ( .DIN1(n559), .DIN2(n3826), .Q(n3883) );
  nnd2s1 U4711 ( .DIN1(n3885), .DIN2(n3886), .Q(\IDinst/n4974 ) );
  nnd2s1 U4712 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][28] ), .Q(n3886) );
  nnd2s1 U4713 ( .DIN1(n561), .DIN2(n3826), .Q(n3885) );
  nnd2s1 U4714 ( .DIN1(n3887), .DIN2(n3888), .Q(\IDinst/n4973 ) );
  nnd2s1 U4715 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][28] ), .Q(n3888) );
  nnd2s1 U4716 ( .DIN1(n563), .DIN2(n3826), .Q(n3887) );
  nnd2s1 U4717 ( .DIN1(n3035), .DIN2(n3889), .Q(n3826) );
  nnd2s1 U4718 ( .DIN1(n3103), .DIN2(n161), .Q(n3889) );
  nnd2s1 U4719 ( .DIN1(n3890), .DIN2(n3891), .Q(\IDinst/n4972 ) );
  nnd2s1 U4720 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][29] ), .Q(n3891) );
  nnd2s1 U4721 ( .DIN1(n596), .DIN2(n724), .Q(n3890) );
  nnd2s1 U4722 ( .DIN1(n3893), .DIN2(n3894), .Q(\IDinst/n4971 ) );
  nnd2s1 U4723 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][29] ), .Q(n3894) );
  nnd2s1 U4724 ( .DIN1(n598), .DIN2(n3892), .Q(n3893) );
  nnd2s1 U4725 ( .DIN1(n3895), .DIN2(n3896), .Q(\IDinst/n4970 ) );
  nnd2s1 U4726 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][29] ), .Q(n3896) );
  nnd2s1 U4727 ( .DIN1(n600), .DIN2(n724), .Q(n3895) );
  nnd2s1 U4728 ( .DIN1(n3897), .DIN2(n3898), .Q(\IDinst/n4969 ) );
  nnd2s1 U4729 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][29] ), .Q(n3898) );
  nnd2s1 U4730 ( .DIN1(n602), .DIN2(n3892), .Q(n3897) );
  nnd2s1 U4731 ( .DIN1(n3899), .DIN2(n3900), .Q(\IDinst/n4968 ) );
  nnd2s1 U4732 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][29] ), .Q(n3900) );
  nnd2s1 U4733 ( .DIN1(n588), .DIN2(n724), .Q(n3899) );
  nnd2s1 U4734 ( .DIN1(n3901), .DIN2(n3902), .Q(\IDinst/n4967 ) );
  nnd2s1 U4735 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][29] ), .Q(n3902) );
  nnd2s1 U4736 ( .DIN1(n590), .DIN2(n3892), .Q(n3901) );
  nnd2s1 U4737 ( .DIN1(n3903), .DIN2(n3904), .Q(\IDinst/n4966 ) );
  nnd2s1 U4738 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][29] ), .Q(n3904) );
  nnd2s1 U4739 ( .DIN1(n592), .DIN2(n724), .Q(n3903) );
  nnd2s1 U4740 ( .DIN1(n3905), .DIN2(n3906), .Q(\IDinst/n4965 ) );
  nnd2s1 U4741 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][29] ), .Q(n3906) );
  nnd2s1 U4742 ( .DIN1(n594), .DIN2(n3892), .Q(n3905) );
  nnd2s1 U4743 ( .DIN1(n3907), .DIN2(n3908), .Q(\IDinst/n4964 ) );
  nnd2s1 U4744 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][29] ), .Q(n3908) );
  nnd2s1 U4745 ( .DIN1(n612), .DIN2(n724), .Q(n3907) );
  nnd2s1 U4746 ( .DIN1(n3909), .DIN2(n3910), .Q(\IDinst/n4963 ) );
  nnd2s1 U4747 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][29] ), .Q(n3910) );
  nnd2s1 U4748 ( .DIN1(n614), .DIN2(n3892), .Q(n3909) );
  nnd2s1 U4749 ( .DIN1(n3911), .DIN2(n3912), .Q(\IDinst/n4962 ) );
  nnd2s1 U4750 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][29] ), .Q(n3912) );
  nnd2s1 U4751 ( .DIN1(n616), .DIN2(n724), .Q(n3911) );
  nnd2s1 U4752 ( .DIN1(n3913), .DIN2(n3914), .Q(\IDinst/n4961 ) );
  nnd2s1 U4753 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][29] ), .Q(n3914) );
  nnd2s1 U4754 ( .DIN1(n618), .DIN2(n3892), .Q(n3913) );
  nnd2s1 U4755 ( .DIN1(n3915), .DIN2(n3916), .Q(\IDinst/n4960 ) );
  nnd2s1 U4756 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][29] ), .Q(n3916) );
  nnd2s1 U4757 ( .DIN1(n604), .DIN2(n724), .Q(n3915) );
  nnd2s1 U4758 ( .DIN1(n3917), .DIN2(n3918), .Q(\IDinst/n4959 ) );
  nnd2s1 U4759 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][29] ), .Q(n3918) );
  nnd2s1 U4760 ( .DIN1(n606), .DIN2(n3892), .Q(n3917) );
  nnd2s1 U4761 ( .DIN1(n3919), .DIN2(n3920), .Q(\IDinst/n4958 ) );
  nnd2s1 U4762 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][29] ), .Q(n3920) );
  nnd2s1 U4763 ( .DIN1(n608), .DIN2(n724), .Q(n3919) );
  nnd2s1 U4764 ( .DIN1(n3921), .DIN2(n3922), .Q(\IDinst/n4957 ) );
  nnd2s1 U4765 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][29] ), .Q(n3922) );
  nnd2s1 U4766 ( .DIN1(n610), .DIN2(n3892), .Q(n3921) );
  nnd2s1 U4767 ( .DIN1(n3923), .DIN2(n3924), .Q(\IDinst/n4956 ) );
  nnd2s1 U4768 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][29] ), .Q(n3924) );
  nnd2s1 U4769 ( .DIN1(n580), .DIN2(n724), .Q(n3923) );
  nnd2s1 U4770 ( .DIN1(n3925), .DIN2(n3926), .Q(\IDinst/n4955 ) );
  nnd2s1 U4771 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][29] ), .Q(n3926) );
  nnd2s1 U4772 ( .DIN1(n582), .DIN2(n3892), .Q(n3925) );
  nnd2s1 U4773 ( .DIN1(n3927), .DIN2(n3928), .Q(\IDinst/n4954 ) );
  nnd2s1 U4774 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][29] ), .Q(n3928) );
  nnd2s1 U4775 ( .DIN1(n584), .DIN2(n724), .Q(n3927) );
  nnd2s1 U4776 ( .DIN1(n3929), .DIN2(n3930), .Q(\IDinst/n4953 ) );
  nnd2s1 U4777 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][29] ), .Q(n3930) );
  nnd2s1 U4778 ( .DIN1(n586), .DIN2(n3892), .Q(n3929) );
  nnd2s1 U4779 ( .DIN1(n3931), .DIN2(n3932), .Q(\IDinst/n4952 ) );
  nnd2s1 U4780 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][29] ), .Q(n3932) );
  nnd2s1 U4781 ( .DIN1(n572), .DIN2(n724), .Q(n3931) );
  nnd2s1 U4782 ( .DIN1(n3933), .DIN2(n3934), .Q(\IDinst/n4951 ) );
  nnd2s1 U4783 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][29] ), .Q(n3934) );
  nnd2s1 U4784 ( .DIN1(n574), .DIN2(n3892), .Q(n3933) );
  nnd2s1 U4785 ( .DIN1(n3935), .DIN2(n3936), .Q(\IDinst/n4950 ) );
  nnd2s1 U4786 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][29] ), .Q(n3936) );
  nnd2s1 U4787 ( .DIN1(n576), .DIN2(n724), .Q(n3935) );
  nnd2s1 U4788 ( .DIN1(n3937), .DIN2(n3938), .Q(\IDinst/n4949 ) );
  nnd2s1 U4789 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][29] ), .Q(n3938) );
  nnd2s1 U4790 ( .DIN1(n578), .DIN2(n3892), .Q(n3937) );
  nnd2s1 U4791 ( .DIN1(n3939), .DIN2(n3940), .Q(\IDinst/n4948 ) );
  nnd2s1 U4792 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][29] ), .Q(n3940) );
  nnd2s1 U4793 ( .DIN1(n564), .DIN2(n724), .Q(n3939) );
  nnd2s1 U4794 ( .DIN1(n3941), .DIN2(n3942), .Q(\IDinst/n4947 ) );
  nnd2s1 U4795 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][29] ), .Q(n3942) );
  nnd2s1 U4796 ( .DIN1(n566), .DIN2(n3892), .Q(n3941) );
  nnd2s1 U4797 ( .DIN1(n3943), .DIN2(n3944), .Q(\IDinst/n4946 ) );
  nnd2s1 U4798 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][29] ), .Q(n3944) );
  nnd2s1 U4799 ( .DIN1(n568), .DIN2(n724), .Q(n3943) );
  nnd2s1 U4800 ( .DIN1(n3945), .DIN2(n3946), .Q(\IDinst/n4945 ) );
  nnd2s1 U4801 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][29] ), .Q(n3946) );
  nnd2s1 U4802 ( .DIN1(n570), .DIN2(n3892), .Q(n3945) );
  nnd2s1 U4803 ( .DIN1(n3947), .DIN2(n3948), .Q(\IDinst/n4944 ) );
  nnd2s1 U4804 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][29] ), .Q(n3948) );
  nnd2s1 U4805 ( .DIN1(n556), .DIN2(n724), .Q(n3947) );
  nnd2s1 U4806 ( .DIN1(n3949), .DIN2(n3950), .Q(\IDinst/n4943 ) );
  nnd2s1 U4807 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][29] ), .Q(n3950) );
  nnd2s1 U4808 ( .DIN1(n558), .DIN2(n3892), .Q(n3949) );
  nnd2s1 U4809 ( .DIN1(n3951), .DIN2(n3952), .Q(\IDinst/n4942 ) );
  nnd2s1 U4810 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][29] ), .Q(n3952) );
  nnd2s1 U4811 ( .DIN1(n560), .DIN2(n724), .Q(n3951) );
  nnd2s1 U4812 ( .DIN1(n3953), .DIN2(n3954), .Q(\IDinst/n4941 ) );
  nnd2s1 U4813 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][29] ), .Q(n3954) );
  nnd2s1 U4814 ( .DIN1(n562), .DIN2(n3892), .Q(n3953) );
  nnd2s1 U4815 ( .DIN1(n3035), .DIN2(n3955), .Q(n3892) );
  nnd2s1 U4816 ( .DIN1(n3103), .DIN2(n159), .Q(n3955) );
  nnd2s1 U4817 ( .DIN1(n3956), .DIN2(n3957), .Q(\IDinst/n4940 ) );
  nnd2s1 U4818 ( .DIN1(n483), .DIN2(\IDinst/RegFile[0][30] ), .Q(n3957) );
  nnd2s1 U4819 ( .DIN1(n597), .DIN2(n738), .Q(n3956) );
  nnd2s1 U4820 ( .DIN1(n3959), .DIN2(n3960), .Q(\IDinst/n4939 ) );
  nnd2s1 U4821 ( .DIN1(n507), .DIN2(\IDinst/RegFile[1][30] ), .Q(n3960) );
  nnd2s1 U4822 ( .DIN1(n599), .DIN2(n3958), .Q(n3959) );
  nnd2s1 U4823 ( .DIN1(n3961), .DIN2(n3962), .Q(\IDinst/n4938 ) );
  nnd2s1 U4824 ( .DIN1(n521), .DIN2(\IDinst/RegFile[2][30] ), .Q(n3962) );
  nnd2s1 U4825 ( .DIN1(n601), .DIN2(n738), .Q(n3961) );
  nnd2s1 U4826 ( .DIN1(n3963), .DIN2(n3964), .Q(\IDinst/n4937 ) );
  nnd2s1 U4827 ( .DIN1(n501), .DIN2(\IDinst/RegFile[3][30] ), .Q(n3964) );
  nnd2s1 U4828 ( .DIN1(n603), .DIN2(n3958), .Q(n3963) );
  nnd2s1 U4829 ( .DIN1(n3965), .DIN2(n3966), .Q(\IDinst/n4936 ) );
  nnd2s1 U4830 ( .DIN1(n523), .DIN2(\IDinst/RegFile[4][30] ), .Q(n3966) );
  nnd2s1 U4831 ( .DIN1(n589), .DIN2(n738), .Q(n3965) );
  nnd2s1 U4832 ( .DIN1(n3967), .DIN2(n3968), .Q(\IDinst/n4935 ) );
  nnd2s1 U4833 ( .DIN1(n503), .DIN2(\IDinst/RegFile[5][30] ), .Q(n3968) );
  nnd2s1 U4834 ( .DIN1(n591), .DIN2(n3958), .Q(n3967) );
  nnd2s1 U4835 ( .DIN1(n3969), .DIN2(n3970), .Q(\IDinst/n4934 ) );
  nnd2s1 U4836 ( .DIN1(n517), .DIN2(\IDinst/RegFile[6][30] ), .Q(n3970) );
  nnd2s1 U4837 ( .DIN1(n593), .DIN2(n738), .Q(n3969) );
  nnd2s1 U4838 ( .DIN1(n3971), .DIN2(n3972), .Q(\IDinst/n4933 ) );
  nnd2s1 U4839 ( .DIN1(n485), .DIN2(\IDinst/RegFile[7][30] ), .Q(n3972) );
  nnd2s1 U4840 ( .DIN1(n595), .DIN2(n3958), .Q(n3971) );
  nnd2s1 U4841 ( .DIN1(n3973), .DIN2(n3974), .Q(\IDinst/n4932 ) );
  nnd2s1 U4842 ( .DIN1(n477), .DIN2(\IDinst/RegFile[8][30] ), .Q(n3974) );
  nnd2s1 U4843 ( .DIN1(n613), .DIN2(n738), .Q(n3973) );
  nnd2s1 U4844 ( .DIN1(n3975), .DIN2(n3976), .Q(\IDinst/n4931 ) );
  nnd2s1 U4845 ( .DIN1(n497), .DIN2(\IDinst/RegFile[9][30] ), .Q(n3976) );
  nnd2s1 U4846 ( .DIN1(n615), .DIN2(n3958), .Q(n3975) );
  nnd2s1 U4847 ( .DIN1(n3977), .DIN2(n3978), .Q(\IDinst/n4930 ) );
  nnd2s1 U4848 ( .DIN1(n519), .DIN2(\IDinst/RegFile[10][30] ), .Q(n3978) );
  nnd2s1 U4849 ( .DIN1(n617), .DIN2(n738), .Q(n3977) );
  nnd2s1 U4850 ( .DIN1(n3979), .DIN2(n3980), .Q(\IDinst/n4929 ) );
  nnd2s1 U4851 ( .DIN1(n499), .DIN2(\IDinst/RegFile[11][30] ), .Q(n3980) );
  nnd2s1 U4852 ( .DIN1(n619), .DIN2(n3958), .Q(n3979) );
  nnd2s1 U4853 ( .DIN1(n3981), .DIN2(n3982), .Q(\IDinst/n4928 ) );
  nnd2s1 U4854 ( .DIN1(n513), .DIN2(\IDinst/RegFile[12][30] ), .Q(n3982) );
  nnd2s1 U4855 ( .DIN1(n605), .DIN2(n738), .Q(n3981) );
  nnd2s1 U4856 ( .DIN1(n3983), .DIN2(n3984), .Q(\IDinst/n4927 ) );
  nnd2s1 U4857 ( .DIN1(n493), .DIN2(\IDinst/RegFile[13][30] ), .Q(n3984) );
  nnd2s1 U4858 ( .DIN1(n607), .DIN2(n3958), .Q(n3983) );
  nnd2s1 U4859 ( .DIN1(n3985), .DIN2(n3986), .Q(\IDinst/n4926 ) );
  nnd2s1 U4860 ( .DIN1(n515), .DIN2(\IDinst/RegFile[14][30] ), .Q(n3986) );
  nnd2s1 U4861 ( .DIN1(n609), .DIN2(n738), .Q(n3985) );
  nnd2s1 U4862 ( .DIN1(n3987), .DIN2(n3988), .Q(\IDinst/n4925 ) );
  nnd2s1 U4863 ( .DIN1(n487), .DIN2(\IDinst/RegFile[15][30] ), .Q(n3988) );
  nnd2s1 U4864 ( .DIN1(n611), .DIN2(n3958), .Q(n3987) );
  nnd2s1 U4865 ( .DIN1(n3989), .DIN2(n3990), .Q(\IDinst/n4924 ) );
  nnd2s1 U4866 ( .DIN1(n479), .DIN2(\IDinst/RegFile[16][30] ), .Q(n3990) );
  nnd2s1 U4867 ( .DIN1(n581), .DIN2(n738), .Q(n3989) );
  nnd2s1 U4868 ( .DIN1(n3991), .DIN2(n3992), .Q(\IDinst/n4923 ) );
  nnd2s1 U4869 ( .DIN1(n495), .DIN2(\IDinst/RegFile[17][30] ), .Q(n3992) );
  nnd2s1 U4870 ( .DIN1(n583), .DIN2(n3958), .Q(n3991) );
  nnd2s1 U4871 ( .DIN1(n3993), .DIN2(n3994), .Q(\IDinst/n4922 ) );
  nnd2s1 U4872 ( .DIN1(n509), .DIN2(\IDinst/RegFile[18][30] ), .Q(n3994) );
  nnd2s1 U4873 ( .DIN1(n585), .DIN2(n738), .Q(n3993) );
  nnd2s1 U4874 ( .DIN1(n3995), .DIN2(n3996), .Q(\IDinst/n4921 ) );
  nnd2s1 U4875 ( .DIN1(n489), .DIN2(\IDinst/RegFile[19][30] ), .Q(n3996) );
  nnd2s1 U4876 ( .DIN1(n587), .DIN2(n3958), .Q(n3995) );
  nnd2s1 U4877 ( .DIN1(n3997), .DIN2(n3998), .Q(\IDinst/n4920 ) );
  nnd2s1 U4878 ( .DIN1(n511), .DIN2(\IDinst/RegFile[20][30] ), .Q(n3998) );
  nnd2s1 U4879 ( .DIN1(n573), .DIN2(n738), .Q(n3997) );
  nnd2s1 U4880 ( .DIN1(n3999), .DIN2(n4000), .Q(\IDinst/n4919 ) );
  nnd2s1 U4881 ( .DIN1(n491), .DIN2(\IDinst/RegFile[21][30] ), .Q(n4000) );
  nnd2s1 U4882 ( .DIN1(n575), .DIN2(n3958), .Q(n3999) );
  nnd2s1 U4883 ( .DIN1(n4001), .DIN2(n4002), .Q(\IDinst/n4918 ) );
  nnd2s1 U4884 ( .DIN1(n505), .DIN2(\IDinst/RegFile[22][30] ), .Q(n4002) );
  nnd2s1 U4885 ( .DIN1(n577), .DIN2(n738), .Q(n4001) );
  nnd2s1 U4886 ( .DIN1(n4003), .DIN2(n4004), .Q(\IDinst/n4917 ) );
  nnd2s1 U4887 ( .DIN1(n481), .DIN2(\IDinst/RegFile[23][30] ), .Q(n4004) );
  nnd2s1 U4888 ( .DIN1(n579), .DIN2(n3958), .Q(n4003) );
  nnd2s1 U4889 ( .DIN1(n4005), .DIN2(n4006), .Q(\IDinst/n4916 ) );
  nnd2s1 U4890 ( .DIN1(n473), .DIN2(\IDinst/RegFile[24][30] ), .Q(n4006) );
  nnd2s1 U4891 ( .DIN1(n565), .DIN2(n738), .Q(n4005) );
  nnd2s1 U4892 ( .DIN1(n4007), .DIN2(n4008), .Q(\IDinst/n4915 ) );
  nnd2s1 U4893 ( .DIN1(n475), .DIN2(\IDinst/RegFile[25][30] ), .Q(n4008) );
  nnd2s1 U4894 ( .DIN1(n567), .DIN2(n3958), .Q(n4007) );
  nnd2s1 U4895 ( .DIN1(n4009), .DIN2(n4010), .Q(\IDinst/n4914 ) );
  nnd2s1 U4896 ( .DIN1(n469), .DIN2(\IDinst/RegFile[26][30] ), .Q(n4010) );
  nnd2s1 U4897 ( .DIN1(n569), .DIN2(n738), .Q(n4009) );
  nnd2s1 U4898 ( .DIN1(n4011), .DIN2(n4012), .Q(\IDinst/n4913 ) );
  nnd2s1 U4899 ( .DIN1(n471), .DIN2(\IDinst/RegFile[27][30] ), .Q(n4012) );
  nnd2s1 U4900 ( .DIN1(n571), .DIN2(n3958), .Q(n4011) );
  nnd2s1 U4901 ( .DIN1(n4013), .DIN2(n4014), .Q(\IDinst/n4912 ) );
  nnd2s1 U4902 ( .DIN1(n465), .DIN2(\IDinst/RegFile[28][30] ), .Q(n4014) );
  nnd2s1 U4903 ( .DIN1(n557), .DIN2(n738), .Q(n4013) );
  nnd2s1 U4904 ( .DIN1(n4015), .DIN2(n4016), .Q(\IDinst/n4911 ) );
  nnd2s1 U4905 ( .DIN1(n467), .DIN2(\IDinst/RegFile[29][30] ), .Q(n4016) );
  nnd2s1 U4906 ( .DIN1(n559), .DIN2(n3958), .Q(n4015) );
  nnd2s1 U4907 ( .DIN1(n4017), .DIN2(n4018), .Q(\IDinst/n4910 ) );
  nnd2s1 U4908 ( .DIN1(n461), .DIN2(\IDinst/RegFile[30][30] ), .Q(n4018) );
  nnd2s1 U4909 ( .DIN1(n561), .DIN2(n738), .Q(n4017) );
  nnd2s1 U4910 ( .DIN1(n4019), .DIN2(n4020), .Q(\IDinst/n4909 ) );
  nnd2s1 U4911 ( .DIN1(n463), .DIN2(\IDinst/RegFile[31][30] ), .Q(n4020) );
  nnd2s1 U4912 ( .DIN1(n563), .DIN2(n3958), .Q(n4019) );
  nnd2s1 U4913 ( .DIN1(n3035), .DIN2(n4021), .Q(n3958) );
  nnd2s1 U4914 ( .DIN1(n3103), .DIN2(n157), .Q(n4021) );
  nnd2s1 U4915 ( .DIN1(n4022), .DIN2(n4023), .Q(\IDinst/n4908 ) );
  nnd2s1 U4916 ( .DIN1(n482), .DIN2(\IDinst/RegFile[0][31] ), .Q(n4023) );
  nnd2s1 U4917 ( .DIN1(n596), .DIN2(n766), .Q(n4022) );
  nnd2s1 U4918 ( .DIN1(n4026), .DIN2(n4027), .Q(\IDinst/n4907 ) );
  nnd2s1 U4919 ( .DIN1(n506), .DIN2(\IDinst/RegFile[1][31] ), .Q(n4027) );
  nnd2s1 U4920 ( .DIN1(n598), .DIN2(n4024), .Q(n4026) );
  nnd2s1 U4921 ( .DIN1(n4029), .DIN2(n4030), .Q(\IDinst/n4906 ) );
  nnd2s1 U4922 ( .DIN1(n520), .DIN2(\IDinst/RegFile[2][31] ), .Q(n4030) );
  nnd2s1 U4923 ( .DIN1(n600), .DIN2(n766), .Q(n4029) );
  nnd2s1 U4924 ( .DIN1(n4032), .DIN2(n4033), .Q(\IDinst/n4905 ) );
  nnd2s1 U4925 ( .DIN1(n500), .DIN2(\IDinst/RegFile[3][31] ), .Q(n4033) );
  nnd2s1 U4926 ( .DIN1(n602), .DIN2(n4024), .Q(n4032) );
  nnd2s1 U4927 ( .DIN1(n4035), .DIN2(n4036), .Q(\IDinst/n4904 ) );
  nnd2s1 U4928 ( .DIN1(n522), .DIN2(\IDinst/RegFile[4][31] ), .Q(n4036) );
  nnd2s1 U4929 ( .DIN1(n588), .DIN2(n766), .Q(n4035) );
  nnd2s1 U4930 ( .DIN1(n4038), .DIN2(n4039), .Q(\IDinst/n4903 ) );
  nnd2s1 U4931 ( .DIN1(n502), .DIN2(\IDinst/RegFile[5][31] ), .Q(n4039) );
  nnd2s1 U4932 ( .DIN1(n590), .DIN2(n4024), .Q(n4038) );
  nnd2s1 U4933 ( .DIN1(n4041), .DIN2(n4042), .Q(\IDinst/n4902 ) );
  nnd2s1 U4934 ( .DIN1(n516), .DIN2(\IDinst/RegFile[6][31] ), .Q(n4042) );
  nnd2s1 U4935 ( .DIN1(n592), .DIN2(n766), .Q(n4041) );
  nnd2s1 U4936 ( .DIN1(n4044), .DIN2(n4045), .Q(\IDinst/n4901 ) );
  nnd2s1 U4937 ( .DIN1(n484), .DIN2(\IDinst/RegFile[7][31] ), .Q(n4045) );
  nnd2s1 U4938 ( .DIN1(n594), .DIN2(n4024), .Q(n4044) );
  and3s1 U4939 ( .DIN1(\IDinst/n1430 ), .DIN2(\IDinst/n1403 ), 
        .DIN3(reg_write_MEM), .Q(n4025) );
  nnd2s1 U4940 ( .DIN1(n4047), .DIN2(n4048), .Q(\IDinst/n4900 ) );
  nnd2s1 U4941 ( .DIN1(n476), .DIN2(\IDinst/RegFile[8][31] ), .Q(n4048) );
  nnd2s1 U4942 ( .DIN1(n612), .DIN2(n766), .Q(n4047) );
  nnd2s1 U4943 ( .DIN1(n4050), .DIN2(n4051), .Q(\IDinst/n4899 ) );
  nnd2s1 U4944 ( .DIN1(n496), .DIN2(\IDinst/RegFile[9][31] ), .Q(n4051) );
  nnd2s1 U4945 ( .DIN1(n614), .DIN2(n4024), .Q(n4050) );
  nnd2s1 U4946 ( .DIN1(n4052), .DIN2(n4053), .Q(\IDinst/n4898 ) );
  nnd2s1 U4947 ( .DIN1(n518), .DIN2(\IDinst/RegFile[10][31] ), .Q(n4053) );
  nnd2s1 U4948 ( .DIN1(n616), .DIN2(n766), .Q(n4052) );
  nnd2s1 U4949 ( .DIN1(n4054), .DIN2(n4055), .Q(\IDinst/n4897 ) );
  nnd2s1 U4950 ( .DIN1(n498), .DIN2(\IDinst/RegFile[11][31] ), .Q(n4055) );
  nnd2s1 U4951 ( .DIN1(n618), .DIN2(n4024), .Q(n4054) );
  nnd2s1 U4952 ( .DIN1(n4056), .DIN2(n4057), .Q(\IDinst/n4896 ) );
  nnd2s1 U4953 ( .DIN1(n512), .DIN2(\IDinst/RegFile[12][31] ), .Q(n4057) );
  nnd2s1 U4954 ( .DIN1(n604), .DIN2(n766), .Q(n4056) );
  nnd2s1 U4955 ( .DIN1(n4058), .DIN2(n4059), .Q(\IDinst/n4895 ) );
  nnd2s1 U4956 ( .DIN1(n492), .DIN2(\IDinst/RegFile[13][31] ), .Q(n4059) );
  nnd2s1 U4957 ( .DIN1(n606), .DIN2(n4024), .Q(n4058) );
  nnd2s1 U4958 ( .DIN1(n4060), .DIN2(n4061), .Q(\IDinst/n4894 ) );
  nnd2s1 U4959 ( .DIN1(n514), .DIN2(\IDinst/RegFile[14][31] ), .Q(n4061) );
  nnd2s1 U4960 ( .DIN1(n608), .DIN2(n766), .Q(n4060) );
  nnd2s1 U4961 ( .DIN1(n4062), .DIN2(n4063), .Q(\IDinst/n4893 ) );
  nnd2s1 U4962 ( .DIN1(n486), .DIN2(\IDinst/RegFile[15][31] ), .Q(n4063) );
  nnd2s1 U4963 ( .DIN1(n610), .DIN2(n4024), .Q(n4062) );
  and3s1 U4964 ( .DIN1(\IDinst/n1403 ), .DIN2(n47), .DIN3(reg_write_MEM), 
        .Q(n4049) );
  nnd2s1 U4965 ( .DIN1(n4064), .DIN2(n4065), .Q(\IDinst/n4892 ) );
  nnd2s1 U4966 ( .DIN1(n478), .DIN2(\IDinst/RegFile[16][31] ), .Q(n4065) );
  nnd2s1 U4967 ( .DIN1(n580), .DIN2(n766), .Q(n4064) );
  nnd2s1 U4968 ( .DIN1(n4067), .DIN2(n4068), .Q(\IDinst/n4891 ) );
  nnd2s1 U4969 ( .DIN1(n494), .DIN2(\IDinst/RegFile[17][31] ), .Q(n4068) );
  nnd2s1 U4970 ( .DIN1(n582), .DIN2(n4024), .Q(n4067) );
  nnd2s1 U4971 ( .DIN1(n4069), .DIN2(n4070), .Q(\IDinst/n4890 ) );
  nnd2s1 U4972 ( .DIN1(n508), .DIN2(\IDinst/RegFile[18][31] ), .Q(n4070) );
  nnd2s1 U4973 ( .DIN1(n584), .DIN2(n766), .Q(n4069) );
  nnd2s1 U4974 ( .DIN1(n4071), .DIN2(n4072), .Q(\IDinst/n4889 ) );
  nnd2s1 U4975 ( .DIN1(n488), .DIN2(\IDinst/RegFile[19][31] ), .Q(n4072) );
  nnd2s1 U4976 ( .DIN1(n586), .DIN2(n4024), .Q(n4071) );
  nnd2s1 U4977 ( .DIN1(n4073), .DIN2(n4074), .Q(\IDinst/n4888 ) );
  nnd2s1 U4978 ( .DIN1(n510), .DIN2(\IDinst/RegFile[20][31] ), .Q(n4074) );
  nnd2s1 U4979 ( .DIN1(n572), .DIN2(n766), .Q(n4073) );
  nnd2s1 U4980 ( .DIN1(n4075), .DIN2(n4076), .Q(\IDinst/n4887 ) );
  nnd2s1 U4981 ( .DIN1(n490), .DIN2(\IDinst/RegFile[21][31] ), .Q(n4076) );
  nnd2s1 U4982 ( .DIN1(n574), .DIN2(n4024), .Q(n4075) );
  nnd2s1 U4983 ( .DIN1(n4077), .DIN2(n4078), .Q(\IDinst/n4886 ) );
  nnd2s1 U4984 ( .DIN1(n504), .DIN2(\IDinst/RegFile[22][31] ), .Q(n4078) );
  nnd2s1 U4985 ( .DIN1(n576), .DIN2(n766), .Q(n4077) );
  nnd2s1 U4986 ( .DIN1(n4079), .DIN2(n4080), .Q(\IDinst/n4885 ) );
  nnd2s1 U4987 ( .DIN1(n480), .DIN2(\IDinst/RegFile[23][31] ), .Q(n4080) );
  nnd2s1 U4988 ( .DIN1(n578), .DIN2(n4024), .Q(n4079) );
  and3s1 U4989 ( .DIN1(\IDinst/n1430 ), .DIN2(n376), .DIN3(reg_write_MEM), 
        .Q(n4066) );
  nnd2s1 U4990 ( .DIN1(n4081), .DIN2(n4082), .Q(\IDinst/n4884 ) );
  nnd2s1 U4991 ( .DIN1(n472), .DIN2(\IDinst/RegFile[24][31] ), .Q(n4082) );
  nnd2s1 U4992 ( .DIN1(n564), .DIN2(n766), .Q(n4081) );
  and3s1 U4993 ( .DIN1(\IDinst/n1432 ), .DIN2(\IDinst/n1431 ), 
        .DIN3(\IDinst/n1433 ), .Q(n1383) );
  nnd2s1 U4994 ( .DIN1(n4084), .DIN2(n4085), .Q(\IDinst/n4883 ) );
  nnd2s1 U4995 ( .DIN1(n474), .DIN2(\IDinst/RegFile[25][31] ), .Q(n4085) );
  nnd2s1 U4996 ( .DIN1(n566), .DIN2(n4024), .Q(n4084) );
  and3s1 U4997 ( .DIN1(\IDinst/n1431 ), .DIN2(n27), .DIN3(\IDinst/n1432 ), 
        .Q(n4028) );
  nnd2s1 U4998 ( .DIN1(n4086), .DIN2(n4087), .Q(\IDinst/n4882 ) );
  nnd2s1 U4999 ( .DIN1(n468), .DIN2(\IDinst/RegFile[26][31] ), .Q(n4087) );
  nnd2s1 U5000 ( .DIN1(n568), .DIN2(n766), .Q(n4086) );
  and3s1 U5001 ( .DIN1(\IDinst/n1431 ), .DIN2(n58), .DIN3(\IDinst/n1433 ), 
        .Q(n4031) );
  nnd2s1 U5002 ( .DIN1(n4088), .DIN2(n4089), .Q(\IDinst/n4881 ) );
  nnd2s1 U5003 ( .DIN1(n470), .DIN2(\IDinst/RegFile[27][31] ), .Q(n4089) );
  nnd2s1 U5004 ( .DIN1(n570), .DIN2(n4024), .Q(n4088) );
  and3s1 U5005 ( .DIN1(n58), .DIN2(n27), .DIN3(\IDinst/n1431 ), .Q(n4034) );
  nnd2s1 U5006 ( .DIN1(n4090), .DIN2(n4091), .Q(\IDinst/n4880 ) );
  nnd2s1 U5007 ( .DIN1(n464), .DIN2(\IDinst/RegFile[28][31] ), .Q(n4091) );
  nnd2s1 U5008 ( .DIN1(n556), .DIN2(n766), .Q(n4090) );
  and3s1 U5009 ( .DIN1(\IDinst/n1432 ), .DIN2(n203), .DIN3(\IDinst/n1433 ), 
        .Q(n4037) );
  nnd2s1 U5010 ( .DIN1(n4092), .DIN2(n4093), .Q(\IDinst/n4879 ) );
  nnd2s1 U5011 ( .DIN1(n466), .DIN2(\IDinst/RegFile[29][31] ), .Q(n4093) );
  nnd2s1 U5012 ( .DIN1(n558), .DIN2(n4024), .Q(n4092) );
  and3s1 U5013 ( .DIN1(n203), .DIN2(n27), .DIN3(\IDinst/n1432 ), .Q(n4040) );
  nnd2s1 U5014 ( .DIN1(n4094), .DIN2(n4095), .Q(\IDinst/n4878 ) );
  nnd2s1 U5015 ( .DIN1(n460), .DIN2(\IDinst/RegFile[30][31] ), .Q(n4095) );
  nnd2s1 U5016 ( .DIN1(n560), .DIN2(n766), .Q(n4094) );
  and3s1 U5017 ( .DIN1(n203), .DIN2(n58), .DIN3(\IDinst/n1433 ), .Q(n4043) );
  nnd2s1 U5018 ( .DIN1(n4096), .DIN2(n4097), .Q(\IDinst/n4877 ) );
  nnd2s1 U5019 ( .DIN1(n462), .DIN2(\IDinst/RegFile[31][31] ), .Q(n4097) );
  nnd2s1 U5020 ( .DIN1(n562), .DIN2(n4024), .Q(n4096) );
  nnd2s1 U5021 ( .DIN1(n3035), .DIN2(n4098), .Q(n4024) );
  nnd2s1 U5022 ( .DIN1(n3103), .DIN2(n155), .Q(n4098) );
  nnd4s1 U5023 ( .DIN1(n3037), .DIN2(n379), .DIN3(n4099), .DIN4(n4100), 
        .Q(n3035) );
  or2s1 U5024 ( .DIN1(n129), .DIN2(n9405), .Q(n4100) );
  nnd2s1 U5025 ( .DIN1(n9404), .DIN2(n9405), .Q(n4099) );
  hi1s1 U5026 ( .DIN(n3103), .Q(n3037) );
  nnd4s1 U5027 ( .DIN1(n9400), .DIN2(n9401), .DIN3(n9402), .DIN4(n9403), 
        .Q(n3103) );
  and3s1 U5028 ( .DIN1(n376), .DIN2(n47), .DIN3(reg_write_MEM), .Q(n4083) );
  and3s1 U5029 ( .DIN1(n58), .DIN2(n27), .DIN3(n203), .Q(n4046) );
  nnd2s1 U5030 ( .DIN1(n4101), .DIN2(n4102), .Q(\IDinst/n4876 ) );
  nnd2s1 U5031 ( .DIN1(n396), .DIN2(n41), .Q(n4102) );
  nnd2s1 U5032 ( .DIN1(n651), .DIN2(n19), .Q(n4101) );
  nnd2s1 U5033 ( .DIN1(n4103), .DIN2(n4104), .Q(\IDinst/n4875 ) );
  nnd2s1 U5034 ( .DIN1(n396), .DIN2(n42), .Q(n4104) );
  nnd2s1 U5035 ( .DIN1(n650), .DIN2(n2), .Q(n4103) );
  nnd2s1 U5036 ( .DIN1(n4105), .DIN2(n4106), .Q(\IDinst/n4874 ) );
  nnd2s1 U5037 ( .DIN1(n396), .DIN2(n100), .Q(n4106) );
  nnd2s1 U5038 ( .DIN1(n649), .DIN2(n17), .Q(n4105) );
  nnd2s1 U5039 ( .DIN1(n4107), .DIN2(n4108), .Q(\IDinst/n4873 ) );
  nnd2s1 U5040 ( .DIN1(n396), .DIN2(n116), .Q(n4108) );
  nnd2s1 U5041 ( .DIN1(n652), .DIN2(n137), .Q(n4107) );
  nnd2s1 U5042 ( .DIN1(n4109), .DIN2(n4110), .Q(\IDinst/n4872 ) );
  nnd2s1 U5043 ( .DIN1(n396), .DIN2(n99), .Q(n4110) );
  or2s1 U5044 ( .DIN1(n130), .DIN2(n9416), .Q(n4109) );
  nnd3s1 U5045 ( .DIN1(n4111), .DIN2(n1964), .DIN3(n4112), .Q(\IDinst/n4871 )
         );
  nnd2s1 U5046 ( .DIN1(n651), .DIN2(n377), .Q(n4112) );
  nnd2s1 U5047 ( .DIN1(n1966), .DIN2(n115), .Q(n4111) );
  nnd2s1 U5048 ( .DIN1(n4113), .DIN2(n4114), .Q(\IDinst/n4870 ) );
  nnd4s1 U5049 ( .DIN1(n4115), .DIN2(n4116), .DIN3(n1927), .DIN4(n4117), 
        .Q(n4114) );
  or2s1 U5050 ( .DIN1(n130), .DIN2(n9414), .Q(n4113) );
  nnd2s1 U5051 ( .DIN1(n4118), .DIN2(n4119), .Q(\IDinst/n4869 ) );
  or2s1 U5052 ( .DIN1(n4120), .DIN2(n4121), .Q(n4119) );
  or2s1 U5053 ( .DIN1(n130), .DIN2(n9415), .Q(n4118) );
  nnd4s1 U5054 ( .DIN1(n4122), .DIN2(n4123), .DIN3(n1910), .DIN4(n1964), 
        .Q(\IDinst/n4868 ) );
  nnd3s1 U5055 ( .DIN1(n4120), .DIN2(n4124), .DIN3(n4115), .Q(n4123) );
  hi1s1 U5056 ( .DIN(n4121), .Q(n4115) );
  nnd2s1 U5057 ( .DIN1(reg_write), .DIN2(n650), .Q(n4122) );
  nnd4s1 U5058 ( .DIN1(n4125), .DIN2(n4126), .DIN3(n1910), .DIN4(n1964), 
        .Q(\IDinst/n4867 ) );
  hi1s1 U5059 ( .DIN(n529), .Q(n1964) );
  nnd2s1 U5060 ( .DIN1(n4127), .DIN2(n1966), .Q(n4126) );
  and2s1 U5061 ( .DIN1(n441), .DIN2(n4128), .Q(n1966) );
  hi1s1 U5062 ( .DIN(n4129), .Q(n4127) );
  nnd2s1 U5063 ( .DIN1(n650), .DIN2(reg_dst), .Q(n4125) );
  nnd2s1 U5064 ( .DIN1(n4130), .DIN2(n4131), .Q(\IDinst/n4866 ) );
  nnd4s1 U5065 ( .DIN1(n4116), .DIN2(n1927), .DIN3(n4117), .DIN4(n396), 
        .Q(n4131) );
  nnd2s1 U5066 ( .DIN1(n1953), .DIN2(n4132), .Q(n4117) );
  nnd2s1 U5067 ( .DIN1(n4133), .DIN2(n1950), .Q(n4132) );
  or2s1 U5068 ( .DIN1(n130), .DIN2(n9413), .Q(n4130) );
  nnd2s1 U5069 ( .DIN1(n4134), .DIN2(n4135), .Q(\IDinst/n4865 ) );
  nnd2s1 U5070 ( .DIN1(n1198), .DIN2(n396), .Q(n4135) );
  nnd2s1 U5071 ( .DIN1(n649), .DIN2(n229), .Q(n4134) );
  nnd2s1 U5072 ( .DIN1(n4136), .DIN2(n4137), .Q(\IDinst/n4864 ) );
  nnd2s1 U5073 ( .DIN1(n1312), .DIN2(n396), .Q(n4137) );
  nnd2s1 U5074 ( .DIN1(n652), .DIN2(n228), .Q(n4136) );
  nnd2s1 U5075 ( .DIN1(n4138), .DIN2(n4139), .Q(\IDinst/n4863 ) );
  nnd2s1 U5076 ( .DIN1(n1372), .DIN2(n396), .Q(n4139) );
  nnd2s1 U5077 ( .DIN1(n651), .DIN2(n227), .Q(n4138) );
  nnd2s1 U5078 ( .DIN1(n4140), .DIN2(n4141), .Q(\IDinst/n4862 ) );
  nnd2s1 U5079 ( .DIN1(n668), .DIN2(n396), .Q(n4141) );
  nnd2s1 U5080 ( .DIN1(n650), .DIN2(n49), .Q(n4140) );
  nnd2s1 U5081 ( .DIN1(n4142), .DIN2(n4143), .Q(\IDinst/n4861 ) );
  nnd2s1 U5082 ( .DIN1(\IDinst/N48 ), .DIN2(n396), .Q(n4143) );
  nnd2s1 U5083 ( .DIN1(n329), .DIN2(n4144), .Q(n4121) );
  nnd2s1 U5084 ( .DIN1(n649), .DIN2(n141), .Q(n4142) );
  nnd2s1 U5085 ( .DIN1(n4145), .DIN2(n4146), .Q(\IDinst/n4860 ) );
  nnd2s1 U5086 ( .DIN1(n4149), .DIN2(n4147), .Q(n4146) );
  nnd3s1 U5087 ( .DIN1(n4148), .DIN2(n1662), .DIN3(n777), .Q(n4145) );
  hi1s1 U5088 ( .DIN(n9459), .Q(n1662) );
  nnd2s1 U5089 ( .DIN1(n4150), .DIN2(n4151), .Q(\IDinst/n4859 ) );
  nnd2s1 U5090 ( .DIN1(n4152), .DIN2(n119), .Q(n4151) );
  nnd3s1 U5091 ( .DIN1(n4148), .DIN2(n4153), .DIN3(n4154), .Q(n4150) );
  nnd4s1 U5092 ( .DIN1(n4155), .DIN2(n4156), .DIN3(n676), .DIN4(n1910), 
        .Q(\IDinst/n4858 ) );
  or2s1 U5093 ( .DIN1(n4157), .DIN2(n383), .Q(n1910) );
  nnd3s1 U5094 ( .DIN1(\IDinst/slot_num[1]), .DIN2(n1919), .DIN3(n4152), 
        .Q(n4156) );
  nnd2s1 U5095 ( .DIN1(n441), .DIN2(n4153), .Q(n4155) );
  nnd2s1 U5096 ( .DIN1(n4158), .DIN2(n4159), .Q(n4153) );
  nnd2s1 U5097 ( .DIN1(n4160), .DIN2(n119), .Q(n4159) );
  nnd3s1 U5098 ( .DIN1(n4161), .DIN2(n1919), .DIN3(n4162), .Q(\IDinst/n4857 )
         );
  nnd2s1 U5099 ( .DIN1(n329), .DIN2(n4147), .Q(n4162) );
  nnd3s1 U5100 ( .DIN1(n4163), .DIN2(n4157), .DIN3(n4158), .Q(n4147) );
  and4s1 U5101 ( .DIN1(n4164), .DIN2(n4165), .DIN3(n4166), .DIN4(n4167), 
        .Q(n4158) );
  nnd2s1 U5102 ( .DIN1(n4168), .DIN2(n4169), .Q(n4165) );
  xnr2s1 U5103 ( .DIN1(n4170), .DIN2(n1950), .Q(n4169) );
  nnd2s1 U5104 ( .DIN1(n4171), .DIN2(n4172), .Q(n4170) );
  nor4s1 U5105 ( .DIN1(n4173), .DIN2(n4174), .DIN3(n4175), .DIN4(n4176), 
        .Q(n4172) );
  or4s1 U5106 ( .DIN1(n4177), .DIN2(n4178), .DIN3(n4179), .DIN4(n4180), 
        .Q(n4176) );
  or4s1 U5107 ( .DIN1(n4181), .DIN2(n4182), .DIN3(n4183), .DIN4(n4184), 
        .Q(n4175) );
  or4s1 U5108 ( .DIN1(n4185), .DIN2(n4186), .DIN3(n4187), .DIN4(n4188), 
        .Q(n4174) );
  or4s1 U5109 ( .DIN1(n4189), .DIN2(n4190), .DIN3(n4191), .DIN4(n4192), 
        .Q(n4173) );
  nor4s1 U5110 ( .DIN1(n4193), .DIN2(n4194), .DIN3(n4195), .DIN4(n4196), 
        .Q(n4171) );
  or4s1 U5111 ( .DIN1(n4197), .DIN2(n4198), .DIN3(n4199), .DIN4(n4200), 
        .Q(n4196) );
  or4s1 U5112 ( .DIN1(n4201), .DIN2(n4202), .DIN3(n4203), .DIN4(n4204), 
        .Q(n4195) );
  or4s1 U5113 ( .DIN1(n4205), .DIN2(n4206), .DIN3(n4207), .DIN4(n4208), 
        .Q(n4194) );
  or4s1 U5114 ( .DIN1(n4209), .DIN2(n4210), .DIN3(n4211), .DIN4(n4212), 
        .Q(n4193) );
  nnd3s1 U5115 ( .DIN1(n4213), .DIN2(n378), .DIN3(\IDinst/slot_num[1]), 
        .Q(n1919) );
  nnd2s1 U5116 ( .DIN1(\IDinst/n1445 ), .DIN2(\IDinst/n1440 ), .Q(n4213) );
  nnd3s1 U5117 ( .DIN1(\IDinst/slot_num[0]), .DIN2(n1915), .DIN3(n4152), 
        .Q(n4161) );
  hi1s1 U5118 ( .DIN(n4154), .Q(n4152) );
  nnd2s1 U5119 ( .DIN1(n383), .DIN2(n1914), .Q(n4154) );
  nnd3s1 U5120 ( .DIN1(n119), .DIN2(n60), .DIN3(\IDinst/slot_num[0]), 
        .Q(n1914) );
  nnd3s1 U5121 ( .DIN1(n215), .DIN2(n60), .DIN3(\IDinst/slot_num[0]), 
        .Q(n1915) );
  nnd2s1 U5122 ( .DIN1(n4214), .DIN2(n4215), .Q(\IDinst/n4856 ) );
  nnd2s1 U5123 ( .DIN1(n637), .DIN2(\IFinst/N7 ), .Q(n4215) );
  nnd2s1 U5124 ( .DIN1(n677), .DIN2(n154), .Q(n4214) );
  nnd2s1 U5125 ( .DIN1(n4216), .DIN2(n4217), .Q(\IDinst/n4855 ) );
  nnd2s1 U5126 ( .DIN1(n640), .DIN2(\IFinst/N8 ), .Q(n4217) );
  nnd2s1 U5127 ( .DIN1(n678), .DIN2(n153), .Q(n4216) );
  nnd2s1 U5128 ( .DIN1(n4218), .DIN2(n4219), .Q(\IDinst/n4854 ) );
  nnd2s1 U5129 ( .DIN1(n639), .DIN2(\NPC[2] ), .Q(n4219) );
  nnd2s1 U5130 ( .DIN1(n675), .DIN2(n152), .Q(n4218) );
  nnd2s1 U5131 ( .DIN1(n4220), .DIN2(n4221), .Q(\IDinst/n4853 ) );
  nnd2s1 U5132 ( .DIN1(n638), .DIN2(\NPC[3] ), .Q(n4221) );
  nnd2s1 U5133 ( .DIN1(n676), .DIN2(n151), .Q(n4220) );
  nnd2s1 U5134 ( .DIN1(n4222), .DIN2(n4223), .Q(\IDinst/n4852 ) );
  nnd2s1 U5135 ( .DIN1(n637), .DIN2(\NPC[4] ), .Q(n4223) );
  nnd2s1 U5136 ( .DIN1(n677), .DIN2(n150), .Q(n4222) );
  nnd2s1 U5137 ( .DIN1(n4224), .DIN2(n4225), .Q(\IDinst/n4851 ) );
  nnd2s1 U5138 ( .DIN1(n640), .DIN2(\NPC[5] ), .Q(n4225) );
  nnd2s1 U5139 ( .DIN1(n678), .DIN2(n149), .Q(n4224) );
  nnd2s1 U5140 ( .DIN1(n4226), .DIN2(n4227), .Q(\IDinst/n4850 ) );
  nnd2s1 U5141 ( .DIN1(n639), .DIN2(\NPC[6] ), .Q(n4227) );
  nnd2s1 U5142 ( .DIN1(n675), .DIN2(n148), .Q(n4226) );
  nnd2s1 U5143 ( .DIN1(n4228), .DIN2(n4229), .Q(\IDinst/n4849 ) );
  nnd2s1 U5144 ( .DIN1(n638), .DIN2(\NPC[7] ), .Q(n4229) );
  nnd2s1 U5145 ( .DIN1(n676), .DIN2(n147), .Q(n4228) );
  nnd2s1 U5146 ( .DIN1(n4230), .DIN2(n4231), .Q(\IDinst/n4848 ) );
  nnd2s1 U5147 ( .DIN1(n637), .DIN2(\NPC[8] ), .Q(n4231) );
  nnd2s1 U5148 ( .DIN1(n677), .DIN2(n201), .Q(n4230) );
  nnd2s1 U5149 ( .DIN1(n4232), .DIN2(n4233), .Q(\IDinst/n4847 ) );
  nnd2s1 U5150 ( .DIN1(n640), .DIN2(\NPC[9] ), .Q(n4233) );
  nnd2s1 U5151 ( .DIN1(n678), .DIN2(n199), .Q(n4232) );
  nnd2s1 U5152 ( .DIN1(n4234), .DIN2(n4235), .Q(\IDinst/n4846 ) );
  nnd2s1 U5153 ( .DIN1(n639), .DIN2(\NPC[10] ), .Q(n4235) );
  nnd2s1 U5154 ( .DIN1(n675), .DIN2(n197), .Q(n4234) );
  nnd2s1 U5155 ( .DIN1(n4236), .DIN2(n4237), .Q(\IDinst/n4845 ) );
  nnd2s1 U5156 ( .DIN1(n638), .DIN2(\NPC[11] ), .Q(n4237) );
  nnd2s1 U5157 ( .DIN1(n676), .DIN2(n195), .Q(n4236) );
  nnd2s1 U5158 ( .DIN1(n4238), .DIN2(n4239), .Q(\IDinst/n4844 ) );
  nnd2s1 U5159 ( .DIN1(n637), .DIN2(\NPC[12] ), .Q(n4239) );
  nnd2s1 U5160 ( .DIN1(n677), .DIN2(n193), .Q(n4238) );
  nnd2s1 U5161 ( .DIN1(n4240), .DIN2(n4241), .Q(\IDinst/n4843 ) );
  nnd2s1 U5162 ( .DIN1(n640), .DIN2(\NPC[13] ), .Q(n4241) );
  nnd2s1 U5163 ( .DIN1(n678), .DIN2(n191), .Q(n4240) );
  nnd2s1 U5164 ( .DIN1(n4242), .DIN2(n4243), .Q(\IDinst/n4842 ) );
  nnd2s1 U5165 ( .DIN1(n639), .DIN2(\NPC[14] ), .Q(n4243) );
  nnd2s1 U5166 ( .DIN1(n675), .DIN2(n189), .Q(n4242) );
  nnd2s1 U5167 ( .DIN1(n4244), .DIN2(n4245), .Q(\IDinst/n4841 ) );
  nnd2s1 U5168 ( .DIN1(n638), .DIN2(\NPC[15] ), .Q(n4245) );
  nnd2s1 U5169 ( .DIN1(n676), .DIN2(n187), .Q(n4244) );
  nnd2s1 U5170 ( .DIN1(n4246), .DIN2(n4247), .Q(\IDinst/n4840 ) );
  nnd2s1 U5171 ( .DIN1(n637), .DIN2(\NPC[16] ), .Q(n4247) );
  nnd2s1 U5172 ( .DIN1(n677), .DIN2(n186), .Q(n4246) );
  nnd2s1 U5173 ( .DIN1(n4248), .DIN2(n4249), .Q(\IDinst/n4839 ) );
  nnd2s1 U5174 ( .DIN1(n640), .DIN2(\NPC[17] ), .Q(n4249) );
  nnd2s1 U5175 ( .DIN1(n678), .DIN2(n184), .Q(n4248) );
  nnd2s1 U5176 ( .DIN1(n4250), .DIN2(n4251), .Q(\IDinst/n4838 ) );
  nnd2s1 U5177 ( .DIN1(n639), .DIN2(\NPC[18] ), .Q(n4251) );
  nnd2s1 U5178 ( .DIN1(n675), .DIN2(n182), .Q(n4250) );
  nnd2s1 U5179 ( .DIN1(n4252), .DIN2(n4253), .Q(\IDinst/n4837 ) );
  nnd2s1 U5180 ( .DIN1(n638), .DIN2(\NPC[19] ), .Q(n4253) );
  nnd2s1 U5181 ( .DIN1(n676), .DIN2(n180), .Q(n4252) );
  nnd2s1 U5182 ( .DIN1(n4254), .DIN2(n4255), .Q(\IDinst/n4836 ) );
  nnd2s1 U5183 ( .DIN1(n637), .DIN2(\NPC[20] ), .Q(n4255) );
  nnd2s1 U5184 ( .DIN1(n677), .DIN2(n178), .Q(n4254) );
  nnd2s1 U5185 ( .DIN1(n4256), .DIN2(n4257), .Q(\IDinst/n4835 ) );
  nnd2s1 U5186 ( .DIN1(n640), .DIN2(\NPC[21] ), .Q(n4257) );
  nnd2s1 U5187 ( .DIN1(n678), .DIN2(n176), .Q(n4256) );
  nnd2s1 U5188 ( .DIN1(n4258), .DIN2(n4259), .Q(\IDinst/n4834 ) );
  nnd2s1 U5189 ( .DIN1(n639), .DIN2(\NPC[22] ), .Q(n4259) );
  nnd2s1 U5190 ( .DIN1(n675), .DIN2(n174), .Q(n4258) );
  nnd2s1 U5191 ( .DIN1(n4260), .DIN2(n4261), .Q(\IDinst/n4833 ) );
  nnd2s1 U5192 ( .DIN1(n638), .DIN2(\NPC[23] ), .Q(n4261) );
  nnd2s1 U5193 ( .DIN1(n676), .DIN2(n172), .Q(n4260) );
  nnd2s1 U5194 ( .DIN1(n4262), .DIN2(n4263), .Q(\IDinst/n4832 ) );
  nnd2s1 U5195 ( .DIN1(n637), .DIN2(\NPC[24] ), .Q(n4263) );
  nnd2s1 U5196 ( .DIN1(n677), .DIN2(n170), .Q(n4262) );
  nnd2s1 U5197 ( .DIN1(n4264), .DIN2(n4265), .Q(\IDinst/n4831 ) );
  nnd2s1 U5198 ( .DIN1(n640), .DIN2(\NPC[25] ), .Q(n4265) );
  nnd2s1 U5199 ( .DIN1(n678), .DIN2(n168), .Q(n4264) );
  nnd2s1 U5200 ( .DIN1(n4266), .DIN2(n4267), .Q(\IDinst/n4830 ) );
  nnd2s1 U5201 ( .DIN1(n639), .DIN2(\NPC[26] ), .Q(n4267) );
  nnd2s1 U5202 ( .DIN1(n675), .DIN2(n166), .Q(n4266) );
  nnd2s1 U5203 ( .DIN1(n4268), .DIN2(n4269), .Q(\IDinst/n4829 ) );
  nnd2s1 U5204 ( .DIN1(n638), .DIN2(\NPC[27] ), .Q(n4269) );
  nnd2s1 U5205 ( .DIN1(n676), .DIN2(n164), .Q(n4268) );
  nnd2s1 U5206 ( .DIN1(n4270), .DIN2(n4271), .Q(\IDinst/n4828 ) );
  nnd2s1 U5207 ( .DIN1(n637), .DIN2(\NPC[28] ), .Q(n4271) );
  nnd2s1 U5208 ( .DIN1(n677), .DIN2(n162), .Q(n4270) );
  nnd2s1 U5209 ( .DIN1(n4272), .DIN2(n4273), .Q(\IDinst/n4827 ) );
  nnd2s1 U5210 ( .DIN1(n640), .DIN2(\NPC[29] ), .Q(n4273) );
  nnd2s1 U5211 ( .DIN1(n678), .DIN2(n160), .Q(n4272) );
  nnd2s1 U5212 ( .DIN1(n4274), .DIN2(n4275), .Q(\IDinst/n4826 ) );
  nnd2s1 U5213 ( .DIN1(n639), .DIN2(\NPC[30] ), .Q(n4275) );
  nnd2s1 U5214 ( .DIN1(n675), .DIN2(n158), .Q(n4274) );
  nnd2s1 U5215 ( .DIN1(n4276), .DIN2(n4277), .Q(\IDinst/n4825 ) );
  nnd2s1 U5216 ( .DIN1(n638), .DIN2(\NPC[31] ), .Q(n4277) );
  nnd2s1 U5217 ( .DIN1(n676), .DIN2(n156), .Q(n4276) );
  nnd4s1 U5218 ( .DIN1(n4278), .DIN2(n4279), .DIN3(n4280), .DIN4(n4281), 
        .Q(\IDinst/n4824 ) );
  nnd2s1 U5219 ( .DIN1(n4282), .DIN2(n781), .Q(n4281) );
  xnr2s1 U5220 ( .DIN1(n41), .DIN2(n9423), .Q(n4282) );
  nnd2s1 U5221 ( .DIN1(n751), .DIN2(n154), .Q(n4280) );
  nnd2s1 U5222 ( .DIN1(n756), .DIN2(n4204), .Q(n4279) );
  nnd2s1 U5223 ( .DIN1(n778), .DIN2(n233), .Q(n4278) );
  nnd4s1 U5224 ( .DIN1(n4286), .DIN2(n4287), .DIN3(n4288), .DIN4(n4289), 
        .Q(\IDinst/n4823 ) );
  nnd2s1 U5225 ( .DIN1(n4290), .DIN2(n781), .Q(n4289) );
  xor2s1 U5226 ( .DIN1(n4291), .DIN2(n4292), .Q(n4290) );
  xnr2s1 U5227 ( .DIN1(n42), .DIN2(n9422), .Q(n4292) );
  nor2s1 U5228 ( .DIN1(n9384), .DIN2(n9423), .Q(n4291) );
  nnd2s1 U5229 ( .DIN1(n750), .DIN2(n153), .Q(n4288) );
  nnd2s1 U5230 ( .DIN1(n757), .DIN2(n4203), .Q(n4287) );
  nnd2s1 U5231 ( .DIN1(n777), .DIN2(n234), .Q(n4286) );
  nnd4s1 U5232 ( .DIN1(n4293), .DIN2(n4294), .DIN3(n4295), .DIN4(n4296), 
        .Q(\IDinst/n4822 ) );
  nnd2s1 U5233 ( .DIN1(n751), .DIN2(n152), .Q(n4296) );
  nnd2s1 U5234 ( .DIN1(n756), .DIN2(n4202), .Q(n4295) );
  or2s1 U5235 ( .DIN1(n4297), .DIN2(n4298), .Q(n4294) );
  nnd2s1 U5236 ( .DIN1(n778), .DIN2(n235), .Q(n4293) );
  nnd4s1 U5237 ( .DIN1(n4299), .DIN2(n4300), .DIN3(n4301), .DIN4(n4302), 
        .Q(\IDinst/n4821 ) );
  nnd2s1 U5238 ( .DIN1(n781), .DIN2(n4303), .Q(n4302) );
  nnd2s1 U5239 ( .DIN1(n4304), .DIN2(n4305), .Q(n4303) );
  nnd2s1 U5240 ( .DIN1(n4306), .DIN2(n4297), .Q(n4305) );
  nnd2s1 U5241 ( .DIN1(n750), .DIN2(n151), .Q(n4301) );
  nnd2s1 U5242 ( .DIN1(n757), .DIN2(n4201), .Q(n4300) );
  nnd2s1 U5243 ( .DIN1(n777), .DIN2(n236), .Q(n4299) );
  nnd4s1 U5244 ( .DIN1(n4307), .DIN2(n4308), .DIN3(n4309), .DIN4(n4310), 
        .Q(\IDinst/n4820 ) );
  nnd2s1 U5245 ( .DIN1(n781), .DIN2(n4311), .Q(n4310) );
  nnd2s1 U5246 ( .DIN1(n4312), .DIN2(n4313), .Q(n4311) );
  nnd2s1 U5247 ( .DIN1(n4314), .DIN2(n4304), .Q(n4313) );
  nnd2s1 U5248 ( .DIN1(n751), .DIN2(n150), .Q(n4309) );
  nnd2s1 U5249 ( .DIN1(n756), .DIN2(n4200), .Q(n4308) );
  nnd2s1 U5250 ( .DIN1(n778), .DIN2(n237), .Q(n4307) );
  nnd4s1 U5251 ( .DIN1(n4315), .DIN2(n4316), .DIN3(n4317), .DIN4(n4318), 
        .Q(\IDinst/n4819 ) );
  nnd2s1 U5252 ( .DIN1(n781), .DIN2(n4319), .Q(n4318) );
  nnd2s1 U5253 ( .DIN1(n4320), .DIN2(n4321), .Q(n4319) );
  nnd2s1 U5254 ( .DIN1(n4322), .DIN2(n4312), .Q(n4321) );
  nnd2s1 U5255 ( .DIN1(n750), .DIN2(n149), .Q(n4317) );
  nnd2s1 U5256 ( .DIN1(n757), .DIN2(n4199), .Q(n4316) );
  nnd2s1 U5257 ( .DIN1(n777), .DIN2(n238), .Q(n4315) );
  nnd4s1 U5258 ( .DIN1(n4323), .DIN2(n4324), .DIN3(n4325), .DIN4(n4326), 
        .Q(\IDinst/n4818 ) );
  nnd2s1 U5259 ( .DIN1(n781), .DIN2(n4327), .Q(n4326) );
  nnd2s1 U5260 ( .DIN1(n4328), .DIN2(n4329), .Q(n4327) );
  nnd2s1 U5261 ( .DIN1(n4330), .DIN2(n4320), .Q(n4329) );
  hi1s1 U5262 ( .DIN(n4331), .Q(n4328) );
  nnd2s1 U5263 ( .DIN1(n751), .DIN2(n148), .Q(n4325) );
  nnd2s1 U5264 ( .DIN1(n756), .DIN2(n4198), .Q(n4324) );
  nnd2s1 U5265 ( .DIN1(n778), .DIN2(n239), .Q(n4323) );
  nnd4s1 U5266 ( .DIN1(n4332), .DIN2(n4333), .DIN3(n4334), .DIN4(n4335), 
        .Q(\IDinst/n4817 ) );
  nnd2s1 U5267 ( .DIN1(n750), .DIN2(n147), .Q(n4335) );
  nor2s1 U5268 ( .DIN1(n4336), .DIN2(n4337), .Q(n4334) );
  nor2s1 U5269 ( .DIN1(n4338), .DIN2(n4298), .Q(n4337) );
  nor2s1 U5270 ( .DIN1(n4339), .DIN2(n4340), .Q(n4338) );
  hi1s1 U5271 ( .DIN(n4341), .Q(n4340) );
  nor2s1 U5272 ( .DIN1(n4331), .DIN2(n4342), .Q(n4339) );
  nnd2s1 U5273 ( .DIN1(n757), .DIN2(n4197), .Q(n4333) );
  nnd2s1 U5274 ( .DIN1(n777), .DIN2(n240), .Q(n4332) );
  nnd4s1 U5275 ( .DIN1(n4343), .DIN2(n4344), .DIN3(n4345), .DIN4(n4346), 
        .Q(\IDinst/n4816 ) );
  nnd2s1 U5276 ( .DIN1(n781), .DIN2(n4347), .Q(n4346) );
  nnd2s1 U5277 ( .DIN1(n4348), .DIN2(n4349), .Q(n4347) );
  nnd2s1 U5278 ( .DIN1(n4350), .DIN2(n4341), .Q(n4349) );
  nnd2s1 U5279 ( .DIN1(n751), .DIN2(n201), .Q(n4345) );
  nnd2s1 U5280 ( .DIN1(n756), .DIN2(n4192), .Q(n4344) );
  nnd2s1 U5281 ( .DIN1(n778), .DIN2(n241), .Q(n4343) );
  nnd4s1 U5282 ( .DIN1(n4351), .DIN2(n4352), .DIN3(n4353), .DIN4(n4354), 
        .Q(\IDinst/n4815 ) );
  nnd2s1 U5283 ( .DIN1(n781), .DIN2(n4355), .Q(n4354) );
  nnd2s1 U5284 ( .DIN1(n4356), .DIN2(n4357), .Q(n4355) );
  nnd2s1 U5285 ( .DIN1(n4358), .DIN2(n4348), .Q(n4357) );
  nnd2s1 U5286 ( .DIN1(n750), .DIN2(n199), .Q(n4353) );
  nnd2s1 U5287 ( .DIN1(n757), .DIN2(n4191), .Q(n4352) );
  nnd2s1 U5288 ( .DIN1(n777), .DIN2(n242), .Q(n4351) );
  nnd4s1 U5289 ( .DIN1(n4359), .DIN2(n4360), .DIN3(n4361), .DIN4(n4362), 
        .Q(\IDinst/n4814 ) );
  nnd2s1 U5290 ( .DIN1(n781), .DIN2(n4363), .Q(n4362) );
  nnd2s1 U5291 ( .DIN1(n4364), .DIN2(n4365), .Q(n4363) );
  nnd2s1 U5292 ( .DIN1(n4366), .DIN2(n4356), .Q(n4365) );
  nnd2s1 U5293 ( .DIN1(n751), .DIN2(n197), .Q(n4361) );
  nnd2s1 U5294 ( .DIN1(n756), .DIN2(n4190), .Q(n4360) );
  nnd2s1 U5295 ( .DIN1(n778), .DIN2(n243), .Q(n4359) );
  nnd4s1 U5296 ( .DIN1(n4367), .DIN2(n4368), .DIN3(n4369), .DIN4(n4370), 
        .Q(\IDinst/n4813 ) );
  nnd2s1 U5297 ( .DIN1(n781), .DIN2(n4371), .Q(n4370) );
  nnd2s1 U5298 ( .DIN1(n4372), .DIN2(n4373), .Q(n4371) );
  nnd2s1 U5299 ( .DIN1(n4374), .DIN2(n4364), .Q(n4373) );
  nnd2s1 U5300 ( .DIN1(n750), .DIN2(n195), .Q(n4369) );
  nnd2s1 U5301 ( .DIN1(n757), .DIN2(n4189), .Q(n4368) );
  nnd2s1 U5302 ( .DIN1(n777), .DIN2(n244), .Q(n4367) );
  nnd4s1 U5303 ( .DIN1(n4375), .DIN2(n4376), .DIN3(n4377), .DIN4(n4378), 
        .Q(\IDinst/n4812 ) );
  nnd2s1 U5304 ( .DIN1(n781), .DIN2(n4379), .Q(n4378) );
  nnd2s1 U5305 ( .DIN1(n4380), .DIN2(n4381), .Q(n4379) );
  nnd2s1 U5306 ( .DIN1(n4382), .DIN2(n4372), .Q(n4381) );
  nnd2s1 U5307 ( .DIN1(n751), .DIN2(n193), .Q(n4377) );
  nnd2s1 U5308 ( .DIN1(n756), .DIN2(n4188), .Q(n4376) );
  nnd2s1 U5309 ( .DIN1(n778), .DIN2(n245), .Q(n4375) );
  nnd4s1 U5310 ( .DIN1(n4383), .DIN2(n4384), .DIN3(n4385), .DIN4(n4386), 
        .Q(\IDinst/n4811 ) );
  nnd2s1 U5311 ( .DIN1(n781), .DIN2(n4387), .Q(n4386) );
  nnd2s1 U5312 ( .DIN1(n4388), .DIN2(n4389), .Q(n4387) );
  nnd2s1 U5313 ( .DIN1(n4390), .DIN2(n4380), .Q(n4389) );
  nnd2s1 U5314 ( .DIN1(n750), .DIN2(n191), .Q(n4385) );
  nnd2s1 U5315 ( .DIN1(n757), .DIN2(n4187), .Q(n4384) );
  nnd2s1 U5316 ( .DIN1(n777), .DIN2(n246), .Q(n4383) );
  nnd4s1 U5317 ( .DIN1(n4391), .DIN2(n4392), .DIN3(n4393), .DIN4(n4394), 
        .Q(\IDinst/n4810 ) );
  nnd2s1 U5318 ( .DIN1(n4283), .DIN2(n4395), .Q(n4394) );
  nnd2s1 U5319 ( .DIN1(n4396), .DIN2(n4397), .Q(n4395) );
  nnd2s1 U5320 ( .DIN1(n4398), .DIN2(n4388), .Q(n4397) );
  nnd2s1 U5321 ( .DIN1(n751), .DIN2(n189), .Q(n4393) );
  nnd2s1 U5322 ( .DIN1(n756), .DIN2(n4186), .Q(n4392) );
  nnd2s1 U5323 ( .DIN1(n778), .DIN2(n247), .Q(n4391) );
  nnd4s1 U5324 ( .DIN1(n4399), .DIN2(n4400), .DIN3(n4401), .DIN4(n4402), 
        .Q(\IDinst/n4809 ) );
  nnd2s1 U5325 ( .DIN1(n4283), .DIN2(n4403), .Q(n4402) );
  nnd2s1 U5326 ( .DIN1(n4404), .DIN2(n4405), .Q(n4403) );
  nnd2s1 U5327 ( .DIN1(n4406), .DIN2(n4396), .Q(n4405) );
  nnd2s1 U5328 ( .DIN1(n750), .DIN2(n187), .Q(n4401) );
  nnd2s1 U5329 ( .DIN1(n757), .DIN2(n4185), .Q(n4400) );
  nnd2s1 U5330 ( .DIN1(n777), .DIN2(n248), .Q(n4399) );
  nnd4s1 U5331 ( .DIN1(n4407), .DIN2(n4408), .DIN3(n4409), .DIN4(n4410), 
        .Q(\IDinst/n4808 ) );
  nnd2s1 U5332 ( .DIN1(n4283), .DIN2(n4411), .Q(n4410) );
  nnd2s1 U5333 ( .DIN1(n4412), .DIN2(n4413), .Q(n4411) );
  nnd2s1 U5334 ( .DIN1(n4414), .DIN2(n4404), .Q(n4413) );
  nnd2s1 U5335 ( .DIN1(n751), .DIN2(n186), .Q(n4409) );
  nnd2s1 U5336 ( .DIN1(n756), .DIN2(n4184), .Q(n4408) );
  nnd2s1 U5337 ( .DIN1(n778), .DIN2(n249), .Q(n4407) );
  nnd4s1 U5338 ( .DIN1(n4415), .DIN2(n4416), .DIN3(n4417), .DIN4(n4418), 
        .Q(\IDinst/n4807 ) );
  nnd2s1 U5339 ( .DIN1(n4283), .DIN2(n4419), .Q(n4418) );
  nnd2s1 U5340 ( .DIN1(n4420), .DIN2(n4421), .Q(n4419) );
  nnd2s1 U5341 ( .DIN1(n4422), .DIN2(n4412), .Q(n4421) );
  nnd2s1 U5342 ( .DIN1(n750), .DIN2(n184), .Q(n4417) );
  nnd2s1 U5343 ( .DIN1(n757), .DIN2(n4183), .Q(n4416) );
  nnd2s1 U5344 ( .DIN1(n777), .DIN2(n250), .Q(n4415) );
  nnd4s1 U5345 ( .DIN1(n4423), .DIN2(n4424), .DIN3(n4425), .DIN4(n4426), 
        .Q(\IDinst/n4806 ) );
  nnd2s1 U5346 ( .DIN1(n4283), .DIN2(n4427), .Q(n4426) );
  nnd2s1 U5347 ( .DIN1(n4428), .DIN2(n4429), .Q(n4427) );
  nnd2s1 U5348 ( .DIN1(n4430), .DIN2(n4420), .Q(n4429) );
  nnd2s1 U5349 ( .DIN1(n751), .DIN2(n182), .Q(n4425) );
  nnd2s1 U5350 ( .DIN1(n756), .DIN2(n4182), .Q(n4424) );
  nnd2s1 U5351 ( .DIN1(n778), .DIN2(n251), .Q(n4423) );
  nnd4s1 U5352 ( .DIN1(n4431), .DIN2(n4432), .DIN3(n4433), .DIN4(n4434), 
        .Q(\IDinst/n4805 ) );
  nnd2s1 U5353 ( .DIN1(n4283), .DIN2(n4435), .Q(n4434) );
  nnd2s1 U5354 ( .DIN1(n4436), .DIN2(n4437), .Q(n4435) );
  nnd2s1 U5355 ( .DIN1(n4438), .DIN2(n4428), .Q(n4437) );
  nnd2s1 U5356 ( .DIN1(n750), .DIN2(n180), .Q(n4433) );
  nnd2s1 U5357 ( .DIN1(n757), .DIN2(n4181), .Q(n4432) );
  nnd2s1 U5358 ( .DIN1(n777), .DIN2(n252), .Q(n4431) );
  nnd4s1 U5359 ( .DIN1(n4439), .DIN2(n4440), .DIN3(n4441), .DIN4(n4442), 
        .Q(\IDinst/n4804 ) );
  nnd2s1 U5360 ( .DIN1(n4283), .DIN2(n4443), .Q(n4442) );
  nnd2s1 U5361 ( .DIN1(n4444), .DIN2(n4445), .Q(n4443) );
  nnd2s1 U5362 ( .DIN1(n4446), .DIN2(n4436), .Q(n4445) );
  nnd2s1 U5363 ( .DIN1(n751), .DIN2(n178), .Q(n4441) );
  nnd2s1 U5364 ( .DIN1(n756), .DIN2(n4180), .Q(n4440) );
  nnd2s1 U5365 ( .DIN1(n778), .DIN2(n253), .Q(n4439) );
  nnd4s1 U5366 ( .DIN1(n4447), .DIN2(n4448), .DIN3(n4449), .DIN4(n4450), 
        .Q(\IDinst/n4803 ) );
  nnd2s1 U5367 ( .DIN1(n4283), .DIN2(n4451), .Q(n4450) );
  nnd2s1 U5368 ( .DIN1(n4452), .DIN2(n4453), .Q(n4451) );
  nnd2s1 U5369 ( .DIN1(n4454), .DIN2(n4444), .Q(n4453) );
  nnd2s1 U5370 ( .DIN1(n750), .DIN2(n176), .Q(n4449) );
  nnd2s1 U5371 ( .DIN1(n757), .DIN2(n4179), .Q(n4448) );
  nnd2s1 U5372 ( .DIN1(n777), .DIN2(n254), .Q(n4447) );
  nnd4s1 U5373 ( .DIN1(n4455), .DIN2(n4456), .DIN3(n4457), .DIN4(n4458), 
        .Q(\IDinst/n4802 ) );
  nnd2s1 U5374 ( .DIN1(n4283), .DIN2(n4459), .Q(n4458) );
  nnd2s1 U5375 ( .DIN1(n4460), .DIN2(n4461), .Q(n4459) );
  nnd2s1 U5376 ( .DIN1(n4462), .DIN2(n4452), .Q(n4461) );
  nnd2s1 U5377 ( .DIN1(n751), .DIN2(n174), .Q(n4457) );
  nnd2s1 U5378 ( .DIN1(n756), .DIN2(n4178), .Q(n4456) );
  nnd2s1 U5379 ( .DIN1(n778), .DIN2(n255), .Q(n4455) );
  nnd4s1 U5380 ( .DIN1(n4463), .DIN2(n4464), .DIN3(n4465), .DIN4(n4466), 
        .Q(\IDinst/n4801 ) );
  nnd2s1 U5381 ( .DIN1(n4283), .DIN2(n4467), .Q(n4466) );
  nnd2s1 U5382 ( .DIN1(n4468), .DIN2(n4469), .Q(n4467) );
  nnd2s1 U5383 ( .DIN1(n4470), .DIN2(n4460), .Q(n4469) );
  nnd2s1 U5384 ( .DIN1(n750), .DIN2(n172), .Q(n4465) );
  nnd2s1 U5385 ( .DIN1(n757), .DIN2(n4177), .Q(n4464) );
  nnd2s1 U5386 ( .DIN1(n777), .DIN2(n256), .Q(n4463) );
  nnd4s1 U5387 ( .DIN1(n4471), .DIN2(n4472), .DIN3(n4473), .DIN4(n4474), 
        .Q(\IDinst/n4800 ) );
  nnd2s1 U5388 ( .DIN1(n4283), .DIN2(n4475), .Q(n4474) );
  nnd2s1 U5389 ( .DIN1(n4476), .DIN2(n4477), .Q(n4475) );
  nnd2s1 U5390 ( .DIN1(n4478), .DIN2(n4468), .Q(n4477) );
  nnd2s1 U5391 ( .DIN1(n751), .DIN2(n170), .Q(n4473) );
  nnd2s1 U5392 ( .DIN1(n756), .DIN2(n4212), .Q(n4472) );
  nnd2s1 U5393 ( .DIN1(n778), .DIN2(n257), .Q(n4471) );
  nnd4s1 U5394 ( .DIN1(n4479), .DIN2(n4480), .DIN3(n4481), .DIN4(n4482), 
        .Q(\IDinst/n4799 ) );
  nnd2s1 U5395 ( .DIN1(n4283), .DIN2(n4483), .Q(n4482) );
  nnd2s1 U5396 ( .DIN1(n4484), .DIN2(n4485), .Q(n4483) );
  nnd2s1 U5397 ( .DIN1(n4486), .DIN2(n4476), .Q(n4485) );
  nnd2s1 U5398 ( .DIN1(n750), .DIN2(n168), .Q(n4481) );
  nnd2s1 U5399 ( .DIN1(n757), .DIN2(n4211), .Q(n4480) );
  nnd2s1 U5400 ( .DIN1(n777), .DIN2(n258), .Q(n4479) );
  nnd4s1 U5401 ( .DIN1(n4487), .DIN2(n4488), .DIN3(n4489), .DIN4(n4490), 
        .Q(\IDinst/n4798 ) );
  nnd2s1 U5402 ( .DIN1(n4283), .DIN2(n4491), .Q(n4490) );
  nnd2s1 U5403 ( .DIN1(n4492), .DIN2(n4493), .Q(n4491) );
  nnd2s1 U5404 ( .DIN1(n4494), .DIN2(n4484), .Q(n4493) );
  nnd2s1 U5405 ( .DIN1(n751), .DIN2(n166), .Q(n4489) );
  nnd2s1 U5406 ( .DIN1(n756), .DIN2(n4210), .Q(n4488) );
  nnd2s1 U5407 ( .DIN1(n778), .DIN2(n259), .Q(n4487) );
  nnd4s1 U5408 ( .DIN1(n4495), .DIN2(n4496), .DIN3(n4497), .DIN4(n4498), 
        .Q(\IDinst/n4797 ) );
  nnd2s1 U5409 ( .DIN1(n4283), .DIN2(n4499), .Q(n4498) );
  nnd2s1 U5410 ( .DIN1(n4500), .DIN2(n4501), .Q(n4499) );
  nnd2s1 U5411 ( .DIN1(n4502), .DIN2(n4492), .Q(n4501) );
  nnd2s1 U5412 ( .DIN1(n750), .DIN2(n164), .Q(n4497) );
  nnd2s1 U5413 ( .DIN1(n757), .DIN2(n4209), .Q(n4496) );
  nnd2s1 U5414 ( .DIN1(n777), .DIN2(n260), .Q(n4495) );
  nnd4s1 U5415 ( .DIN1(n4503), .DIN2(n4504), .DIN3(n4505), .DIN4(n4506), 
        .Q(\IDinst/n4796 ) );
  nnd2s1 U5416 ( .DIN1(n4283), .DIN2(n4507), .Q(n4506) );
  nnd2s1 U5417 ( .DIN1(n4508), .DIN2(n4509), .Q(n4507) );
  nnd2s1 U5418 ( .DIN1(n4510), .DIN2(n4500), .Q(n4509) );
  nnd2s1 U5419 ( .DIN1(n751), .DIN2(n162), .Q(n4505) );
  nnd2s1 U5420 ( .DIN1(n756), .DIN2(n4208), .Q(n4504) );
  nnd2s1 U5421 ( .DIN1(n778), .DIN2(n261), .Q(n4503) );
  nnd4s1 U5422 ( .DIN1(n4511), .DIN2(n4512), .DIN3(n4513), .DIN4(n4514), 
        .Q(\IDinst/n4795 ) );
  nnd2s1 U5423 ( .DIN1(n4283), .DIN2(n4515), .Q(n4514) );
  nnd2s1 U5424 ( .DIN1(n4516), .DIN2(n4517), .Q(n4515) );
  nnd2s1 U5425 ( .DIN1(n4518), .DIN2(n4508), .Q(n4517) );
  hi1s1 U5426 ( .DIN(n4519), .Q(n4516) );
  nnd2s1 U5427 ( .DIN1(n750), .DIN2(n160), .Q(n4513) );
  nnd2s1 U5428 ( .DIN1(n757), .DIN2(n4207), .Q(n4512) );
  nnd2s1 U5429 ( .DIN1(n777), .DIN2(n262), .Q(n4511) );
  nnd4s1 U5430 ( .DIN1(n4520), .DIN2(n4521), .DIN3(n4522), .DIN4(n4523), 
        .Q(\IDinst/n4794 ) );
  nnd2s1 U5431 ( .DIN1(n4283), .DIN2(n4524), .Q(n4523) );
  nnd2s1 U5432 ( .DIN1(n4525), .DIN2(n4526), .Q(n4524) );
  or2s1 U5433 ( .DIN1(n4527), .DIN2(n4519), .Q(n4526) );
  nnd2s1 U5434 ( .DIN1(n751), .DIN2(n158), .Q(n4522) );
  nnd2s1 U5435 ( .DIN1(n756), .DIN2(n4206), .Q(n4521) );
  nnd2s1 U5436 ( .DIN1(n778), .DIN2(n263), .Q(n4520) );
  nnd4s1 U5437 ( .DIN1(n4528), .DIN2(n4529), .DIN3(n4530), .DIN4(n4531), 
        .Q(\IDinst/n4793 ) );
  nor2s1 U5438 ( .DIN1(n4532), .DIN2(n4533), .Q(n4531) );
  nor2s1 U5439 ( .DIN1(n9406), .DIN2(n4149), .Q(n4533) );
  and2s1 U5440 ( .DIN1(n4205), .DIN2(n757), .Q(n4532) );
  nnd2s1 U5441 ( .DIN1(n750), .DIN2(n156), .Q(n4530) );
  hi1s1 U5442 ( .DIN(n4336), .Q(n4529) );
  nor2s1 U5443 ( .DIN1(n777), .DIN2(n4535), .Q(n4336) );
  nnd2s1 U5444 ( .DIN1(n4283), .DIN2(n4536), .Q(n4528) );
  xor2s1 U5445 ( .DIN1(n4537), .DIN2(n4538), .Q(n4536) );
  xor2s1 U5446 ( .DIN1(n4525), .DIN2(n4539), .Q(n4538) );
  nnd2s1 U5447 ( .DIN1(n4540), .DIN2(n4541), .Q(n4539) );
  nnd2s1 U5448 ( .DIN1(n9520), .DIN2(n4542), .Q(n4541) );
  nnd2s1 U5449 ( .DIN1(n4543), .DIN2(n4544), .Q(n4542) );
  or2s1 U5450 ( .DIN1(n4544), .DIN2(n732), .Q(n4540) );
  nnd2s1 U5451 ( .DIN1(n4519), .DIN2(n4527), .Q(n4525) );
  xnr2s1 U5452 ( .DIN1(n4544), .DIN2(n4545), .Q(n4527) );
  xnr2s1 U5453 ( .DIN1(n9520), .DIN2(n4543), .Q(n4545) );
  nnd2s1 U5454 ( .DIN1(n4546), .DIN2(n4547), .Q(n4544) );
  nnd2s1 U5455 ( .DIN1(n4548), .DIN2(\NPC[29] ), .Q(n4547) );
  or2s1 U5456 ( .DIN1(n4549), .DIN2(n732), .Q(n4548) );
  nnd2s1 U5457 ( .DIN1(n4549), .DIN2(n732), .Q(n4546) );
  nor2s1 U5458 ( .DIN1(n4508), .DIN2(n4518), .Q(n4519) );
  xnr2s1 U5459 ( .DIN1(n4550), .DIN2(n4549), .Q(n4518) );
  nnd2s1 U5460 ( .DIN1(n4551), .DIN2(n4552), .Q(n4549) );
  nnd2s1 U5461 ( .DIN1(n4553), .DIN2(\NPC[28] ), .Q(n4552) );
  or2s1 U5462 ( .DIN1(n4554), .DIN2(n732), .Q(n4553) );
  nnd2s1 U5463 ( .DIN1(n4554), .DIN2(n732), .Q(n4551) );
  xnr2s1 U5464 ( .DIN1(n9425), .DIN2(n4555), .Q(n4550) );
  or2s1 U5465 ( .DIN1(n4500), .DIN2(n4510), .Q(n4508) );
  xor2s1 U5466 ( .DIN1(n4554), .DIN2(n4556), .Q(n4510) );
  xnr2s1 U5467 ( .DIN1(n9426), .DIN2(n4543), .Q(n4556) );
  nnd2s1 U5468 ( .DIN1(n4557), .DIN2(n4558), .Q(n4554) );
  nnd2s1 U5469 ( .DIN1(n4559), .DIN2(\NPC[27] ), .Q(n4558) );
  or2s1 U5470 ( .DIN1(n4560), .DIN2(n732), .Q(n4559) );
  nnd2s1 U5471 ( .DIN1(n4560), .DIN2(n4543), .Q(n4557) );
  or2s1 U5472 ( .DIN1(n4492), .DIN2(n4502), .Q(n4500) );
  xnr2s1 U5473 ( .DIN1(n4561), .DIN2(n4560), .Q(n4502) );
  nnd2s1 U5474 ( .DIN1(n4562), .DIN2(n4563), .Q(n4560) );
  nnd2s1 U5475 ( .DIN1(n4564), .DIN2(\NPC[26] ), .Q(n4563) );
  or2s1 U5476 ( .DIN1(n4565), .DIN2(n732), .Q(n4564) );
  nnd2s1 U5477 ( .DIN1(n4565), .DIN2(n4543), .Q(n4562) );
  xnr2s1 U5478 ( .DIN1(n9427), .DIN2(n4555), .Q(n4561) );
  or2s1 U5479 ( .DIN1(n4484), .DIN2(n4494), .Q(n4492) );
  xor2s1 U5480 ( .DIN1(n4565), .DIN2(n4566), .Q(n4494) );
  xnr2s1 U5481 ( .DIN1(n9428), .DIN2(n4543), .Q(n4566) );
  nnd2s1 U5482 ( .DIN1(n4567), .DIN2(n4568), .Q(n4565) );
  nnd2s1 U5483 ( .DIN1(n4569), .DIN2(\NPC[25] ), .Q(n4568) );
  or2s1 U5484 ( .DIN1(n4570), .DIN2(n732), .Q(n4569) );
  nnd2s1 U5485 ( .DIN1(n4570), .DIN2(n4543), .Q(n4567) );
  or2s1 U5486 ( .DIN1(n4476), .DIN2(n4486), .Q(n4484) );
  xnr2s1 U5487 ( .DIN1(n4571), .DIN2(n4570), .Q(n4486) );
  nnd2s1 U5488 ( .DIN1(n4572), .DIN2(n4573), .Q(n4570) );
  nnd2s1 U5489 ( .DIN1(n4574), .DIN2(\NPC[24] ), .Q(n4573) );
  or2s1 U5490 ( .DIN1(n4575), .DIN2(n4576), .Q(n4574) );
  nnd2s1 U5491 ( .DIN1(n4575), .DIN2(n4576), .Q(n4572) );
  xnr2s1 U5492 ( .DIN1(n9429), .DIN2(n4555), .Q(n4571) );
  hi1s1 U5493 ( .DIN(n4543), .Q(n4555) );
  or2s1 U5494 ( .DIN1(n4468), .DIN2(n4478), .Q(n4476) );
  xor2s1 U5495 ( .DIN1(n4575), .DIN2(n4577), .Q(n4478) );
  xnr2s1 U5496 ( .DIN1(n9430), .DIN2(n4576), .Q(n4577) );
  nnd2s1 U5497 ( .DIN1(n4578), .DIN2(n4579), .Q(n4576) );
  nnd2s1 U5498 ( .DIN1(n4580), .DIN2(\NPC[23] ), .Q(n4579) );
  or2s1 U5499 ( .DIN1(n4581), .DIN2(n4582), .Q(n4580) );
  nnd2s1 U5500 ( .DIN1(n4581), .DIN2(n4582), .Q(n4578) );
  nnd2s1 U5501 ( .DIN1(n4583), .DIN2(n4584), .Q(n4575) );
  nnd2s1 U5502 ( .DIN1(n643), .DIN2(n4585), .Q(n4584) );
  or2s1 U5503 ( .DIN1(n4460), .DIN2(n4470), .Q(n4468) );
  xor2s1 U5504 ( .DIN1(n4581), .DIN2(n4586), .Q(n4470) );
  xnr2s1 U5505 ( .DIN1(n9431), .DIN2(n4582), .Q(n4586) );
  nnd2s1 U5506 ( .DIN1(n4587), .DIN2(n4588), .Q(n4582) );
  nnd2s1 U5507 ( .DIN1(n4589), .DIN2(\NPC[22] ), .Q(n4588) );
  or2s1 U5508 ( .DIN1(n4590), .DIN2(n4591), .Q(n4589) );
  nnd2s1 U5509 ( .DIN1(n4590), .DIN2(n4591), .Q(n4587) );
  nnd2s1 U5510 ( .DIN1(n4583), .DIN2(n4592), .Q(n4581) );
  nnd2s1 U5511 ( .DIN1(n1197), .DIN2(n4585), .Q(n4592) );
  or2s1 U5512 ( .DIN1(n4452), .DIN2(n4462), .Q(n4460) );
  xor2s1 U5513 ( .DIN1(n4590), .DIN2(n4593), .Q(n4462) );
  xnr2s1 U5514 ( .DIN1(n9432), .DIN2(n4591), .Q(n4593) );
  nnd2s1 U5515 ( .DIN1(n4594), .DIN2(n4595), .Q(n4591) );
  nnd2s1 U5516 ( .DIN1(n4596), .DIN2(\NPC[21] ), .Q(n4595) );
  or2s1 U5517 ( .DIN1(n4597), .DIN2(n4598), .Q(n4596) );
  nnd2s1 U5518 ( .DIN1(n4597), .DIN2(n4598), .Q(n4594) );
  nnd2s1 U5519 ( .DIN1(n4583), .DIN2(n4599), .Q(n4590) );
  nnd2s1 U5520 ( .DIN1(n1153), .DIN2(n4585), .Q(n4599) );
  or2s1 U5521 ( .DIN1(n4444), .DIN2(n4454), .Q(n4452) );
  xor2s1 U5522 ( .DIN1(n4597), .DIN2(n4600), .Q(n4454) );
  xnr2s1 U5523 ( .DIN1(n9433), .DIN2(n4598), .Q(n4600) );
  nnd2s1 U5524 ( .DIN1(n4601), .DIN2(n4602), .Q(n4598) );
  nnd2s1 U5525 ( .DIN1(n4603), .DIN2(\NPC[20] ), .Q(n4602) );
  or2s1 U5526 ( .DIN1(n4604), .DIN2(n4605), .Q(n4603) );
  nnd2s1 U5527 ( .DIN1(n4604), .DIN2(n4605), .Q(n4601) );
  nnd2s1 U5528 ( .DIN1(n4583), .DIN2(n4606), .Q(n4597) );
  nnd2s1 U5529 ( .DIN1(n1065), .DIN2(n4585), .Q(n4606) );
  or2s1 U5530 ( .DIN1(n4436), .DIN2(n4446), .Q(n4444) );
  xor2s1 U5531 ( .DIN1(n4604), .DIN2(n4607), .Q(n4446) );
  xnr2s1 U5532 ( .DIN1(n9434), .DIN2(n4605), .Q(n4607) );
  nnd2s1 U5533 ( .DIN1(n4608), .DIN2(n4609), .Q(n4605) );
  nnd2s1 U5534 ( .DIN1(n4610), .DIN2(\NPC[19] ), .Q(n4609) );
  or2s1 U5535 ( .DIN1(n4611), .DIN2(n4612), .Q(n4610) );
  nnd2s1 U5536 ( .DIN1(n4611), .DIN2(n4612), .Q(n4608) );
  nnd2s1 U5537 ( .DIN1(n4583), .DIN2(n4613), .Q(n4604) );
  nnd2s1 U5538 ( .DIN1(n534), .DIN2(n4585), .Q(n4613) );
  or2s1 U5539 ( .DIN1(n4428), .DIN2(n4438), .Q(n4436) );
  xor2s1 U5540 ( .DIN1(n4611), .DIN2(n4614), .Q(n4438) );
  xnr2s1 U5541 ( .DIN1(n9435), .DIN2(n4612), .Q(n4614) );
  nnd2s1 U5542 ( .DIN1(n4615), .DIN2(n4616), .Q(n4612) );
  nnd2s1 U5543 ( .DIN1(n4617), .DIN2(\NPC[18] ), .Q(n4616) );
  or2s1 U5544 ( .DIN1(n4618), .DIN2(n4619), .Q(n4617) );
  nnd2s1 U5545 ( .DIN1(n4618), .DIN2(n4619), .Q(n4615) );
  nnd2s1 U5546 ( .DIN1(n4583), .DIN2(n4620), .Q(n4611) );
  nnd2s1 U5547 ( .DIN1(n665), .DIN2(n4585), .Q(n4620) );
  or2s1 U5548 ( .DIN1(n4420), .DIN2(n4430), .Q(n4428) );
  xor2s1 U5549 ( .DIN1(n4618), .DIN2(n4621), .Q(n4430) );
  xnr2s1 U5550 ( .DIN1(n9436), .DIN2(n4619), .Q(n4621) );
  nnd2s1 U5551 ( .DIN1(n4622), .DIN2(n4623), .Q(n4619) );
  nnd2s1 U5552 ( .DIN1(n4624), .DIN2(\NPC[17] ), .Q(n4623) );
  or2s1 U5553 ( .DIN1(n4625), .DIN2(n4626), .Q(n4624) );
  nnd2s1 U5554 ( .DIN1(n4625), .DIN2(n4626), .Q(n4622) );
  nnd2s1 U5555 ( .DIN1(n4583), .DIN2(n4627), .Q(n4618) );
  nnd2s1 U5556 ( .DIN1(n1372), .DIN2(n4585), .Q(n4627) );
  or2s1 U5557 ( .DIN1(n4412), .DIN2(n4422), .Q(n4420) );
  xor2s1 U5558 ( .DIN1(n4625), .DIN2(n4628), .Q(n4422) );
  xnr2s1 U5559 ( .DIN1(n9437), .DIN2(n4626), .Q(n4628) );
  nnd2s1 U5560 ( .DIN1(n4629), .DIN2(n4630), .Q(n4626) );
  nnd2s1 U5561 ( .DIN1(n4631), .DIN2(\NPC[16] ), .Q(n4630) );
  or2s1 U5562 ( .DIN1(n4632), .DIN2(n4633), .Q(n4631) );
  nnd2s1 U5563 ( .DIN1(n4632), .DIN2(n4633), .Q(n4629) );
  nnd2s1 U5564 ( .DIN1(n4583), .DIN2(n4634), .Q(n4625) );
  nnd2s1 U5565 ( .DIN1(n1312), .DIN2(n4585), .Q(n4634) );
  or2s1 U5566 ( .DIN1(n4404), .DIN2(n4414), .Q(n4412) );
  xor2s1 U5567 ( .DIN1(n4632), .DIN2(n4635), .Q(n4414) );
  xnr2s1 U5568 ( .DIN1(n9438), .DIN2(n4633), .Q(n4635) );
  nnd2s1 U5569 ( .DIN1(n4636), .DIN2(n4637), .Q(n4633) );
  nnd2s1 U5570 ( .DIN1(n4638), .DIN2(\NPC[15] ), .Q(n4637) );
  or2s1 U5571 ( .DIN1(n92), .DIN2(n4639), .Q(n4638) );
  nnd2s1 U5572 ( .DIN1(n4639), .DIN2(n92), .Q(n4636) );
  nnd2s1 U5573 ( .DIN1(n4583), .DIN2(n4640), .Q(n4632) );
  nnd2s1 U5574 ( .DIN1(n1198), .DIN2(n4585), .Q(n4640) );
  or2s1 U5575 ( .DIN1(n4396), .DIN2(n4406), .Q(n4404) );
  xnr2s1 U5576 ( .DIN1(n4641), .DIN2(n4639), .Q(n4406) );
  nnd2s1 U5577 ( .DIN1(n4642), .DIN2(n4643), .Q(n4639) );
  nnd2s1 U5578 ( .DIN1(n4644), .DIN2(\NPC[14] ), .Q(n4643) );
  or2s1 U5579 ( .DIN1(n97), .DIN2(n4645), .Q(n4644) );
  nnd2s1 U5580 ( .DIN1(n4645), .DIN2(n97), .Q(n4642) );
  xnr2s1 U5581 ( .DIN1(n9439), .DIN2(n9387), .Q(n4641) );
  or2s1 U5582 ( .DIN1(n4388), .DIN2(n4398), .Q(n4396) );
  xor2s1 U5583 ( .DIN1(n4645), .DIN2(n4646), .Q(n4398) );
  xnr2s1 U5584 ( .DIN1(n97), .DIN2(n9440), .Q(n4646) );
  nnd2s1 U5585 ( .DIN1(n4647), .DIN2(n4648), .Q(n4645) );
  nnd2s1 U5586 ( .DIN1(n4649), .DIN2(\NPC[13] ), .Q(n4648) );
  or2s1 U5587 ( .DIN1(n113), .DIN2(n4650), .Q(n4649) );
  nnd2s1 U5588 ( .DIN1(n4650), .DIN2(n113), .Q(n4647) );
  or2s1 U5589 ( .DIN1(n4380), .DIN2(n4390), .Q(n4388) );
  xnr2s1 U5590 ( .DIN1(n4651), .DIN2(n4650), .Q(n4390) );
  nnd2s1 U5591 ( .DIN1(n4652), .DIN2(n4653), .Q(n4650) );
  nnd2s1 U5592 ( .DIN1(n4654), .DIN2(\NPC[12] ), .Q(n4653) );
  or2s1 U5593 ( .DIN1(n98), .DIN2(n4655), .Q(n4654) );
  nnd2s1 U5594 ( .DIN1(n4655), .DIN2(n98), .Q(n4652) );
  xnr2s1 U5595 ( .DIN1(n9441), .DIN2(n9386), .Q(n4651) );
  or2s1 U5596 ( .DIN1(n4372), .DIN2(n4382), .Q(n4380) );
  xor2s1 U5597 ( .DIN1(n4655), .DIN2(n4656), .Q(n4382) );
  xnr2s1 U5598 ( .DIN1(n98), .DIN2(n9442), .Q(n4656) );
  nnd2s1 U5599 ( .DIN1(n4657), .DIN2(n4658), .Q(n4655) );
  nnd2s1 U5600 ( .DIN1(n4659), .DIN2(\NPC[11] ), .Q(n4658) );
  or2s1 U5601 ( .DIN1(n114), .DIN2(n4660), .Q(n4659) );
  nnd2s1 U5602 ( .DIN1(n4660), .DIN2(n114), .Q(n4657) );
  or2s1 U5603 ( .DIN1(n4364), .DIN2(n4374), .Q(n4372) );
  xnr2s1 U5604 ( .DIN1(n4661), .DIN2(n4660), .Q(n4374) );
  nnd2s1 U5605 ( .DIN1(n4662), .DIN2(n4663), .Q(n4660) );
  nnd2s1 U5606 ( .DIN1(n4664), .DIN2(\NPC[10] ), .Q(n4663) );
  or2s1 U5607 ( .DIN1(n110), .DIN2(n4665), .Q(n4664) );
  nnd2s1 U5608 ( .DIN1(n4665), .DIN2(n110), .Q(n4662) );
  xnr2s1 U5609 ( .DIN1(n9443), .DIN2(n9385), .Q(n4661) );
  or2s1 U5610 ( .DIN1(n4356), .DIN2(n4366), .Q(n4364) );
  xor2s1 U5611 ( .DIN1(n4665), .DIN2(n4666), .Q(n4366) );
  xnr2s1 U5612 ( .DIN1(n110), .DIN2(n9444), .Q(n4666) );
  nnd2s1 U5613 ( .DIN1(n4667), .DIN2(n4668), .Q(n4665) );
  nnd2s1 U5614 ( .DIN1(n4669), .DIN2(\NPC[9] ), .Q(n4668) );
  or2s1 U5615 ( .DIN1(n125), .DIN2(n4670), .Q(n4669) );
  nnd2s1 U5616 ( .DIN1(n4670), .DIN2(n125), .Q(n4667) );
  or2s1 U5617 ( .DIN1(n4348), .DIN2(n4358), .Q(n4356) );
  xnr2s1 U5618 ( .DIN1(n4671), .DIN2(n4670), .Q(n4358) );
  nnd2s1 U5619 ( .DIN1(n4672), .DIN2(n4673), .Q(n4670) );
  nnd2s1 U5620 ( .DIN1(n4674), .DIN2(\NPC[8] ), .Q(n4673) );
  or2s1 U5621 ( .DIN1(n111), .DIN2(n4675), .Q(n4674) );
  nnd2s1 U5622 ( .DIN1(n4675), .DIN2(n111), .Q(n4672) );
  xnr2s1 U5623 ( .DIN1(n9445), .DIN2(n9392), .Q(n4671) );
  or2s1 U5624 ( .DIN1(n4341), .DIN2(n4350), .Q(n4348) );
  xor2s1 U5625 ( .DIN1(n4675), .DIN2(n4676), .Q(n4350) );
  xnr2s1 U5626 ( .DIN1(n111), .DIN2(n9446), .Q(n4676) );
  nnd2s1 U5627 ( .DIN1(n4677), .DIN2(n4678), .Q(n4675) );
  nnd2s1 U5628 ( .DIN1(n4679), .DIN2(\NPC[7] ), .Q(n4678) );
  or2s1 U5629 ( .DIN1(n126), .DIN2(n4680), .Q(n4679) );
  nnd2s1 U5630 ( .DIN1(n4680), .DIN2(n126), .Q(n4677) );
  nnd2s1 U5631 ( .DIN1(n4331), .DIN2(n4342), .Q(n4341) );
  xor2s1 U5632 ( .DIN1(n4681), .DIN2(n4680), .Q(n4342) );
  nnd2s1 U5633 ( .DIN1(n4682), .DIN2(n4683), .Q(n4680) );
  nnd2s1 U5634 ( .DIN1(n4684), .DIN2(\NPC[6] ), .Q(n4683) );
  or2s1 U5635 ( .DIN1(n112), .DIN2(n4685), .Q(n4684) );
  nnd2s1 U5636 ( .DIN1(n4685), .DIN2(n112), .Q(n4682) );
  xnr2s1 U5637 ( .DIN1(n9447), .DIN2(n9391), .Q(n4681) );
  nor2s1 U5638 ( .DIN1(n4320), .DIN2(n4330), .Q(n4331) );
  xor2s1 U5639 ( .DIN1(n4685), .DIN2(n4686), .Q(n4330) );
  xnr2s1 U5640 ( .DIN1(n112), .DIN2(n9448), .Q(n4686) );
  nnd2s1 U5641 ( .DIN1(n4687), .DIN2(n4688), .Q(n4685) );
  nnd2s1 U5642 ( .DIN1(n4689), .DIN2(\NPC[5] ), .Q(n4688) );
  or2s1 U5643 ( .DIN1(n115), .DIN2(n4690), .Q(n4689) );
  nnd2s1 U5644 ( .DIN1(n4690), .DIN2(n115), .Q(n4687) );
  or2s1 U5645 ( .DIN1(n4312), .DIN2(n4322), .Q(n4320) );
  xnr2s1 U5646 ( .DIN1(n4691), .DIN2(n4690), .Q(n4322) );
  nnd2s1 U5647 ( .DIN1(n4692), .DIN2(n4693), .Q(n4690) );
  nnd2s1 U5648 ( .DIN1(n4694), .DIN2(\NPC[4] ), .Q(n4693) );
  or2s1 U5649 ( .DIN1(n99), .DIN2(n4695), .Q(n4694) );
  nnd2s1 U5650 ( .DIN1(n4695), .DIN2(n99), .Q(n4692) );
  xnr2s1 U5651 ( .DIN1(n9449), .DIN2(n9390), .Q(n4691) );
  or2s1 U5652 ( .DIN1(n4304), .DIN2(n4314), .Q(n4312) );
  xor2s1 U5653 ( .DIN1(n4695), .DIN2(n4696), .Q(n4314) );
  xnr2s1 U5654 ( .DIN1(n99), .DIN2(n9450), .Q(n4696) );
  nnd2s1 U5655 ( .DIN1(n4697), .DIN2(n4698), .Q(n4695) );
  nnd2s1 U5656 ( .DIN1(n4699), .DIN2(\NPC[3] ), .Q(n4698) );
  or2s1 U5657 ( .DIN1(n116), .DIN2(n4700), .Q(n4699) );
  nnd2s1 U5658 ( .DIN1(n4700), .DIN2(n116), .Q(n4697) );
  or2s1 U5659 ( .DIN1(n4306), .DIN2(n4297), .Q(n4304) );
  xor2s1 U5660 ( .DIN1(n4701), .DIN2(n4702), .Q(n4297) );
  xnr2s1 U5661 ( .DIN1(n100), .DIN2(n9491), .Q(n4702) );
  xnr2s1 U5662 ( .DIN1(n4703), .DIN2(n4700), .Q(n4306) );
  nnd2s1 U5663 ( .DIN1(n4704), .DIN2(n4705), .Q(n4700) );
  nnd2s1 U5664 ( .DIN1(n4706), .DIN2(\NPC[2] ), .Q(n4705) );
  or2s1 U5665 ( .DIN1(n100), .DIN2(n4701), .Q(n4706) );
  nnd2s1 U5666 ( .DIN1(n4701), .DIN2(n100), .Q(n4704) );
  nnd2s1 U5667 ( .DIN1(n4707), .DIN2(n4708), .Q(n4701) );
  nnd3s1 U5668 ( .DIN1(\IFinst/N7 ), .DIN2(n41), .DIN3(n4709), .Q(n4708) );
  nnd2s1 U5669 ( .DIN1(n9388), .DIN2(n9422), .Q(n4709) );
  nnd2s1 U5670 ( .DIN1(\IFinst/N8 ), .DIN2(n42), .Q(n4707) );
  xnr2s1 U5671 ( .DIN1(n9451), .DIN2(n9389), .Q(n4703) );
  xnr2s1 U5672 ( .DIN1(n9424), .DIN2(n4543), .Q(n4537) );
  nnd2s1 U5673 ( .DIN1(n4583), .DIN2(n4710), .Q(n4543) );
  nnd2s1 U5674 ( .DIN1(\IDinst/N43 ), .DIN2(n4585), .Q(n4710) );
  nnd2s1 U5675 ( .DIN1(n4168), .DIN2(n92), .Q(n4583) );
  hi1s1 U5676 ( .DIN(n4298), .Q(n4283) );
  nnd2s1 U5677 ( .DIN1(n4149), .DIN2(n4711), .Q(n4298) );
  or4s1 U5678 ( .DIN1(n4534), .DIN2(n4711), .DIN3(n1921), .DIN4(n4713), 
        .Q(n4712) );
  nnd3s1 U5679 ( .DIN1(n4535), .DIN2(n4157), .DIN3(n4714), .Q(n4713) );
  nnd3s1 U5680 ( .DIN1(n4715), .DIN2(n4716), .DIN3(n4163), .Q(n4157) );
  nnd4s1 U5681 ( .DIN1(n4717), .DIN2(n4718), .DIN3(n1924), .DIN4(n1923), 
        .Q(n1921) );
  nnd3s1 U5682 ( .DIN1(n4719), .DIN2(n4720), .DIN3(n4160), .Q(n1923) );
  nnd3s1 U5683 ( .DIN1(n4160), .DIN2(n4721), .DIN3(n4722), .Q(n1924) );
  nnd2s1 U5684 ( .DIN1(n4723), .DIN2(n4724), .Q(n4718) );
  nnd2s1 U5685 ( .DIN1(n4725), .DIN2(n4726), .Q(n4717) );
  or2s1 U5686 ( .DIN1(n4585), .DIN2(n4168), .Q(n4711) );
  nor2s1 U5687 ( .DIN1(n4727), .DIN2(n4728), .Q(n4168) );
  nnd2s1 U5688 ( .DIN1(n4729), .DIN2(n4166), .Q(n4585) );
  nnd4s1 U5689 ( .DIN1(n4730), .DIN2(n4731), .DIN3(n4732), .DIN4(n1953), 
        .Q(n4166) );
  nnd2s1 U5690 ( .DIN1(n4733), .DIN2(n4167), .Q(n4534) );
  nnd2s1 U5691 ( .DIN1(n4734), .DIN2(n4716), .Q(n4167) );
  nnd2s1 U5692 ( .DIN1(n4735), .DIN2(n4736), .Q(\IDinst/n4792 ) );
  nnd2s1 U5693 ( .DIN1(n652), .DIN2(n124), .Q(n4736) );
  nnd2s1 U5694 ( .DIN1(n4737), .DIN2(n4738), .Q(\IDinst/n4791 ) );
  nnd2s1 U5695 ( .DIN1(n637), .DIN2(n124), .Q(n4738) );
  nnd2s1 U5696 ( .DIN1(n677), .DIN2(n282), .Q(n4737) );
  nnd2s1 U5697 ( .DIN1(n4735), .DIN2(n4739), .Q(\IDinst/n4790 ) );
  nnd2s1 U5698 ( .DIN1(n651), .DIN2(n96), .Q(n4739) );
  nnd2s1 U5699 ( .DIN1(n4740), .DIN2(n4741), .Q(\IDinst/n4789 ) );
  nnd2s1 U5700 ( .DIN1(n640), .DIN2(n96), .Q(n4741) );
  nnd2s1 U5701 ( .DIN1(n678), .DIN2(n283), .Q(n4740) );
  nnd2s1 U5702 ( .DIN1(n4735), .DIN2(n4742), .Q(\IDinst/n4788 ) );
  nnd2s1 U5703 ( .DIN1(n650), .DIN2(n14), .Q(n4742) );
  nnd2s1 U5704 ( .DIN1(n4743), .DIN2(n4744), .Q(\IDinst/n4787 ) );
  nnd2s1 U5705 ( .DIN1(n639), .DIN2(n14), .Q(n4744) );
  nnd2s1 U5706 ( .DIN1(n675), .DIN2(n284), .Q(n4743) );
  nnd2s1 U5707 ( .DIN1(n4735), .DIN2(n4745), .Q(\IDinst/n4786 ) );
  nnd2s1 U5708 ( .DIN1(n649), .DIN2(n102), .Q(n4745) );
  nnd2s1 U5709 ( .DIN1(n4746), .DIN2(n4747), .Q(\IDinst/n4785 ) );
  nnd2s1 U5710 ( .DIN1(n638), .DIN2(n102), .Q(n4747) );
  nnd2s1 U5711 ( .DIN1(n676), .DIN2(n285), .Q(n4746) );
  nnd2s1 U5712 ( .DIN1(n4735), .DIN2(n4748), .Q(\IDinst/n4784 ) );
  nnd2s1 U5713 ( .DIN1(n652), .DIN2(n95), .Q(n4748) );
  nnd2s1 U5714 ( .DIN1(n4749), .DIN2(n4750), .Q(\IDinst/n4783 ) );
  nnd2s1 U5715 ( .DIN1(n637), .DIN2(n95), .Q(n4750) );
  nnd2s1 U5716 ( .DIN1(n677), .DIN2(n286), .Q(n4749) );
  nnd2s1 U5717 ( .DIN1(n4735), .DIN2(n4751), .Q(\IDinst/n4782 ) );
  nnd2s1 U5718 ( .DIN1(n651), .DIN2(n103), .Q(n4751) );
  nnd2s1 U5719 ( .DIN1(n4752), .DIN2(n4753), .Q(\IDinst/n4781 ) );
  nnd2s1 U5720 ( .DIN1(n640), .DIN2(n103), .Q(n4753) );
  nnd2s1 U5721 ( .DIN1(n678), .DIN2(n287), .Q(n4752) );
  nnd2s1 U5722 ( .DIN1(n4735), .DIN2(n4754), .Q(\IDinst/n4780 ) );
  nnd2s1 U5723 ( .DIN1(n650), .DIN2(n15), .Q(n4754) );
  nnd2s1 U5724 ( .DIN1(n4755), .DIN2(n4756), .Q(\IDinst/n4779 ) );
  nnd2s1 U5725 ( .DIN1(n639), .DIN2(n15), .Q(n4756) );
  nnd2s1 U5726 ( .DIN1(n675), .DIN2(n288), .Q(n4755) );
  nnd2s1 U5727 ( .DIN1(n4735), .DIN2(n4757), .Q(\IDinst/n4778 ) );
  nnd2s1 U5728 ( .DIN1(n649), .DIN2(n120), .Q(n4757) );
  nnd2s1 U5729 ( .DIN1(n4758), .DIN2(n4759), .Q(\IDinst/n4777 ) );
  nnd2s1 U5730 ( .DIN1(n638), .DIN2(n120), .Q(n4759) );
  nnd2s1 U5731 ( .DIN1(n676), .DIN2(n289), .Q(n4758) );
  nnd2s1 U5732 ( .DIN1(n4735), .DIN2(n4760), .Q(\IDinst/n4776 ) );
  nnd2s1 U5733 ( .DIN1(n652), .DIN2(n93), .Q(n4760) );
  nnd2s1 U5734 ( .DIN1(n4761), .DIN2(n4762), .Q(\IDinst/n4775 ) );
  nnd2s1 U5735 ( .DIN1(n637), .DIN2(n93), .Q(n4762) );
  nnd2s1 U5736 ( .DIN1(n677), .DIN2(n290), .Q(n4761) );
  nnd2s1 U5737 ( .DIN1(n4735), .DIN2(n4763), .Q(\IDinst/n4774 ) );
  nnd2s1 U5738 ( .DIN1(n651), .DIN2(n121), .Q(n4763) );
  nnd2s1 U5739 ( .DIN1(n4764), .DIN2(n4765), .Q(\IDinst/n4773 ) );
  nnd2s1 U5740 ( .DIN1(n640), .DIN2(n121), .Q(n4765) );
  nnd2s1 U5741 ( .DIN1(n678), .DIN2(n291), .Q(n4764) );
  nnd2s1 U5742 ( .DIN1(n4735), .DIN2(n4766), .Q(\IDinst/n4772 ) );
  nnd2s1 U5743 ( .DIN1(n650), .DIN2(n16), .Q(n4766) );
  nnd2s1 U5744 ( .DIN1(n4767), .DIN2(n4768), .Q(\IDinst/n4771 ) );
  nnd2s1 U5745 ( .DIN1(n639), .DIN2(n16), .Q(n4768) );
  nnd2s1 U5746 ( .DIN1(n675), .DIN2(n292), .Q(n4767) );
  nnd2s1 U5747 ( .DIN1(n4735), .DIN2(n4769), .Q(\IDinst/n4770 ) );
  nnd2s1 U5748 ( .DIN1(n649), .DIN2(n123), .Q(n4769) );
  nnd2s1 U5749 ( .DIN1(n4770), .DIN2(n4771), .Q(\IDinst/n4769 ) );
  nnd2s1 U5750 ( .DIN1(n638), .DIN2(n123), .Q(n4771) );
  nnd2s1 U5751 ( .DIN1(n676), .DIN2(n293), .Q(n4770) );
  nnd2s1 U5752 ( .DIN1(n4735), .DIN2(n4772), .Q(\IDinst/n4768 ) );
  nnd2s1 U5753 ( .DIN1(n652), .DIN2(n94), .Q(n4772) );
  nnd2s1 U5754 ( .DIN1(n4773), .DIN2(n4774), .Q(\IDinst/n4767 ) );
  nnd2s1 U5755 ( .DIN1(n637), .DIN2(n94), .Q(n4774) );
  nnd2s1 U5756 ( .DIN1(n677), .DIN2(n294), .Q(n4773) );
  nnd2s1 U5757 ( .DIN1(n4735), .DIN2(n4775), .Q(\IDinst/n4766 ) );
  nnd2s1 U5758 ( .DIN1(n651), .DIN2(n122), .Q(n4775) );
  nnd2s1 U5759 ( .DIN1(n4776), .DIN2(n4777), .Q(\IDinst/n4765 ) );
  nnd2s1 U5760 ( .DIN1(n640), .DIN2(n122), .Q(n4777) );
  nnd2s1 U5761 ( .DIN1(n678), .DIN2(n295), .Q(n4776) );
  nnd2s1 U5762 ( .DIN1(n4735), .DIN2(n4778), .Q(\IDinst/n4764 ) );
  nnd2s1 U5763 ( .DIN1(n650), .DIN2(n13), .Q(n4778) );
  nnd2s1 U5764 ( .DIN1(n4779), .DIN2(n4780), .Q(\IDinst/n4763 ) );
  nnd2s1 U5765 ( .DIN1(n639), .DIN2(n13), .Q(n4780) );
  nnd2s1 U5766 ( .DIN1(n675), .DIN2(n296), .Q(n4779) );
  nnd2s1 U5767 ( .DIN1(n4735), .DIN2(n4781), .Q(\IDinst/n4762 ) );
  nnd2s1 U5768 ( .DIN1(n649), .DIN2(n109), .Q(n4781) );
  nnd3s1 U5769 ( .DIN1(n4782), .DIN2(n92), .DIN3(n436), .Q(n4735) );
  nnd4s1 U5770 ( .DIN1(n4783), .DIN2(n4730), .DIN3(n4784), .DIN4(n4133), 
        .Q(n4782) );
  nor2s1 U5771 ( .DIN1(n4785), .DIN2(n4786), .Q(n4784) );
  nnd2s1 U5772 ( .DIN1(n4787), .DIN2(n4788), .Q(\IDinst/n4761 ) );
  nnd2s1 U5773 ( .DIN1(n638), .DIN2(n109), .Q(n4788) );
  nnd2s1 U5774 ( .DIN1(n676), .DIN2(n297), .Q(n4787) );
  nnd2s1 U5775 ( .DIN1(n4789), .DIN2(n4790), .Q(\IDinst/n4760 ) );
  nnd2s1 U5776 ( .DIN1(n436), .DIN2(n92), .Q(n4790) );
  nnd2s1 U5777 ( .DIN1(n652), .DIN2(n7), .Q(n4789) );
  nnd2s1 U5778 ( .DIN1(n4791), .DIN2(n4792), .Q(\IDinst/n4759 ) );
  nnd2s1 U5779 ( .DIN1(n637), .DIN2(n7), .Q(n4792) );
  nnd2s1 U5780 ( .DIN1(n677), .DIN2(n298), .Q(n4791) );
  nnd2s1 U5781 ( .DIN1(n4793), .DIN2(n4794), .Q(\IDinst/n4758 ) );
  nnd2s1 U5782 ( .DIN1(n437), .DIN2(n97), .Q(n4794) );
  nnd2s1 U5783 ( .DIN1(n651), .DIN2(n108), .Q(n4793) );
  nnd2s1 U5784 ( .DIN1(n4795), .DIN2(n4796), .Q(\IDinst/n4757 ) );
  nnd2s1 U5785 ( .DIN1(n640), .DIN2(n108), .Q(n4796) );
  nnd2s1 U5786 ( .DIN1(n678), .DIN2(n299), .Q(n4795) );
  nnd2s1 U5787 ( .DIN1(n4797), .DIN2(n4798), .Q(\IDinst/n4756 ) );
  nnd2s1 U5788 ( .DIN1(n436), .DIN2(n113), .Q(n4798) );
  nnd2s1 U5789 ( .DIN1(n650), .DIN2(n9), .Q(n4797) );
  nnd2s1 U5790 ( .DIN1(n4799), .DIN2(n4800), .Q(\IDinst/n4755 ) );
  nnd2s1 U5791 ( .DIN1(n639), .DIN2(n9), .Q(n4800) );
  nnd2s1 U5792 ( .DIN1(n675), .DIN2(n300), .Q(n4799) );
  nnd2s1 U5793 ( .DIN1(n4801), .DIN2(n4802), .Q(\IDinst/n4754 ) );
  nnd2s1 U5794 ( .DIN1(n437), .DIN2(n98), .Q(n4802) );
  nnd2s1 U5795 ( .DIN1(n649), .DIN2(n106), .Q(n4801) );
  nnd2s1 U5796 ( .DIN1(n4803), .DIN2(n4804), .Q(\IDinst/n4753 ) );
  nnd2s1 U5797 ( .DIN1(n638), .DIN2(n106), .Q(n4804) );
  nnd2s1 U5798 ( .DIN1(n676), .DIN2(n301), .Q(n4803) );
  nnd2s1 U5799 ( .DIN1(n4805), .DIN2(n4806), .Q(\IDinst/n4752 ) );
  nnd2s1 U5800 ( .DIN1(n436), .DIN2(n114), .Q(n4806) );
  nnd2s1 U5801 ( .DIN1(n652), .DIN2(n8), .Q(n4805) );
  nnd2s1 U5802 ( .DIN1(n4807), .DIN2(n4808), .Q(\IDinst/n4751 ) );
  nnd2s1 U5803 ( .DIN1(n637), .DIN2(n8), .Q(n4808) );
  nnd2s1 U5804 ( .DIN1(n677), .DIN2(n302), .Q(n4807) );
  nnd2s1 U5805 ( .DIN1(n4809), .DIN2(n4810), .Q(\IDinst/n4750 ) );
  nnd2s1 U5806 ( .DIN1(n437), .DIN2(n110), .Q(n4810) );
  nnd2s1 U5807 ( .DIN1(n651), .DIN2(n104), .Q(n4809) );
  nnd2s1 U5808 ( .DIN1(n4811), .DIN2(n4812), .Q(\IDinst/n4749 ) );
  nnd2s1 U5809 ( .DIN1(n640), .DIN2(n104), .Q(n4812) );
  nnd2s1 U5810 ( .DIN1(n678), .DIN2(n303), .Q(n4811) );
  nnd2s1 U5811 ( .DIN1(n4813), .DIN2(n4814), .Q(\IDinst/n4748 ) );
  nnd2s1 U5812 ( .DIN1(n436), .DIN2(n125), .Q(n4814) );
  nnd2s1 U5813 ( .DIN1(n650), .DIN2(n75), .Q(n4813) );
  nnd2s1 U5814 ( .DIN1(n4815), .DIN2(n4816), .Q(\IDinst/n4747 ) );
  nnd2s1 U5815 ( .DIN1(n639), .DIN2(n75), .Q(n4816) );
  nnd2s1 U5816 ( .DIN1(n675), .DIN2(n304), .Q(n4815) );
  nnd2s1 U5817 ( .DIN1(n4817), .DIN2(n4818), .Q(\IDinst/n4746 ) );
  nnd2s1 U5818 ( .DIN1(n437), .DIN2(n111), .Q(n4818) );
  nnd2s1 U5819 ( .DIN1(n649), .DIN2(n107), .Q(n4817) );
  nnd2s1 U5820 ( .DIN1(n4819), .DIN2(n4820), .Q(\IDinst/n4745 ) );
  nnd2s1 U5821 ( .DIN1(n638), .DIN2(n107), .Q(n4820) );
  nnd2s1 U5822 ( .DIN1(n676), .DIN2(n305), .Q(n4819) );
  nnd2s1 U5823 ( .DIN1(n4821), .DIN2(n4822), .Q(\IDinst/n4744 ) );
  nnd2s1 U5824 ( .DIN1(n436), .DIN2(n126), .Q(n4822) );
  nnd2s1 U5825 ( .DIN1(n652), .DIN2(n76), .Q(n4821) );
  nnd2s1 U5826 ( .DIN1(n4823), .DIN2(n4824), .Q(\IDinst/n4743 ) );
  nnd2s1 U5827 ( .DIN1(n637), .DIN2(n76), .Q(n4824) );
  nnd2s1 U5828 ( .DIN1(n677), .DIN2(n264), .Q(n4823) );
  nnd2s1 U5829 ( .DIN1(n4825), .DIN2(n4826), .Q(\IDinst/n4742 ) );
  nnd2s1 U5830 ( .DIN1(n437), .DIN2(n112), .Q(n4826) );
  nnd2s1 U5831 ( .DIN1(n651), .DIN2(n105), .Q(n4825) );
  nnd2s1 U5832 ( .DIN1(n4827), .DIN2(n4828), .Q(\IDinst/n4741 ) );
  nnd2s1 U5833 ( .DIN1(n640), .DIN2(n105), .Q(n4828) );
  nnd2s1 U5834 ( .DIN1(n678), .DIN2(n265), .Q(n4827) );
  nnd2s1 U5835 ( .DIN1(n4829), .DIN2(n4830), .Q(\IDinst/n4740 ) );
  nnd2s1 U5836 ( .DIN1(n436), .DIN2(n115), .Q(n4830) );
  nnd2s1 U5837 ( .DIN1(n650), .DIN2(n4831), .Q(n4829) );
  nnd2s1 U5838 ( .DIN1(n4832), .DIN2(n4833), .Q(\IDinst/n4739 ) );
  nnd2s1 U5839 ( .DIN1(n639), .DIN2(n4831), .Q(n4833) );
  nnd2s1 U5840 ( .DIN1(n675), .DIN2(n266), .Q(n4832) );
  nnd2s1 U5841 ( .DIN1(n4834), .DIN2(n4835), .Q(\IDinst/n4738 ) );
  nnd2s1 U5842 ( .DIN1(n437), .DIN2(n99), .Q(n4835) );
  nnd2s1 U5843 ( .DIN1(n649), .DIN2(n805), .Q(n4834) );
  nnd2s1 U5844 ( .DIN1(n4836), .DIN2(n4837), .Q(\IDinst/n4737 ) );
  nnd2s1 U5845 ( .DIN1(n638), .DIN2(n806), .Q(n4837) );
  nnd2s1 U5846 ( .DIN1(n676), .DIN2(n267), .Q(n4836) );
  nnd2s1 U5847 ( .DIN1(n4838), .DIN2(n4839), .Q(\IDinst/n4736 ) );
  nnd2s1 U5848 ( .DIN1(n436), .DIN2(n116), .Q(n4839) );
  nnd2s1 U5849 ( .DIN1(n652), .DIN2(n4840), .Q(n4838) );
  nnd2s1 U5850 ( .DIN1(n4841), .DIN2(n4842), .Q(\IDinst/n4735 ) );
  nnd2s1 U5851 ( .DIN1(n637), .DIN2(n803), .Q(n4842) );
  nnd2s1 U5852 ( .DIN1(n677), .DIN2(n268), .Q(n4841) );
  nnd2s1 U5853 ( .DIN1(n4843), .DIN2(n4844), .Q(\IDinst/n4734 ) );
  nnd2s1 U5854 ( .DIN1(n437), .DIN2(n100), .Q(n4844) );
  nnd2s1 U5855 ( .DIN1(n651), .DIN2(n792), .Q(n4843) );
  nnd2s1 U5856 ( .DIN1(n4846), .DIN2(n4847), .Q(\IDinst/n4733 ) );
  nnd2s1 U5857 ( .DIN1(n640), .DIN2(n792), .Q(n4847) );
  nnd2s1 U5858 ( .DIN1(n678), .DIN2(n269), .Q(n4846) );
  nnd2s1 U5859 ( .DIN1(n4848), .DIN2(n4849), .Q(\IDinst/n4732 ) );
  nnd2s1 U5860 ( .DIN1(n436), .DIN2(n42), .Q(n4849) );
  nnd2s1 U5861 ( .DIN1(n650), .DIN2(n707), .Q(n4848) );
  nnd2s1 U5862 ( .DIN1(n4850), .DIN2(n4851), .Q(\IDinst/n4731 ) );
  nnd2s1 U5863 ( .DIN1(n639), .DIN2(n707), .Q(n4851) );
  nnd2s1 U5864 ( .DIN1(n675), .DIN2(n270), .Q(n4850) );
  nnd2s1 U5865 ( .DIN1(n4852), .DIN2(n4853), .Q(\IDinst/n4730 ) );
  nnd2s1 U5866 ( .DIN1(n437), .DIN2(n41), .Q(n4853) );
  or2s1 U5867 ( .DIN1(n4144), .DIN2(n4854), .Q(n4128) );
  nnd4s1 U5868 ( .DIN1(n4855), .DIN2(n4856), .DIN3(n4857), .DIN4(n4714), 
        .Q(n4144) );
  nnd3s1 U5869 ( .DIN1(n4124), .DIN2(n4727), .DIN3(n4734), .Q(n4714) );
  hi1s1 U5870 ( .DIN(n4728), .Q(n4734) );
  nnd2s1 U5871 ( .DIN1(n4858), .DIN2(n4859), .Q(n4728) );
  hi1s1 U5872 ( .DIN(n4860), .Q(n4858) );
  nnd4s1 U5873 ( .DIN1(n4715), .DIN2(n4116), .DIN3(n4783), .DIN4(n1956), 
        .Q(n4727) );
  nor2s1 U5874 ( .DIN1(n1962), .DIN2(n1959), .Q(n4116) );
  nnd3s1 U5875 ( .DIN1(n4861), .DIN2(n4862), .DIN3(n4160), .Q(n4857) );
  nnd2s1 U5876 ( .DIN1(n4722), .DIN2(n4721), .Q(n4862) );
  nnd2s1 U5877 ( .DIN1(n4863), .DIN2(n4864), .Q(n4721) );
  nnd3s1 U5878 ( .DIN1(n4865), .DIN2(n40), .DIN3(n4866), .Q(n4864) );
  nnd2s1 U5879 ( .DIN1(n4867), .DIN2(n4868), .Q(n4861) );
  or2s1 U5880 ( .DIN1(n4720), .DIN2(n4869), .Q(n4867) );
  nnd2s1 U5881 ( .DIN1(n4863), .DIN2(n4870), .Q(n4720) );
  nnd3s1 U5882 ( .DIN1(n4871), .DIN2(n40), .DIN3(n4866), .Q(n4870) );
  and2s1 U5883 ( .DIN1(n4872), .DIN2(n4873), .Q(n4863) );
  nnd4s1 U5884 ( .DIN1(n4874), .DIN2(n4875), .DIN3(n4876), .DIN4(n4877), 
        .Q(n4873) );
  hi1s1 U5885 ( .DIN(n4878), .Q(n4877) );
  nor2s1 U5886 ( .DIN1(IR_opcode_field[4]), .DIN2(IR_opcode_field[3]), 
        .Q(n4876) );
  nnd2s1 U5887 ( .DIN1(n4879), .DIN2(n117), .Q(n4875) );
  nnd2s1 U5888 ( .DIN1(n39), .DIN2(n132), .Q(n4879) );
  nnd2s1 U5889 ( .DIN1(IR_opcode_field[2]), .DIN2(IR_opcode_field[1]), 
        .Q(n4874) );
  nnd3s1 U5890 ( .DIN1(n4880), .DIN2(n4881), .DIN3(n117), .Q(n4872) );
  nnd2s1 U5891 ( .DIN1(n4882), .DIN2(n4883), .Q(n4881) );
  nnd2s1 U5892 ( .DIN1(n4884), .DIN2(n4885), .Q(n4883) );
  nnd2s1 U5893 ( .DIN1(IR_opcode_field[3]), .DIN2(IR_opcode_field[1]), 
        .Q(n4885) );
  or2s1 U5894 ( .DIN1(n4882), .DIN2(IR_opcode_field[3]), .Q(n4880) );
  nor2s1 U5895 ( .DIN1(n101), .DIN2(n39), .Q(n4882) );
  nnd2s1 U5896 ( .DIN1(n4886), .DIN2(n4723), .Q(n4856) );
  and3s1 U5897 ( .DIN1(n4887), .DIN2(n4160), .DIN3(n4888), .Q(n4723) );
  hi1s1 U5898 ( .DIN(n4889), .Q(n4888) );
  hi1s1 U5899 ( .DIN(n4724), .Q(n4886) );
  nnd2s1 U5900 ( .DIN1(n4890), .DIN2(n4891), .Q(n4724) );
  nnd2s1 U5901 ( .DIN1(n4892), .DIN2(n4865), .Q(n4891) );
  nnd2s1 U5902 ( .DIN1(n4893), .DIN2(n4894), .Q(n4865) );
  nnd4s1 U5903 ( .DIN1(n4133), .DIN2(n4730), .DIN3(n4895), .DIN4(n4896), 
        .Q(n4894) );
  nnd2s1 U5904 ( .DIN1(n1950), .DIN2(n4783), .Q(n4895) );
  nnd2s1 U5905 ( .DIN1(n4783), .DIN2(n4897), .Q(n4893) );
  nnd3s1 U5906 ( .DIN1(n4898), .DIN2(n4899), .DIN3(n4900), .Q(n4897) );
  or3s1 U5907 ( .DIN1(n4133), .DIN2(n4901), .DIN3(n1953), .Q(n4900) );
  nnd3s1 U5908 ( .DIN1(n1953), .DIN2(n1962), .DIN3(n4785), .Q(n4899) );
  nnd2s1 U5909 ( .DIN1(n1959), .DIN2(n4902), .Q(n4898) );
  nnd3s1 U5910 ( .DIN1(n1956), .DIN2(n4903), .DIN3(n1953), .Q(n4902) );
  nnd2s1 U5911 ( .DIN1(n4730), .DIN2(n4786), .Q(n4903) );
  nnd2s1 U5912 ( .DIN1(n4904), .DIN2(n4725), .Q(n4855) );
  nor2s1 U5913 ( .DIN1(n4859), .DIN2(n4860), .Q(n4725) );
  nnd3s1 U5914 ( .DIN1(n4160), .DIN2(n4889), .DIN3(n4887), .Q(n4860) );
  nor2s1 U5915 ( .DIN1(n4719), .DIN2(n4722), .Q(n4887) );
  hi1s1 U5916 ( .DIN(n4868), .Q(n4722) );
  nnd4s1 U5917 ( .DIN1(n4905), .DIN2(n4906), .DIN3(n4907), .DIN4(n4908), 
        .Q(n4868) );
  and3s1 U5918 ( .DIN1(n4909), .DIN2(n4910), .DIN3(n4911), .Q(n4908) );
  xnr2s1 U5919 ( .DIN1(\IDinst/reg_dst_of_EX[3]), .DIN2(n641), .Q(n4911) );
  xnr2s1 U5920 ( .DIN1(\IDinst/reg_dst_of_EX[4]), .DIN2(\IDinst/N43 ), 
        .Q(n4910) );
  xnr2s1 U5921 ( .DIN1(\IDinst/reg_dst_of_EX[2]), .DIN2(\IDinst/N41 ), 
        .Q(n4909) );
  xnr2s1 U5922 ( .DIN1(\IDinst/reg_dst_of_EX[0]), .DIN2(n1065), .Q(n4907) );
  xnr2s1 U5923 ( .DIN1(\IDinst/reg_dst_of_EX[1]), .DIN2(n1153), .Q(n4905) );
  hi1s1 U5924 ( .DIN(n4869), .Q(n4719) );
  nnd4s1 U5925 ( .DIN1(n4912), .DIN2(n4913), .DIN3(n4914), .DIN4(n4915), 
        .Q(n4869) );
  and3s1 U5926 ( .DIN1(n4916), .DIN2(n4917), .DIN3(n4918), .Q(n4915) );
  xnr2s1 U5927 ( .DIN1(\IDinst/reg_dst_of_EX[3]), .DIN2(n666), .Q(n4918) );
  nnd2s1 U5928 ( .DIN1(n4919), .DIN2(n4920), .Q(\IDinst/reg_dst_of_EX[3]) );
  nnd2s1 U5929 ( .DIN1(n49), .DIN2(n11), .Q(n4920) );
  nnd2s1 U5930 ( .DIN1(reg_dst), .DIN2(n50), .Q(n4919) );
  xnr2s1 U5931 ( .DIN1(\IDinst/reg_dst_of_EX[4]), .DIN2(n534), .Q(n4917) );
  nnd2s1 U5932 ( .DIN1(n4921), .DIN2(n4922), .Q(\IDinst/reg_dst_of_EX[4]) );
  nnd2s1 U5933 ( .DIN1(n141), .DIN2(n11), .Q(n4922) );
  nnd2s1 U5934 ( .DIN1(reg_dst), .DIN2(n142), .Q(n4921) );
  xnr2s1 U5935 ( .DIN1(\IDinst/reg_dst_of_EX[2]), .DIN2(n1372), .Q(n4916) );
  nnd2s1 U5936 ( .DIN1(n4923), .DIN2(n4924), .Q(\IDinst/reg_dst_of_EX[2]) );
  nnd2s1 U5937 ( .DIN1(n227), .DIN2(n11), .Q(n4924) );
  nnd2s1 U5938 ( .DIN1(reg_dst), .DIN2(n230), .Q(n4923) );
  xnr2s1 U5939 ( .DIN1(\IDinst/reg_dst_of_EX[0]), .DIN2(n1198), .Q(n4914) );
  nnd2s1 U5940 ( .DIN1(n4925), .DIN2(n4926), .Q(\IDinst/reg_dst_of_EX[0]) );
  nnd2s1 U5941 ( .DIN1(n229), .DIN2(n11), .Q(n4926) );
  nnd2s1 U5942 ( .DIN1(reg_dst), .DIN2(n232), .Q(n4925) );
  xnr2s1 U5943 ( .DIN1(\IDinst/reg_dst_of_EX[1]), .DIN2(n1312), .Q(n4912) );
  nnd2s1 U5944 ( .DIN1(n4927), .DIN2(n4928), .Q(\IDinst/reg_dst_of_EX[1]) );
  nnd2s1 U5945 ( .DIN1(n228), .DIN2(n11), .Q(n4928) );
  nnd2s1 U5946 ( .DIN1(reg_dst), .DIN2(n231), .Q(n4927) );
  nnd4s1 U5947 ( .DIN1(n4929), .DIN2(n4906), .DIN3(n4930), .DIN4(n4931), 
        .Q(n4889) );
  and3s1 U5948 ( .DIN1(n4932), .DIN2(n728), .DIN3(n4934), .Q(n4931) );
  xnr2s1 U5949 ( .DIN1(n9420), .DIN2(n671), .Q(n4934) );
  xnr2s1 U5950 ( .DIN1(n9421), .DIN2(n1181), .Q(n4932) );
  xnr2s1 U5951 ( .DIN1(n9452), .DIN2(n1025), .Q(n4930) );
  xnr2s1 U5952 ( .DIN1(n9455), .DIN2(n1133), .Q(n4929) );
  and2s1 U5953 ( .DIN1(n4731), .DIN2(n4935), .Q(n4160) );
  nnd3s1 U5954 ( .DIN1(n4732), .DIN2(n1953), .DIN3(n4730), .Q(n4935) );
  hi1s1 U5955 ( .DIN(n4936), .Q(n4731) );
  nnd4s1 U5956 ( .DIN1(n4937), .DIN2(n4913), .DIN3(n4938), .DIN4(n4939), 
        .Q(n4859) );
  and3s1 U5957 ( .DIN1(n4940), .DIN2(n762), .DIN3(n4942), .Q(n4939) );
  xnr2s1 U5958 ( .DIN1(n9420), .DIN2(n681), .Q(n4942) );
  xnr2s1 U5959 ( .DIN1(n9421), .DIN2(n1364), .Q(n4940) );
  xnr2s1 U5960 ( .DIN1(n9452), .DIN2(n1238), .Q(n4938) );
  xnr2s1 U5961 ( .DIN1(n9455), .DIN2(n1332), .Q(n4937) );
  hi1s1 U5962 ( .DIN(n4726), .Q(n4904) );
  nnd2s1 U5963 ( .DIN1(n4890), .DIN2(n4943), .Q(n4726) );
  nnd2s1 U5964 ( .DIN1(n4892), .DIN2(n4871), .Q(n4943) );
  nnd2s1 U5965 ( .DIN1(n4120), .DIN2(n4129), .Q(n4871) );
  nnd3s1 U5966 ( .DIN1(n4715), .DIN2(n4732), .DIN3(n4730), .Q(n4129) );
  nnd4s1 U5967 ( .DIN1(n1927), .DIN2(n4896), .DIN3(n1959), .DIN4(n4944), 
        .Q(n4120) );
  nor2s1 U5968 ( .DIN1(n1962), .DIN2(n1956), .Q(n4944) );
  nnd2s1 U5969 ( .DIN1(n1953), .DIN2(n4786), .Q(n4896) );
  and3s1 U5970 ( .DIN1(n225), .DIN2(n57), .DIN3(\IDinst/opcode_of_MEM[3]), 
        .Q(n4892) );
  and2s1 U5971 ( .DIN1(n4945), .DIN2(n4946), .Q(n4890) );
  nnd4s1 U5972 ( .DIN1(n4947), .DIN2(n4948), .DIN3(n375), .DIN4(n59), 
        .Q(n4946) );
  nnd2s1 U5973 ( .DIN1(\IDinst/opcode_of_MEM[1]), .DIN2(n4949), .Q(n4948) );
  nnd2s1 U5974 ( .DIN1(\IDinst/opcode_of_MEM[0]), .DIN2(n209), .Q(n4949) );
  nnd2s1 U5975 ( .DIN1(n4950), .DIN2(n57), .Q(n4947) );
  or2s1 U5976 ( .DIN1(\IDinst/opcode_of_MEM[2]), 
        .DIN2(\IDinst/opcode_of_MEM[0]), .Q(n4950) );
  nnd3s1 U5977 ( .DIN1(n4951), .DIN2(n4952), .DIN3(n57), .Q(n4945) );
  or2s1 U5978 ( .DIN1(n4953), .DIN2(\IDinst/opcode_of_MEM[3]), .Q(n4952) );
  nnd2s1 U5979 ( .DIN1(n4953), .DIN2(n4954), .Q(n4951) );
  nnd2s1 U5980 ( .DIN1(n4955), .DIN2(n4956), .Q(n4954) );
  nnd2s1 U5981 ( .DIN1(\IDinst/opcode_of_MEM[0]), .DIN2(n225), .Q(n4956) );
  nnd2s1 U5982 ( .DIN1(\IDinst/opcode_of_MEM[3]), 
        .DIN2(\IDinst/opcode_of_MEM[1]), .Q(n4955) );
  nor2s1 U5983 ( .DIN1(n59), .DIN2(n209), .Q(n4953) );
  nnd2s1 U5984 ( .DIN1(n649), .DIN2(n439), .Q(n4852) );
  nnd2s1 U5985 ( .DIN1(n4957), .DIN2(n4958), .Q(\IDinst/n4729 ) );
  nnd2s1 U5986 ( .DIN1(n638), .DIN2(n440), .Q(n4958) );
  nnd2s1 U5987 ( .DIN1(n675), .DIN2(n271), .Q(n4957) );
  nnd4s1 U5988 ( .DIN1(n4959), .DIN2(n4960), .DIN3(n4961), .DIN4(n4962), 
        .Q(\IDinst/N999 ) );
  nnd2s1 U5989 ( .DIN1(n748), .DIN2(n4197), .Q(n4962) );
  nnd2s1 U5990 ( .DIN1(n4964), .DIN2(n4965), .Q(n4197) );
  nnd2s1 U5991 ( .DIN1(n627), .DIN2(n1998), .Q(n4965) );
  nnd2s1 U5992 ( .DIN1(\IDinst/N78 ), .DIN2(n525), .Q(n4964) );
  nnd2s1 U5993 ( .DIN1(n543), .DIN2(n264), .Q(n4961) );
  nnd2s1 U5994 ( .DIN1(n541), .DIN2(n147), .Q(n4960) );
  nnd2s1 U5995 ( .DIN1(n530), .DIN2(\NPC[7] ), .Q(n4959) );
  nnd4s1 U5996 ( .DIN1(n4966), .DIN2(n4967), .DIN3(n4968), .DIN4(n4969), 
        .Q(\IDinst/N998 ) );
  nnd2s1 U5997 ( .DIN1(n4963), .DIN2(n4198), .Q(n4969) );
  nnd2s1 U5998 ( .DIN1(n4970), .DIN2(n4971), .Q(n4198) );
  nnd2s1 U5999 ( .DIN1(n626), .DIN2(n1995), .Q(n4971) );
  nnd2s1 U6000 ( .DIN1(\IDinst/N79 ), .DIN2(n524), .Q(n4970) );
  nnd2s1 U6001 ( .DIN1(n542), .DIN2(n265), .Q(n4968) );
  nnd2s1 U6002 ( .DIN1(n540), .DIN2(n148), .Q(n4967) );
  nnd2s1 U6003 ( .DIN1(n529), .DIN2(\NPC[6] ), .Q(n4966) );
  nnd4s1 U6004 ( .DIN1(n4972), .DIN2(n4973), .DIN3(n4974), .DIN4(n4975), 
        .Q(\IDinst/N997 ) );
  nnd2s1 U6005 ( .DIN1(n748), .DIN2(n4199), .Q(n4975) );
  nnd2s1 U6006 ( .DIN1(n4976), .DIN2(n4977), .Q(n4199) );
  nnd2s1 U6007 ( .DIN1(n627), .DIN2(n1992), .Q(n4977) );
  nnd2s1 U6008 ( .DIN1(\IDinst/N80 ), .DIN2(n525), .Q(n4976) );
  nnd2s1 U6009 ( .DIN1(n543), .DIN2(n266), .Q(n4974) );
  nnd2s1 U6010 ( .DIN1(n541), .DIN2(n149), .Q(n4973) );
  nnd2s1 U6011 ( .DIN1(n530), .DIN2(\NPC[5] ), .Q(n4972) );
  nnd4s1 U6012 ( .DIN1(n4978), .DIN2(n4979), .DIN3(n4980), .DIN4(n4981), 
        .Q(\IDinst/N996 ) );
  nnd2s1 U6013 ( .DIN1(n4963), .DIN2(n4200), .Q(n4981) );
  nnd2s1 U6014 ( .DIN1(n4982), .DIN2(n4983), .Q(n4200) );
  nnd2s1 U6015 ( .DIN1(n626), .DIN2(n1989), .Q(n4983) );
  nnd2s1 U6016 ( .DIN1(\IDinst/N81 ), .DIN2(n524), .Q(n4982) );
  nnd2s1 U6017 ( .DIN1(n542), .DIN2(n267), .Q(n4980) );
  nnd2s1 U6018 ( .DIN1(n540), .DIN2(n150), .Q(n4979) );
  nnd2s1 U6019 ( .DIN1(n529), .DIN2(\NPC[4] ), .Q(n4978) );
  nnd4s1 U6020 ( .DIN1(n4984), .DIN2(n4985), .DIN3(n4986), .DIN4(n4987), 
        .Q(\IDinst/N995 ) );
  nnd2s1 U6021 ( .DIN1(n748), .DIN2(n4201), .Q(n4987) );
  nnd2s1 U6022 ( .DIN1(n4988), .DIN2(n4989), .Q(n4201) );
  nnd2s1 U6023 ( .DIN1(n627), .DIN2(n1986), .Q(n4989) );
  nnd2s1 U6024 ( .DIN1(\IDinst/N82 ), .DIN2(n525), .Q(n4988) );
  nnd2s1 U6025 ( .DIN1(n543), .DIN2(n268), .Q(n4986) );
  nnd2s1 U6026 ( .DIN1(n541), .DIN2(n151), .Q(n4985) );
  nnd2s1 U6027 ( .DIN1(n530), .DIN2(\NPC[3] ), .Q(n4984) );
  nnd4s1 U6028 ( .DIN1(n4990), .DIN2(n4991), .DIN3(n4992), .DIN4(n4993), 
        .Q(\IDinst/N994 ) );
  nnd2s1 U6029 ( .DIN1(n4963), .DIN2(n4202), .Q(n4993) );
  nnd2s1 U6030 ( .DIN1(n4994), .DIN2(n4995), .Q(n4202) );
  nnd2s1 U6031 ( .DIN1(n626), .DIN2(n1983), .Q(n4995) );
  nnd2s1 U6032 ( .DIN1(\IDinst/N83 ), .DIN2(n524), .Q(n4994) );
  nnd2s1 U6033 ( .DIN1(n542), .DIN2(n269), .Q(n4992) );
  nnd2s1 U6034 ( .DIN1(n540), .DIN2(n152), .Q(n4991) );
  nnd2s1 U6035 ( .DIN1(n529), .DIN2(\NPC[2] ), .Q(n4990) );
  nnd4s1 U6036 ( .DIN1(n4996), .DIN2(n4997), .DIN3(n4998), .DIN4(n4999), 
        .Q(\IDinst/N993 ) );
  nnd2s1 U6037 ( .DIN1(n748), .DIN2(n4203), .Q(n4999) );
  nnd2s1 U6038 ( .DIN1(n5000), .DIN2(n5001), .Q(n4203) );
  nnd2s1 U6039 ( .DIN1(n627), .DIN2(n1980), .Q(n5001) );
  nnd2s1 U6040 ( .DIN1(\IDinst/N84 ), .DIN2(n525), .Q(n5000) );
  nnd2s1 U6041 ( .DIN1(n543), .DIN2(n270), .Q(n4998) );
  nnd2s1 U6042 ( .DIN1(n541), .DIN2(n153), .Q(n4997) );
  nnd2s1 U6043 ( .DIN1(n530), .DIN2(\IFinst/N8 ), .Q(n4996) );
  nnd4s1 U6044 ( .DIN1(n5002), .DIN2(n5003), .DIN3(n5004), .DIN4(n5005), 
        .Q(\IDinst/N992 ) );
  nnd2s1 U6045 ( .DIN1(n4963), .DIN2(n4204), .Q(n5005) );
  nnd2s1 U6046 ( .DIN1(n5006), .DIN2(n5007), .Q(n4204) );
  nnd2s1 U6047 ( .DIN1(n626), .DIN2(n1977), .Q(n5007) );
  nnd2s1 U6048 ( .DIN1(\IDinst/N85 ), .DIN2(n524), .Q(n5006) );
  nnd2s1 U6049 ( .DIN1(n542), .DIN2(n271), .Q(n5004) );
  nnd2s1 U6050 ( .DIN1(n540), .DIN2(n154), .Q(n5003) );
  nnd2s1 U6051 ( .DIN1(n529), .DIN2(\IFinst/N7 ), .Q(n5002) );
  nnd2s1 U6052 ( .DIN1(n5008), .DIN2(n5009), .Q(\IDinst/N1055 ) );
  nnd2s1 U6053 ( .DIN1(\IDinst/N89 ), .DIN2(n537), .Q(n5009) );
  nnd2s1 U6054 ( .DIN1(n770), .DIN2(n155), .Q(n5008) );
  nnd2s1 U6055 ( .DIN1(n5011), .DIN2(n5012), .Q(\IDinst/N1054 ) );
  nnd2s1 U6056 ( .DIN1(\IDinst/N90 ), .DIN2(n536), .Q(n5012) );
  nnd2s1 U6057 ( .DIN1(n5010), .DIN2(n157), .Q(n5011) );
  nnd2s1 U6058 ( .DIN1(n5013), .DIN2(n5014), .Q(\IDinst/N1053 ) );
  nnd2s1 U6059 ( .DIN1(\IDinst/N91 ), .DIN2(n537), .Q(n5014) );
  nnd2s1 U6060 ( .DIN1(n770), .DIN2(n159), .Q(n5013) );
  nnd2s1 U6061 ( .DIN1(n5015), .DIN2(n5016), .Q(\IDinst/N1052 ) );
  nnd2s1 U6062 ( .DIN1(\IDinst/N92 ), .DIN2(n536), .Q(n5016) );
  nnd2s1 U6063 ( .DIN1(n5010), .DIN2(n161), .Q(n5015) );
  nnd2s1 U6064 ( .DIN1(n5017), .DIN2(n5018), .Q(\IDinst/N1051 ) );
  nnd2s1 U6065 ( .DIN1(\IDinst/N93 ), .DIN2(n537), .Q(n5018) );
  nnd2s1 U6066 ( .DIN1(n770), .DIN2(n163), .Q(n5017) );
  nnd2s1 U6067 ( .DIN1(n5019), .DIN2(n5020), .Q(\IDinst/N1050 ) );
  nnd2s1 U6068 ( .DIN1(\IDinst/N94 ), .DIN2(n536), .Q(n5020) );
  nnd2s1 U6069 ( .DIN1(n5010), .DIN2(n165), .Q(n5019) );
  nnd2s1 U6070 ( .DIN1(n5021), .DIN2(n5022), .Q(\IDinst/N1049 ) );
  nnd2s1 U6071 ( .DIN1(\IDinst/N95 ), .DIN2(n537), .Q(n5022) );
  nnd2s1 U6072 ( .DIN1(n770), .DIN2(n167), .Q(n5021) );
  nnd2s1 U6073 ( .DIN1(n5023), .DIN2(n5024), .Q(\IDinst/N1048 ) );
  nnd2s1 U6074 ( .DIN1(\IDinst/N96 ), .DIN2(n536), .Q(n5024) );
  nnd2s1 U6075 ( .DIN1(n5010), .DIN2(n169), .Q(n5023) );
  nnd2s1 U6076 ( .DIN1(n5025), .DIN2(n5026), .Q(\IDinst/N1047 ) );
  nnd2s1 U6077 ( .DIN1(\IDinst/N97 ), .DIN2(n537), .Q(n5026) );
  nnd2s1 U6078 ( .DIN1(n770), .DIN2(n171), .Q(n5025) );
  nnd2s1 U6079 ( .DIN1(n5027), .DIN2(n5028), .Q(\IDinst/N1046 ) );
  nnd2s1 U6080 ( .DIN1(\IDinst/N98 ), .DIN2(n536), .Q(n5028) );
  nnd2s1 U6081 ( .DIN1(n5010), .DIN2(n173), .Q(n5027) );
  nnd2s1 U6082 ( .DIN1(n5029), .DIN2(n5030), .Q(\IDinst/N1045 ) );
  nnd2s1 U6083 ( .DIN1(\IDinst/N99 ), .DIN2(n537), .Q(n5030) );
  nnd2s1 U6084 ( .DIN1(n770), .DIN2(n175), .Q(n5029) );
  nnd2s1 U6085 ( .DIN1(n5031), .DIN2(n5032), .Q(\IDinst/N1044 ) );
  nnd2s1 U6086 ( .DIN1(\IDinst/N100 ), .DIN2(n536), .Q(n5032) );
  nnd2s1 U6087 ( .DIN1(n5010), .DIN2(n177), .Q(n5031) );
  nnd2s1 U6088 ( .DIN1(n5033), .DIN2(n5034), .Q(\IDinst/N1043 ) );
  nnd2s1 U6089 ( .DIN1(\IDinst/N101 ), .DIN2(n537), .Q(n5034) );
  nnd2s1 U6090 ( .DIN1(n770), .DIN2(n179), .Q(n5033) );
  nnd2s1 U6091 ( .DIN1(n5035), .DIN2(n5036), .Q(\IDinst/N1042 ) );
  nnd2s1 U6092 ( .DIN1(\IDinst/N102 ), .DIN2(n536), .Q(n5036) );
  nnd2s1 U6093 ( .DIN1(n5010), .DIN2(n181), .Q(n5035) );
  nnd2s1 U6094 ( .DIN1(n5037), .DIN2(n5038), .Q(\IDinst/N1041 ) );
  nnd2s1 U6095 ( .DIN1(\IDinst/N103 ), .DIN2(n537), .Q(n5038) );
  nnd2s1 U6096 ( .DIN1(n770), .DIN2(n183), .Q(n5037) );
  nnd2s1 U6097 ( .DIN1(n5039), .DIN2(n5040), .Q(\IDinst/N1040 ) );
  nnd2s1 U6098 ( .DIN1(\IDinst/N104 ), .DIN2(n536), .Q(n5040) );
  nnd2s1 U6099 ( .DIN1(n5010), .DIN2(n185), .Q(n5039) );
  nnd2s1 U6100 ( .DIN1(n5041), .DIN2(n5042), .Q(\IDinst/N1039 ) );
  nnd2s1 U6101 ( .DIN1(\IDinst/N105 ), .DIN2(n537), .Q(n5042) );
  nnd2s1 U6102 ( .DIN1(n770), .DIN2(n129), .Q(n5041) );
  nnd2s1 U6103 ( .DIN1(n5043), .DIN2(n5044), .Q(\IDinst/N1038 ) );
  nnd2s1 U6104 ( .DIN1(\IDinst/N106 ), .DIN2(n536), .Q(n5044) );
  nnd2s1 U6105 ( .DIN1(n5010), .DIN2(n188), .Q(n5043) );
  nnd2s1 U6106 ( .DIN1(n5045), .DIN2(n5046), .Q(\IDinst/N1037 ) );
  nnd2s1 U6107 ( .DIN1(\IDinst/N107 ), .DIN2(n537), .Q(n5046) );
  nnd2s1 U6108 ( .DIN1(n770), .DIN2(n190), .Q(n5045) );
  nnd2s1 U6109 ( .DIN1(n5047), .DIN2(n5048), .Q(\IDinst/N1036 ) );
  nnd2s1 U6110 ( .DIN1(\IDinst/N108 ), .DIN2(n536), .Q(n5048) );
  nnd2s1 U6111 ( .DIN1(n5010), .DIN2(n192), .Q(n5047) );
  nnd2s1 U6112 ( .DIN1(n5049), .DIN2(n5050), .Q(\IDinst/N1035 ) );
  nnd2s1 U6113 ( .DIN1(\IDinst/N109 ), .DIN2(n537), .Q(n5050) );
  nnd2s1 U6114 ( .DIN1(n770), .DIN2(n194), .Q(n5049) );
  nnd2s1 U6115 ( .DIN1(n5051), .DIN2(n5052), .Q(\IDinst/N1034 ) );
  nnd2s1 U6116 ( .DIN1(\IDinst/N110 ), .DIN2(n536), .Q(n5052) );
  nnd2s1 U6117 ( .DIN1(n5010), .DIN2(n196), .Q(n5051) );
  nnd2s1 U6118 ( .DIN1(n5053), .DIN2(n5054), .Q(\IDinst/N1033 ) );
  nnd2s1 U6119 ( .DIN1(\IDinst/N111 ), .DIN2(n537), .Q(n5054) );
  nnd2s1 U6120 ( .DIN1(n770), .DIN2(n198), .Q(n5053) );
  nnd2s1 U6121 ( .DIN1(n5055), .DIN2(n5056), .Q(\IDinst/N1032 ) );
  nnd2s1 U6122 ( .DIN1(\IDinst/N112 ), .DIN2(n536), .Q(n5056) );
  nnd2s1 U6123 ( .DIN1(n5010), .DIN2(n200), .Q(n5055) );
  nnd2s1 U6124 ( .DIN1(n5057), .DIN2(n5058), .Q(\IDinst/N1031 ) );
  nnd2s1 U6125 ( .DIN1(\IDinst/N113 ), .DIN2(n537), .Q(n5058) );
  nnd2s1 U6126 ( .DIN1(n770), .DIN2(n1998), .Q(n5057) );
  hi1s1 U6127 ( .DIN(n9404), .Q(n1998) );
  nnd2s1 U6128 ( .DIN1(n5059), .DIN2(n5060), .Q(\IDinst/N1030 ) );
  nnd2s1 U6129 ( .DIN1(\IDinst/N114 ), .DIN2(n536), .Q(n5060) );
  nnd2s1 U6130 ( .DIN1(n5010), .DIN2(n1995), .Q(n5059) );
  hi1s1 U6131 ( .DIN(n9399), .Q(n1995) );
  nnd2s1 U6132 ( .DIN1(n5061), .DIN2(n5062), .Q(\IDinst/N1029 ) );
  nnd2s1 U6133 ( .DIN1(\IDinst/N115 ), .DIN2(n537), .Q(n5062) );
  nnd2s1 U6134 ( .DIN1(n770), .DIN2(n1992), .Q(n5061) );
  hi1s1 U6135 ( .DIN(n9398), .Q(n1992) );
  nnd2s1 U6136 ( .DIN1(n5063), .DIN2(n5064), .Q(\IDinst/N1028 ) );
  nnd2s1 U6137 ( .DIN1(\IDinst/N116 ), .DIN2(n536), .Q(n5064) );
  nnd2s1 U6138 ( .DIN1(n5010), .DIN2(n1989), .Q(n5063) );
  hi1s1 U6139 ( .DIN(n9397), .Q(n1989) );
  nnd2s1 U6140 ( .DIN1(n5065), .DIN2(n5066), .Q(\IDinst/N1027 ) );
  nnd2s1 U6141 ( .DIN1(\IDinst/N117 ), .DIN2(n537), .Q(n5066) );
  nnd2s1 U6142 ( .DIN1(n770), .DIN2(n1986), .Q(n5065) );
  hi1s1 U6143 ( .DIN(n9396), .Q(n1986) );
  nnd2s1 U6144 ( .DIN1(n5067), .DIN2(n5068), .Q(\IDinst/N1026 ) );
  nnd2s1 U6145 ( .DIN1(\IDinst/N118 ), .DIN2(n536), .Q(n5068) );
  nnd2s1 U6146 ( .DIN1(n5010), .DIN2(n1983), .Q(n5067) );
  hi1s1 U6147 ( .DIN(n9395), .Q(n1983) );
  nnd2s1 U6148 ( .DIN1(n5069), .DIN2(n5070), .Q(\IDinst/N1025 ) );
  nnd2s1 U6149 ( .DIN1(\IDinst/N119 ), .DIN2(n537), .Q(n5070) );
  nnd2s1 U6150 ( .DIN1(n770), .DIN2(n1980), .Q(n5069) );
  hi1s1 U6151 ( .DIN(n9394), .Q(n1980) );
  nnd2s1 U6152 ( .DIN1(n5071), .DIN2(n5072), .Q(\IDinst/N1024 ) );
  nnd2s1 U6153 ( .DIN1(\IDinst/N120 ), .DIN2(n536), .Q(n5072) );
  nnd2s1 U6154 ( .DIN1(n5010), .DIN2(n1977), .Q(n5071) );
  hi1s1 U6155 ( .DIN(n9393), .Q(n1977) );
  nor2s1 U6156 ( .DIN1(n5073), .DIN2(n5075), .Q(n5010) );
  nnd4s1 U6157 ( .DIN1(n729), .DIN2(n5077), .DIN3(reg_write_MEM), .DIN4(n5078), 
        .Q(n5073) );
  and4s1 U6158 ( .DIN1(n713), .DIN2(n5080), .DIN3(n5081), .DIN4(n4913), 
        .Q(n5078) );
  nnd4s1 U6159 ( .DIN1(n634), .DIN2(n683), .DIN3(n5082), .DIN4(n1364), 
        .Q(n4913) );
  nor2s1 U6160 ( .DIN1(n1198), .DIN2(n1312), .Q(n5082) );
  xnr2s1 U6161 ( .DIN1(\IDinst/n1433 ), .DIN2(n1238), .Q(n5081) );
  nnd2s1 U6162 ( .DIN1(n5083), .DIN2(n5084), .Q(\IDinst/N44 ) );
  nnd2s1 U6163 ( .DIN1(n9453), .DIN2(n272), .Q(n5084) );
  nnd2s1 U6164 ( .DIN1(n528), .DIN2(n273), .Q(n5083) );
  xnr2s1 U6165 ( .DIN1(\IDinst/n1432 ), .DIN2(n1332), .Q(n5080) );
  nnd2s1 U6166 ( .DIN1(n5085), .DIN2(n5086), .Q(\IDinst/N45 ) );
  nnd2s1 U6167 ( .DIN1(n9453), .DIN2(n274), .Q(n5086) );
  nnd2s1 U6168 ( .DIN1(n528), .DIN2(n275), .Q(n5085) );
  nnd2s1 U6169 ( .DIN1(n5087), .DIN2(n5088), .Q(\IDinst/N48 ) );
  nnd2s1 U6170 ( .DIN1(n551), .DIN2(n276), .Q(n5088) );
  nnd2s1 U6171 ( .DIN1(n527), .DIN2(n277), .Q(n5087) );
  xnr2s1 U6172 ( .DIN1(\IDinst/n1431 ), .DIN2(n1364), .Q(n5077) );
  nnd2s1 U6173 ( .DIN1(n5089), .DIN2(n5090), .Q(\IDinst/N46 ) );
  nnd2s1 U6174 ( .DIN1(n9453), .DIN2(n278), .Q(n5090) );
  nnd2s1 U6175 ( .DIN1(n527), .DIN2(n279), .Q(n5089) );
  nnd2s1 U6176 ( .DIN1(n551), .DIN2(n280), .Q(n5092) );
  nnd2s1 U6177 ( .DIN1(n528), .DIN2(n281), .Q(n5091) );
  nnd4s1 U6178 ( .DIN1(n5093), .DIN2(n5094), .DIN3(n5095), .DIN4(n5096), 
        .Q(\IDinst/N1023 ) );
  nnd2s1 U6179 ( .DIN1(n748), .DIN2(n4205), .Q(n5096) );
  nnd2s1 U6180 ( .DIN1(n5097), .DIN2(n5098), .Q(n4205) );
  nnd2s1 U6181 ( .DIN1(n627), .DIN2(n155), .Q(n5098) );
  nnd2s1 U6182 ( .DIN1(\IDinst/N54 ), .DIN2(n525), .Q(n5097) );
  nnd2s1 U6183 ( .DIN1(n543), .DIN2(n282), .Q(n5095) );
  nnd2s1 U6184 ( .DIN1(n541), .DIN2(n156), .Q(n5094) );
  nnd2s1 U6185 ( .DIN1(n530), .DIN2(\NPC[31] ), .Q(n5093) );
  nnd4s1 U6186 ( .DIN1(n5099), .DIN2(n5100), .DIN3(n5101), .DIN4(n5102), 
        .Q(\IDinst/N1022 ) );
  nnd2s1 U6187 ( .DIN1(n4963), .DIN2(n4206), .Q(n5102) );
  nnd2s1 U6188 ( .DIN1(n5103), .DIN2(n5104), .Q(n4206) );
  nnd2s1 U6189 ( .DIN1(n626), .DIN2(n157), .Q(n5104) );
  nnd2s1 U6190 ( .DIN1(\IDinst/N55 ), .DIN2(n524), .Q(n5103) );
  nnd2s1 U6191 ( .DIN1(n542), .DIN2(n283), .Q(n5101) );
  nnd2s1 U6192 ( .DIN1(n540), .DIN2(n158), .Q(n5100) );
  nnd2s1 U6193 ( .DIN1(n529), .DIN2(\NPC[30] ), .Q(n5099) );
  nnd4s1 U6194 ( .DIN1(n5105), .DIN2(n5106), .DIN3(n5107), .DIN4(n5108), 
        .Q(\IDinst/N1021 ) );
  nnd2s1 U6195 ( .DIN1(n748), .DIN2(n4207), .Q(n5108) );
  nnd2s1 U6196 ( .DIN1(n5109), .DIN2(n5110), .Q(n4207) );
  nnd2s1 U6197 ( .DIN1(n627), .DIN2(n159), .Q(n5110) );
  nnd2s1 U6198 ( .DIN1(\IDinst/N56 ), .DIN2(n525), .Q(n5109) );
  nnd2s1 U6199 ( .DIN1(n543), .DIN2(n284), .Q(n5107) );
  nnd2s1 U6200 ( .DIN1(n541), .DIN2(n160), .Q(n5106) );
  nnd2s1 U6201 ( .DIN1(n530), .DIN2(\NPC[29] ), .Q(n5105) );
  nnd4s1 U6202 ( .DIN1(n5111), .DIN2(n5112), .DIN3(n5113), .DIN4(n5114), 
        .Q(\IDinst/N1020 ) );
  nnd2s1 U6203 ( .DIN1(n4963), .DIN2(n4208), .Q(n5114) );
  nnd2s1 U6204 ( .DIN1(n5115), .DIN2(n5116), .Q(n4208) );
  nnd2s1 U6205 ( .DIN1(n626), .DIN2(n161), .Q(n5116) );
  nnd2s1 U6206 ( .DIN1(\IDinst/N57 ), .DIN2(n524), .Q(n5115) );
  nnd2s1 U6207 ( .DIN1(n542), .DIN2(n285), .Q(n5113) );
  nnd2s1 U6208 ( .DIN1(n540), .DIN2(n162), .Q(n5112) );
  nnd2s1 U6209 ( .DIN1(n529), .DIN2(\NPC[28] ), .Q(n5111) );
  nnd4s1 U6210 ( .DIN1(n5117), .DIN2(n5118), .DIN3(n5119), .DIN4(n5120), 
        .Q(\IDinst/N1019 ) );
  nnd2s1 U6211 ( .DIN1(n748), .DIN2(n4209), .Q(n5120) );
  nnd2s1 U6212 ( .DIN1(n5121), .DIN2(n5122), .Q(n4209) );
  nnd2s1 U6213 ( .DIN1(n627), .DIN2(n163), .Q(n5122) );
  nnd2s1 U6214 ( .DIN1(\IDinst/N58 ), .DIN2(n525), .Q(n5121) );
  nnd2s1 U6215 ( .DIN1(n543), .DIN2(n286), .Q(n5119) );
  nnd2s1 U6216 ( .DIN1(n541), .DIN2(n164), .Q(n5118) );
  nnd2s1 U6217 ( .DIN1(n530), .DIN2(\NPC[27] ), .Q(n5117) );
  nnd4s1 U6218 ( .DIN1(n5123), .DIN2(n5124), .DIN3(n5125), .DIN4(n5126), 
        .Q(\IDinst/N1018 ) );
  nnd2s1 U6219 ( .DIN1(n4963), .DIN2(n4210), .Q(n5126) );
  nnd2s1 U6220 ( .DIN1(n5127), .DIN2(n5128), .Q(n4210) );
  nnd2s1 U6221 ( .DIN1(n626), .DIN2(n165), .Q(n5128) );
  nnd2s1 U6222 ( .DIN1(\IDinst/N59 ), .DIN2(n524), .Q(n5127) );
  nnd2s1 U6223 ( .DIN1(n542), .DIN2(n287), .Q(n5125) );
  nnd2s1 U6224 ( .DIN1(n540), .DIN2(n166), .Q(n5124) );
  nnd2s1 U6225 ( .DIN1(n529), .DIN2(\NPC[26] ), .Q(n5123) );
  nnd4s1 U6226 ( .DIN1(n5129), .DIN2(n5130), .DIN3(n5131), .DIN4(n5132), 
        .Q(\IDinst/N1017 ) );
  nnd2s1 U6227 ( .DIN1(n748), .DIN2(n4211), .Q(n5132) );
  nnd2s1 U6228 ( .DIN1(n5133), .DIN2(n5134), .Q(n4211) );
  nnd2s1 U6229 ( .DIN1(n627), .DIN2(n167), .Q(n5134) );
  nnd2s1 U6230 ( .DIN1(\IDinst/N60 ), .DIN2(n525), .Q(n5133) );
  nnd2s1 U6231 ( .DIN1(n543), .DIN2(n288), .Q(n5131) );
  nnd2s1 U6232 ( .DIN1(n541), .DIN2(n168), .Q(n5130) );
  nnd2s1 U6233 ( .DIN1(n530), .DIN2(\NPC[25] ), .Q(n5129) );
  nnd4s1 U6234 ( .DIN1(n5135), .DIN2(n5136), .DIN3(n5137), .DIN4(n5138), 
        .Q(\IDinst/N1016 ) );
  nnd2s1 U6235 ( .DIN1(n4963), .DIN2(n4212), .Q(n5138) );
  nnd2s1 U6236 ( .DIN1(n5139), .DIN2(n5140), .Q(n4212) );
  nnd2s1 U6237 ( .DIN1(n626), .DIN2(n169), .Q(n5140) );
  nnd2s1 U6238 ( .DIN1(\IDinst/N61 ), .DIN2(n524), .Q(n5139) );
  nnd2s1 U6239 ( .DIN1(n542), .DIN2(n289), .Q(n5137) );
  nnd2s1 U6240 ( .DIN1(n540), .DIN2(n170), .Q(n5136) );
  nnd2s1 U6241 ( .DIN1(n529), .DIN2(\NPC[24] ), .Q(n5135) );
  nnd4s1 U6242 ( .DIN1(n5141), .DIN2(n5142), .DIN3(n5143), .DIN4(n5144), 
        .Q(\IDinst/N1015 ) );
  nnd2s1 U6243 ( .DIN1(n748), .DIN2(n4177), .Q(n5144) );
  nnd2s1 U6244 ( .DIN1(n5145), .DIN2(n5146), .Q(n4177) );
  nnd2s1 U6245 ( .DIN1(n627), .DIN2(n171), .Q(n5146) );
  nnd2s1 U6246 ( .DIN1(\IDinst/N62 ), .DIN2(n525), .Q(n5145) );
  nnd2s1 U6247 ( .DIN1(n543), .DIN2(n290), .Q(n5143) );
  nnd2s1 U6248 ( .DIN1(n541), .DIN2(n172), .Q(n5142) );
  nnd2s1 U6249 ( .DIN1(n530), .DIN2(\NPC[23] ), .Q(n5141) );
  nnd4s1 U6250 ( .DIN1(n5147), .DIN2(n5148), .DIN3(n5149), .DIN4(n5150), 
        .Q(\IDinst/N1014 ) );
  nnd2s1 U6251 ( .DIN1(n4963), .DIN2(n4178), .Q(n5150) );
  nnd2s1 U6252 ( .DIN1(n5151), .DIN2(n5152), .Q(n4178) );
  nnd2s1 U6253 ( .DIN1(n626), .DIN2(n173), .Q(n5152) );
  nnd2s1 U6254 ( .DIN1(\IDinst/N63 ), .DIN2(n524), .Q(n5151) );
  nnd2s1 U6255 ( .DIN1(n542), .DIN2(n291), .Q(n5149) );
  nnd2s1 U6256 ( .DIN1(n540), .DIN2(n174), .Q(n5148) );
  nnd2s1 U6257 ( .DIN1(n529), .DIN2(\NPC[22] ), .Q(n5147) );
  nnd4s1 U6258 ( .DIN1(n5153), .DIN2(n5154), .DIN3(n5155), .DIN4(n5156), 
        .Q(\IDinst/N1013 ) );
  nnd2s1 U6259 ( .DIN1(n748), .DIN2(n4179), .Q(n5156) );
  nnd2s1 U6260 ( .DIN1(n5157), .DIN2(n5158), .Q(n4179) );
  nnd2s1 U6261 ( .DIN1(n627), .DIN2(n175), .Q(n5158) );
  nnd2s1 U6262 ( .DIN1(\IDinst/N64 ), .DIN2(n525), .Q(n5157) );
  nnd2s1 U6263 ( .DIN1(n543), .DIN2(n292), .Q(n5155) );
  nnd2s1 U6264 ( .DIN1(n541), .DIN2(n176), .Q(n5154) );
  nnd2s1 U6265 ( .DIN1(n530), .DIN2(\NPC[21] ), .Q(n5153) );
  nnd4s1 U6266 ( .DIN1(n5159), .DIN2(n5160), .DIN3(n5161), .DIN4(n5162), 
        .Q(\IDinst/N1012 ) );
  nnd2s1 U6267 ( .DIN1(n4963), .DIN2(n4180), .Q(n5162) );
  nnd2s1 U6268 ( .DIN1(n5163), .DIN2(n5164), .Q(n4180) );
  nnd2s1 U6269 ( .DIN1(n626), .DIN2(n177), .Q(n5164) );
  nnd2s1 U6270 ( .DIN1(\IDinst/N65 ), .DIN2(n524), .Q(n5163) );
  nnd2s1 U6271 ( .DIN1(n542), .DIN2(n293), .Q(n5161) );
  nnd2s1 U6272 ( .DIN1(n540), .DIN2(n178), .Q(n5160) );
  nnd2s1 U6273 ( .DIN1(n529), .DIN2(\NPC[20] ), .Q(n5159) );
  nnd4s1 U6274 ( .DIN1(n5165), .DIN2(n5166), .DIN3(n5167), .DIN4(n5168), 
        .Q(\IDinst/N1011 ) );
  nnd2s1 U6275 ( .DIN1(n748), .DIN2(n4181), .Q(n5168) );
  nnd2s1 U6276 ( .DIN1(n5169), .DIN2(n5170), .Q(n4181) );
  nnd2s1 U6277 ( .DIN1(n627), .DIN2(n179), .Q(n5170) );
  nnd2s1 U6278 ( .DIN1(\IDinst/N66 ), .DIN2(n525), .Q(n5169) );
  nnd2s1 U6279 ( .DIN1(n543), .DIN2(n294), .Q(n5167) );
  nnd2s1 U6280 ( .DIN1(n541), .DIN2(n180), .Q(n5166) );
  nnd2s1 U6281 ( .DIN1(n530), .DIN2(\NPC[19] ), .Q(n5165) );
  nnd4s1 U6282 ( .DIN1(n5171), .DIN2(n5172), .DIN3(n5173), .DIN4(n5174), 
        .Q(\IDinst/N1010 ) );
  nnd2s1 U6283 ( .DIN1(n4963), .DIN2(n4182), .Q(n5174) );
  nnd2s1 U6284 ( .DIN1(n5175), .DIN2(n5176), .Q(n4182) );
  nnd2s1 U6285 ( .DIN1(n626), .DIN2(n181), .Q(n5176) );
  nnd2s1 U6286 ( .DIN1(\IDinst/N67 ), .DIN2(n524), .Q(n5175) );
  nnd2s1 U6287 ( .DIN1(n542), .DIN2(n295), .Q(n5173) );
  nnd2s1 U6288 ( .DIN1(n540), .DIN2(n182), .Q(n5172) );
  nnd2s1 U6289 ( .DIN1(n529), .DIN2(\NPC[18] ), .Q(n5171) );
  nnd4s1 U6290 ( .DIN1(n5177), .DIN2(n5178), .DIN3(n5179), .DIN4(n5180), 
        .Q(\IDinst/N1009 ) );
  nnd2s1 U6291 ( .DIN1(n748), .DIN2(n4183), .Q(n5180) );
  nnd2s1 U6292 ( .DIN1(n5181), .DIN2(n5182), .Q(n4183) );
  nnd2s1 U6293 ( .DIN1(n627), .DIN2(n183), .Q(n5182) );
  nnd2s1 U6294 ( .DIN1(\IDinst/N68 ), .DIN2(n525), .Q(n5181) );
  nnd2s1 U6295 ( .DIN1(n543), .DIN2(n296), .Q(n5179) );
  nnd2s1 U6296 ( .DIN1(n541), .DIN2(n184), .Q(n5178) );
  nnd2s1 U6297 ( .DIN1(n530), .DIN2(\NPC[17] ), .Q(n5177) );
  nnd4s1 U6298 ( .DIN1(n5183), .DIN2(n5184), .DIN3(n5185), .DIN4(n5186), 
        .Q(\IDinst/N1008 ) );
  nnd2s1 U6299 ( .DIN1(n4963), .DIN2(n4184), .Q(n5186) );
  nnd2s1 U6300 ( .DIN1(n5187), .DIN2(n5188), .Q(n4184) );
  nnd2s1 U6301 ( .DIN1(n626), .DIN2(n185), .Q(n5188) );
  nnd2s1 U6302 ( .DIN1(\IDinst/N69 ), .DIN2(n524), .Q(n5187) );
  nnd2s1 U6303 ( .DIN1(n542), .DIN2(n297), .Q(n5185) );
  nnd2s1 U6304 ( .DIN1(n540), .DIN2(n186), .Q(n5184) );
  nnd2s1 U6305 ( .DIN1(n529), .DIN2(\NPC[16] ), .Q(n5183) );
  nnd4s1 U6306 ( .DIN1(n5189), .DIN2(n5190), .DIN3(n5191), .DIN4(n5192), 
        .Q(\IDinst/N1007 ) );
  nnd2s1 U6307 ( .DIN1(n748), .DIN2(n4185), .Q(n5192) );
  nnd2s1 U6308 ( .DIN1(n5193), .DIN2(n5194), .Q(n4185) );
  nnd2s1 U6309 ( .DIN1(n627), .DIN2(n129), .Q(n5194) );
  nnd2s1 U6310 ( .DIN1(\IDinst/N70 ), .DIN2(n525), .Q(n5193) );
  nnd2s1 U6311 ( .DIN1(n543), .DIN2(n298), .Q(n5191) );
  nnd2s1 U6312 ( .DIN1(n541), .DIN2(n187), .Q(n5190) );
  nnd2s1 U6313 ( .DIN1(n530), .DIN2(\NPC[15] ), .Q(n5189) );
  nnd4s1 U6314 ( .DIN1(n5195), .DIN2(n5196), .DIN3(n5197), .DIN4(n5198), 
        .Q(\IDinst/N1006 ) );
  nnd2s1 U6315 ( .DIN1(n4963), .DIN2(n4186), .Q(n5198) );
  nnd2s1 U6316 ( .DIN1(n5199), .DIN2(n5200), .Q(n4186) );
  nnd2s1 U6317 ( .DIN1(n626), .DIN2(n188), .Q(n5200) );
  nnd2s1 U6318 ( .DIN1(\IDinst/N71 ), .DIN2(n524), .Q(n5199) );
  nnd2s1 U6319 ( .DIN1(n542), .DIN2(n299), .Q(n5197) );
  nnd2s1 U6320 ( .DIN1(n540), .DIN2(n189), .Q(n5196) );
  nnd2s1 U6321 ( .DIN1(n529), .DIN2(\NPC[14] ), .Q(n5195) );
  nnd4s1 U6322 ( .DIN1(n5201), .DIN2(n5202), .DIN3(n5203), .DIN4(n5204), 
        .Q(\IDinst/N1005 ) );
  nnd2s1 U6323 ( .DIN1(n748), .DIN2(n4187), .Q(n5204) );
  nnd2s1 U6324 ( .DIN1(n5205), .DIN2(n5206), .Q(n4187) );
  nnd2s1 U6325 ( .DIN1(n627), .DIN2(n190), .Q(n5206) );
  nnd2s1 U6326 ( .DIN1(\IDinst/N72 ), .DIN2(n525), .Q(n5205) );
  nnd2s1 U6327 ( .DIN1(n543), .DIN2(n300), .Q(n5203) );
  nnd2s1 U6328 ( .DIN1(n541), .DIN2(n191), .Q(n5202) );
  nnd2s1 U6329 ( .DIN1(n530), .DIN2(\NPC[13] ), .Q(n5201) );
  nnd4s1 U6330 ( .DIN1(n5207), .DIN2(n5208), .DIN3(n5209), .DIN4(n5210), 
        .Q(\IDinst/N1004 ) );
  nnd2s1 U6331 ( .DIN1(n4963), .DIN2(n4188), .Q(n5210) );
  nnd2s1 U6332 ( .DIN1(n5211), .DIN2(n5212), .Q(n4188) );
  nnd2s1 U6333 ( .DIN1(n626), .DIN2(n192), .Q(n5212) );
  nnd2s1 U6334 ( .DIN1(\IDinst/N73 ), .DIN2(n524), .Q(n5211) );
  nnd2s1 U6335 ( .DIN1(n542), .DIN2(n301), .Q(n5209) );
  nnd2s1 U6336 ( .DIN1(n540), .DIN2(n193), .Q(n5208) );
  nnd2s1 U6337 ( .DIN1(n529), .DIN2(\NPC[12] ), .Q(n5207) );
  nnd4s1 U6338 ( .DIN1(n5213), .DIN2(n5214), .DIN3(n5215), .DIN4(n5216), 
        .Q(\IDinst/N1003 ) );
  nnd2s1 U6339 ( .DIN1(n748), .DIN2(n4189), .Q(n5216) );
  nnd2s1 U6340 ( .DIN1(n5217), .DIN2(n5218), .Q(n4189) );
  nnd2s1 U6341 ( .DIN1(n627), .DIN2(n194), .Q(n5218) );
  nnd2s1 U6342 ( .DIN1(\IDinst/N74 ), .DIN2(n525), .Q(n5217) );
  nnd2s1 U6343 ( .DIN1(n543), .DIN2(n302), .Q(n5215) );
  nnd2s1 U6344 ( .DIN1(n541), .DIN2(n195), .Q(n5214) );
  nnd2s1 U6345 ( .DIN1(n530), .DIN2(\NPC[11] ), .Q(n5213) );
  nnd4s1 U6346 ( .DIN1(n5219), .DIN2(n5220), .DIN3(n5221), .DIN4(n5222), 
        .Q(\IDinst/N1002 ) );
  nnd2s1 U6347 ( .DIN1(n4963), .DIN2(n4190), .Q(n5222) );
  nnd2s1 U6348 ( .DIN1(n5223), .DIN2(n5224), .Q(n4190) );
  nnd2s1 U6349 ( .DIN1(n626), .DIN2(n196), .Q(n5224) );
  nnd2s1 U6350 ( .DIN1(\IDinst/N75 ), .DIN2(n524), .Q(n5223) );
  nnd2s1 U6351 ( .DIN1(n542), .DIN2(n303), .Q(n5221) );
  nnd2s1 U6352 ( .DIN1(n540), .DIN2(n197), .Q(n5220) );
  nnd2s1 U6353 ( .DIN1(n529), .DIN2(\NPC[10] ), .Q(n5219) );
  nnd4s1 U6354 ( .DIN1(n5225), .DIN2(n5226), .DIN3(n5227), .DIN4(n5228), 
        .Q(\IDinst/N1001 ) );
  nnd2s1 U6355 ( .DIN1(n748), .DIN2(n4191), .Q(n5228) );
  nnd2s1 U6356 ( .DIN1(n5229), .DIN2(n5230), .Q(n4191) );
  nnd2s1 U6357 ( .DIN1(n627), .DIN2(n198), .Q(n5230) );
  nnd2s1 U6358 ( .DIN1(\IDinst/N76 ), .DIN2(n525), .Q(n5229) );
  nnd2s1 U6359 ( .DIN1(n543), .DIN2(n304), .Q(n5227) );
  nnd2s1 U6360 ( .DIN1(n541), .DIN2(n199), .Q(n5226) );
  nnd2s1 U6361 ( .DIN1(n530), .DIN2(\NPC[9] ), .Q(n5225) );
  nnd4s1 U6362 ( .DIN1(n5231), .DIN2(n5232), .DIN3(n5233), .DIN4(n5234), 
        .Q(\IDinst/N1000 ) );
  nnd2s1 U6363 ( .DIN1(n4963), .DIN2(n4192), .Q(n5234) );
  nnd2s1 U6364 ( .DIN1(n5235), .DIN2(n5236), .Q(n4192) );
  nnd2s1 U6365 ( .DIN1(n626), .DIN2(n200), .Q(n5236) );
  nnd2s1 U6366 ( .DIN1(\IDinst/N77 ), .DIN2(n524), .Q(n5235) );
  and4s1 U6367 ( .DIN1(n761), .DIN2(n5241), .DIN3(n5242), .DIN4(n4906), 
        .Q(n5239) );
  nnd3s1 U6368 ( .DIN1(n1133), .DIN2(n1025), .DIN3(n5243), .Q(n4906) );
  xnr2s1 U6369 ( .DIN1(\IDinst/n1433 ), .DIN2(n1025), .Q(n5242) );
  xnr2s1 U6370 ( .DIN1(\IDinst/n1432 ), .DIN2(n1133), .Q(n5241) );
  xnr2s1 U6371 ( .DIN1(\IDinst/n1431 ), .DIN2(n1181), .Q(n5238) );
  xnr2s1 U6372 ( .DIN1(\IDinst/n1430 ), .DIN2(n672), .Q(n5237) );
  nor2s1 U6373 ( .DIN1(n5075), .DIN2(n5244), .Q(n4963) );
  hi1s1 U6374 ( .DIN(n5074), .Q(n5075) );
  nnd3s1 U6375 ( .DIN1(n4936), .DIN2(n678), .DIN3(n441), .Q(n5074) );
  hi1s1 U6376 ( .DIN(n4854), .Q(n4535) );
  nor2s1 U6377 ( .DIN1(n5245), .DIN2(n4163), .Q(n4854) );
  nnd3s1 U6378 ( .DIN1(n4163), .DIN2(n5246), .DIN3(n4164), .Q(n4936) );
  nnd2s1 U6379 ( .DIN1(n4716), .DIN2(n4715), .Q(n5246) );
  hi1s1 U6380 ( .DIN(n4124), .Q(n4716) );
  nnd2s1 U6381 ( .DIN1(n4732), .DIN2(n1962), .Q(n4124) );
  and2s1 U6382 ( .DIN1(n4786), .DIN2(n5247), .Q(n4732) );
  and2s1 U6383 ( .DIN1(n5248), .DIN2(n5249), .Q(n4163) );
  nnd3s1 U6384 ( .DIN1(\IDinst/n1444 ), .DIN2(\IDinst/n1440 ), .DIN3(INT), 
        .Q(n5249) );
  nnd2s1 U6385 ( .DIN1(n5247), .DIN2(n4901), .Q(n5248) );
  nnd2s1 U6386 ( .DIN1(n542), .DIN2(n305), .Q(n5233) );
  nnd2s1 U6387 ( .DIN1(n540), .DIN2(n201), .Q(n5232) );
  nnd2s1 U6388 ( .DIN1(n5250), .DIN2(n5251), .Q(\IDinst/N40 ) );
  nnd2s1 U6389 ( .DIN1(n9453), .DIN2(n306), .Q(n5251) );
  nnd2s1 U6390 ( .DIN1(n528), .DIN2(n307), .Q(n5250) );
  nnd2s1 U6391 ( .DIN1(n5252), .DIN2(n5253), .Q(\IDinst/N39 ) );
  nnd2s1 U6392 ( .DIN1(n551), .DIN2(n308), .Q(n5253) );
  nnd2s1 U6393 ( .DIN1(n527), .DIN2(n309), .Q(n5252) );
  and3s1 U6394 ( .DIN1(n670), .DIN2(n1183), .DIN3(n635), .Q(n5243) );
  nnd2s1 U6395 ( .DIN1(n5254), .DIN2(n5255), .Q(\IDinst/N43 ) );
  nnd2s1 U6396 ( .DIN1(n550), .DIN2(n310), .Q(n5255) );
  nnd2s1 U6397 ( .DIN1(n527), .DIN2(n311), .Q(n5254) );
  nnd2s1 U6398 ( .DIN1(n5256), .DIN2(n5257), .Q(\IDinst/N41 ) );
  nnd2s1 U6399 ( .DIN1(n9453), .DIN2(n312), .Q(n5257) );
  nnd2s1 U6400 ( .DIN1(n528), .DIN2(n313), .Q(n5256) );
  nnd2s1 U6401 ( .DIN1(n551), .DIN2(n314), .Q(n5259) );
  nnd2s1 U6402 ( .DIN1(n528), .DIN2(n315), .Q(n5258) );
  and4s1 U6403 ( .DIN1(n4715), .DIN2(n4901), .DIN3(n5260), .DIN4(n4785), 
        .Q(n5244) );
  nor2s1 U6404 ( .DIN1(n4783), .DIN2(n1956), .Q(n5260) );
  hi1s1 U6405 ( .DIN(n1953), .Q(n4715) );
  nnd2s1 U6406 ( .DIN1(n529), .DIN2(\NPC[8] ), .Q(n5231) );
  hi1s1 U6407 ( .DIN(n5245), .Q(n4164) );
  nnd2s1 U6408 ( .DIN1(n4729), .DIN2(n4733), .Q(n5245) );
  nnd2s1 U6409 ( .DIN1(n5261), .DIN2(n4901), .Q(n4733) );
  nor2s1 U6410 ( .DIN1(n4730), .DIN2(n4786), .Q(n4901) );
  hi1s1 U6411 ( .DIN(n1950), .Q(n4786) );
  nnd3s1 U6412 ( .DIN1(n5261), .DIN2(n1950), .DIN3(n4730), .Q(n4729) );
  hi1s1 U6413 ( .DIN(n1962), .Q(n4730) );
  nnd2s1 U6414 ( .DIN1(n5262), .DIN2(n5263), .Q(n1962) );
  nnd2s1 U6415 ( .DIN1(n550), .DIN2(n316), .Q(n5263) );
  nnd2s1 U6416 ( .DIN1(n527), .DIN2(n317), .Q(n5262) );
  nnd2s1 U6417 ( .DIN1(n5264), .DIN2(n5265), .Q(n1950) );
  nnd2s1 U6418 ( .DIN1(n9453), .DIN2(n318), .Q(n5265) );
  nnd2s1 U6419 ( .DIN1(n527), .DIN2(n319), .Q(n5264) );
  and2s1 U6420 ( .DIN1(n5247), .DIN2(n1953), .Q(n5261) );
  nnd2s1 U6421 ( .DIN1(n5266), .DIN2(n5267), .Q(n1953) );
  nnd2s1 U6422 ( .DIN1(n551), .DIN2(n320), .Q(n5267) );
  nnd2s1 U6423 ( .DIN1(n528), .DIN2(n321), .Q(n5266) );
  and3s1 U6424 ( .DIN1(n4785), .DIN2(n4133), .DIN3(n4783), .Q(n5247) );
  hi1s1 U6425 ( .DIN(n1927), .Q(n4783) );
  nnd2s1 U6426 ( .DIN1(n5268), .DIN2(n5269), .Q(n1927) );
  nnd2s1 U6427 ( .DIN1(n550), .DIN2(n322), .Q(n5269) );
  nnd2s1 U6428 ( .DIN1(n528), .DIN2(n323), .Q(n5268) );
  hi1s1 U6429 ( .DIN(n1956), .Q(n4133) );
  nnd2s1 U6430 ( .DIN1(n5270), .DIN2(n5271), .Q(n1956) );
  nnd2s1 U6431 ( .DIN1(n9453), .DIN2(n324), .Q(n5271) );
  nnd2s1 U6432 ( .DIN1(n527), .DIN2(n325), .Q(n5270) );
  hi1s1 U6433 ( .DIN(n1959), .Q(n4785) );
  nnd2s1 U6434 ( .DIN1(n5272), .DIN2(n5273), .Q(n1959) );
  nnd2s1 U6435 ( .DIN1(n551), .DIN2(n326), .Q(n5273) );
  nnd2s1 U6436 ( .DIN1(n527), .DIN2(n327), .Q(n5272) );
  nnd2s1 U6437 ( .DIN1(stall), .DIN2(\IDinst/n1440 ), .Q(n5274) );
  hi1s1 U6438 ( .DIN(n1918), .Q(n4148) );
  nnd4s1 U6439 ( .DIN1(\IDinst/n1445 ), .DIN2(n9453), .DIN3(n5275), 
        .DIN4(n5276), .Q(n1918) );
  nnd2s1 U6440 ( .DIN1(\IDinst/n1440 ), .DIN2(FREEZE), .Q(n5276) );
  nnd2s1 U6441 ( .DIN1(n5277), .DIN2(n119), .Q(n5275) );
  nnd2s1 U6442 ( .DIN1(\IDinst/slot_num[1]), .DIN2(\IDinst/slot_num[0]), 
        .Q(n5277) );
  or4s1 U6443 ( .DIN1(n5278), .DIN2(n5279), .DIN3(n5280), .DIN4(n5281), 
        .Q(\EXinst/n1463 ) );
  nnd4s1 U6444 ( .DIN1(n5282), .DIN2(n5283), .DIN3(n5284), .DIN4(n5285), 
        .Q(n5281) );
  nnd2s1 U6445 ( .DIN1(n5286), .DIN2(n5287), .Q(n5285) );
  nnd2s1 U6446 ( .DIN1(n5288), .DIN2(n5289), .Q(n5286) );
  or2s1 U6447 ( .DIN1(n5290), .DIN2(n5291), .Q(n5289) );
  nnd4s1 U6448 ( .DIN1(n5292), .DIN2(n5293), .DIN3(n5294), .DIN4(n5295), 
        .Q(n5284) );
  nor2s1 U6449 ( .DIN1(n5296), .DIN2(n5297), .Q(n5295) );
  nor2s1 U6450 ( .DIN1(n5298), .DIN2(n5299), .Q(n5297) );
  and2s1 U6451 ( .DIN1(n5300), .DIN2(n5301), .Q(n5298) );
  nor2s1 U6452 ( .DIN1(n5302), .DIN2(n5303), .Q(n5296) );
  nnd2s1 U6453 ( .DIN1(n719), .DIN2(n5305), .Q(n5294) );
  nnd2s1 U6454 ( .DIN1(n5306), .DIN2(n5307), .Q(n5293) );
  nnd4s1 U6455 ( .DIN1(n5308), .DIN2(n5309), .DIN3(n5310), .DIN4(n5311), 
        .Q(n5307) );
  nnd2s1 U6456 ( .DIN1(n783), .DIN2(n79), .Q(n5311) );
  nnd2s1 U6457 ( .DIN1(n758), .DIN2(n335), .Q(n5310) );
  nnd2s1 U6458 ( .DIN1(n789), .DIN2(n717), .Q(n5309) );
  nnd2s1 U6459 ( .DIN1(n553), .DIN2(n62), .Q(n5308) );
  nnd2s1 U6460 ( .DIN1(n5315), .DIN2(n5316), .Q(n5292) );
  nnd2s1 U6461 ( .DIN1(n5317), .DIN2(n5318), .Q(n5283) );
  nnd2s1 U6462 ( .DIN1(n5319), .DIN2(n5320), .Q(n5318) );
  nnd2s1 U6463 ( .DIN1(n5321), .DIN2(n5322), .Q(n5320) );
  hi1s1 U6464 ( .DIN(n5323), .Q(n5319) );
  nnd2s1 U6465 ( .DIN1(n782), .DIN2(n5325), .Q(n5282) );
  nnd4s1 U6466 ( .DIN1(n5326), .DIN2(n5327), .DIN3(n5328), .DIN4(n5329), 
        .Q(n5325) );
  and3s1 U6467 ( .DIN1(n5330), .DIN2(n5331), .DIN3(n5332), .Q(n5329) );
  nnd2s1 U6468 ( .DIN1(n734), .DIN2(n5333), .Q(n5332) );
  nnd3s1 U6469 ( .DIN1(n5334), .DIN2(n5335), .DIN3(n5469), .Q(n5333) );
  nnd2s1 U6470 ( .DIN1(n769), .DIN2(n5337), .Q(n5335) );
  nnd2s1 U6471 ( .DIN1(reg_out_B[31]), .DIN2(n776), .Q(n5334) );
  nnd3s1 U6472 ( .DIN1(n5339), .DIN2(n5340), .DIN3(n5341), .Q(n5331) );
  nnd2s1 U6473 ( .DIN1(n5342), .DIN2(n5343), .Q(n5341) );
  nnd2s1 U6474 ( .DIN1(n387), .DIN2(n5344), .Q(n5343) );
  nnd2s1 U6475 ( .DIN1(n5345), .DIN2(n5346), .Q(n5340) );
  nnd4s1 U6476 ( .DIN1(n5347), .DIN2(n5348), .DIN3(n5349), .DIN4(n5350), 
        .Q(n5346) );
  nnd2s1 U6477 ( .DIN1(n771), .DIN2(n79), .Q(n5350) );
  nnd2s1 U6478 ( .DIN1(n531), .DIN2(n335), .Q(n5349) );
  nnd2s1 U6479 ( .DIN1(n773), .DIN2(n717), .Q(n5348) );
  nnd2s1 U6480 ( .DIN1(n755), .DIN2(n401), .Q(n5347) );
  nnd2s1 U6481 ( .DIN1(n5354), .DIN2(n808), .Q(n5339) );
  nnd3s1 U6482 ( .DIN1(n5355), .DIN2(n5356), .DIN3(n5357), .Q(n5354) );
  or2s1 U6483 ( .DIN1(n140), .DIN2(n5358), .Q(n5357) );
  or2s1 U6484 ( .DIN1(n5359), .DIN2(n5360), .Q(n5356) );
  or2s1 U6485 ( .DIN1(n208), .DIN2(n5361), .Q(n5355) );
  nnd2s1 U6486 ( .DIN1(n5362), .DIN2(n5363), .Q(n5330) );
  nnd2s1 U6487 ( .DIN1(n5364), .DIN2(n5365), .Q(n5363) );
  nnd2s1 U6488 ( .DIN1(n5336), .DIN2(n5366), .Q(n5365) );
  hi1s1 U6489 ( .DIN(n5367), .Q(n5364) );
  nnd2s1 U6490 ( .DIN1(n5368), .DIN2(reg_out_B[31]), .Q(n5328) );
  nnd2s1 U6491 ( .DIN1(n5369), .DIN2(n5370), .Q(n5327) );
  nnd3s1 U6492 ( .DIN1(n5371), .DIN2(n749), .DIN3(n5373), .Q(n5369) );
  or2s1 U6493 ( .DIN1(n5374), .DIN2(n706), .Q(n5373) );
  nnd2s1 U6494 ( .DIN1(n653), .DIN2(n5376), .Q(n5371) );
  nnd2s1 U6495 ( .DIN1(n5377), .DIN2(n5378), .Q(n5326) );
  nnd2s1 U6496 ( .DIN1(n5379), .DIN2(n5380), .Q(n5378) );
  or2s1 U6497 ( .DIN1(n5381), .DIN2(n5376), .Q(n5380) );
  nnd2s1 U6498 ( .DIN1(n5382), .DIN2(n5383), .Q(n5376) );
  nnd2s1 U6499 ( .DIN1(n5384), .DIN2(n18), .Q(n5383) );
  nnd2s1 U6500 ( .DIN1(reg_out_A[30]), .DIN2(n5385), .Q(n5384) );
  nnd2s1 U6501 ( .DIN1(n5386), .DIN2(n717), .Q(n5382) );
  nnd2s1 U6502 ( .DIN1(n620), .DIN2(n5374), .Q(n5379) );
  nnd2s1 U6503 ( .DIN1(n5387), .DIN2(n5388), .Q(n5374) );
  nnd2s1 U6504 ( .DIN1(n5389), .DIN2(n5390), .Q(n5388) );
  nnd3s1 U6505 ( .DIN1(n5391), .DIN2(n5392), .DIN3(n5393), .Q(n5280) );
  nnd2s1 U6506 ( .DIN1(n727), .DIN2(\DM_addr[31] ), .Q(n5393) );
  nnd2s1 U6507 ( .DIN1(n734), .DIN2(n5395), .Q(n5392) );
  nnd4s1 U6508 ( .DIN1(n5396), .DIN2(n5397), .DIN3(n5398), .DIN4(n5399), 
        .Q(n5395) );
  nor2s1 U6509 ( .DIN1(n5400), .DIN2(n402), .Q(n5399) );
  nnd2s1 U6510 ( .DIN1(n5401), .DIN2(n124), .Q(n5398) );
  nnd2s1 U6511 ( .DIN1(n5402), .DIN2(n5403), .Q(n5401) );
  nnd2s1 U6512 ( .DIN1(n385), .DIN2(n5291), .Q(n5403) );
  hi1s1 U6513 ( .DIN(n5405), .Q(n5402) );
  nnd2s1 U6514 ( .DIN1(n791), .DIN2(n5407), .Q(n5397) );
  nnd2s1 U6515 ( .DIN1(n5408), .DIN2(n548), .Q(n5396) );
  nnd2s1 U6516 ( .DIN1(n5409), .DIN2(n62), .Q(n5391) );
  nnd3s1 U6517 ( .DIN1(n5410), .DIN2(n5411), .DIN3(n5412), .Q(n5409) );
  nnd3s1 U6518 ( .DIN1(n9460), .DIN2(n5291), .DIN3(n385), .Q(n5412) );
  xor2s1 U6519 ( .DIN1(n744), .DIN2(n5414), .Q(n5291) );
  nor2s1 U6520 ( .DIN1(n5415), .DIN2(n5416), .Q(n5414) );
  and2s1 U6521 ( .DIN1(n5417), .DIN2(n5418), .Q(n5416) );
  nor2s1 U6522 ( .DIN1(reg_out_A[30]), .DIN2(n5419), .Q(n5415) );
  nor2s1 U6523 ( .DIN1(n5418), .DIN2(n5417), .Q(n5419) );
  nnd2s1 U6524 ( .DIN1(n549), .DIN2(n5407), .Q(n5411) );
  nnd2s1 U6525 ( .DIN1(n791), .DIN2(n5408), .Q(n5410) );
  hi1s1 U6526 ( .DIN(n5407), .Q(n5408) );
  nnd2s1 U6527 ( .DIN1(n5420), .DIN2(n5421), .Q(n5407) );
  nnd2s1 U6528 ( .DIN1(n5422), .DIN2(n717), .Q(n5421) );
  nnd2s1 U6529 ( .DIN1(n633), .DIN2(n5424), .Q(n5422) );
  nnd2s1 U6530 ( .DIN1(n5425), .DIN2(n5426), .Q(n5420) );
  nor2s1 U6531 ( .DIN1(n9460), .DIN2(n5427), .Q(n5279) );
  nor2s1 U6532 ( .DIN1(n9476), .DIN2(n5428), .Q(n5278) );
  or4s1 U6533 ( .DIN1(n5429), .DIN2(n5430), .DIN3(n5431), .DIN4(n5432), 
        .Q(\EXinst/n1462 ) );
  nnd4s1 U6534 ( .DIN1(n5433), .DIN2(n5434), .DIN3(n5435), .DIN4(n5436), 
        .Q(n5432) );
  and3s1 U6535 ( .DIN1(n5437), .DIN2(n5438), .DIN3(n5439), .Q(n5436) );
  nnd2s1 U6536 ( .DIN1(n405), .DIN2(n96), .Q(n5439) );
  nnd2s1 U6537 ( .DIN1(n782), .DIN2(n5440), .Q(n5438) );
  nnd4s1 U6538 ( .DIN1(n5441), .DIN2(n5442), .DIN3(n5443), .DIN4(n5444), 
        .Q(n5440) );
  and4s1 U6539 ( .DIN1(n5445), .DIN2(n5446), .DIN3(n5447), .DIN4(n5448), 
        .Q(n5444) );
  nnd2s1 U6540 ( .DIN1(n5449), .DIN2(n5450), .Q(n5448) );
  nnd3s1 U6541 ( .DIN1(n5451), .DIN2(n5372), .DIN3(n5452), .Q(n5449) );
  nnd2s1 U6542 ( .DIN1(n705), .DIN2(n5453), .Q(n5452) );
  nnd2s1 U6543 ( .DIN1(n656), .DIN2(n5386), .Q(n5451) );
  hi1s1 U6544 ( .DIN(n5385), .Q(n5386) );
  nnd2s1 U6545 ( .DIN1(n5454), .DIN2(n5455), .Q(n5447) );
  nnd2s1 U6546 ( .DIN1(n5456), .DIN2(n5457), .Q(n5455) );
  nnd2s1 U6547 ( .DIN1(n655), .DIN2(n5385), .Q(n5457) );
  nnd2s1 U6548 ( .DIN1(n5458), .DIN2(n5459), .Q(n5385) );
  nnd2s1 U6549 ( .DIN1(reg_out_B[29]), .DIN2(n5460), .Q(n5459) );
  nnd2s1 U6550 ( .DIN1(n5461), .DIN2(n79), .Q(n5460) );
  nnd2s1 U6551 ( .DIN1(n406), .DIN2(n5462), .Q(n5458) );
  nnd2s1 U6552 ( .DIN1(n620), .DIN2(n5389), .Q(n5456) );
  hi1s1 U6553 ( .DIN(n5453), .Q(n5389) );
  nnd2s1 U6554 ( .DIN1(n5463), .DIN2(n5464), .Q(n5453) );
  nnd2s1 U6555 ( .DIN1(n5465), .DIN2(n5466), .Q(n5464) );
  nnd2s1 U6556 ( .DIN1(n5467), .DIN2(n5468), .Q(n5446) );
  nnd2s1 U6557 ( .DIN1(reg_out_A[30]), .DIN2(n768), .Q(n5445) );
  nnd2s1 U6558 ( .DIN1(reg_out_B[30]), .DIN2(n5470), .Q(n5443) );
  nnd2s1 U6559 ( .DIN1(n723), .DIN2(n5472), .Q(n5470) );
  nnd2s1 U6560 ( .DIN1(reg_out_A[30]), .DIN2(n775), .Q(n5472) );
  nnd3s1 U6561 ( .DIN1(n5473), .DIN2(n5474), .DIN3(n769), .Q(n5442) );
  nnd2s1 U6562 ( .DIN1(n5475), .DIN2(n5476), .Q(n5474) );
  nnd3s1 U6563 ( .DIN1(n5477), .DIN2(n337), .DIN3(n5478), .Q(n5476) );
  nnd2s1 U6564 ( .DIN1(reg_out_B[5]), .DIN2(n5479), .Q(n5473) );
  nnd3s1 U6565 ( .DIN1(n714), .DIN2(n801), .DIN3(n5480), .Q(n5479) );
  nnd2s1 U6566 ( .DIN1(n5481), .DIN2(n5482), .Q(n5441) );
  nnd3s1 U6567 ( .DIN1(n5483), .DIN2(n5484), .DIN3(n204), .Q(n5482) );
  nnd2s1 U6568 ( .DIN1(n5485), .DIN2(n801), .Q(n5484) );
  nnd2s1 U6569 ( .DIN1(n5486), .DIN2(n5487), .Q(n5485) );
  nnd2s1 U6570 ( .DIN1(n741), .DIN2(n5488), .Q(n5487) );
  nnd2s1 U6571 ( .DIN1(n5489), .DIN2(n205), .Q(n5486) );
  nnd4s1 U6572 ( .DIN1(n5491), .DIN2(n5492), .DIN3(n5493), .DIN4(n5494), 
        .Q(n5489) );
  hi1s1 U6573 ( .DIN(n5495), .Q(n5494) );
  nnd2s1 U6574 ( .DIN1(n5496), .DIN2(n61), .Q(n5483) );
  nnd2s1 U6575 ( .DIN1(n5497), .DIN2(n5498), .Q(n5496) );
  nnd2s1 U6576 ( .DIN1(n742), .DIN2(n5499), .Q(n5498) );
  nnd2s1 U6577 ( .DIN1(n5500), .DIN2(n205), .Q(n5497) );
  nnd2s1 U6578 ( .DIN1(n5342), .DIN2(n5501), .Q(n5481) );
  nnd2s1 U6579 ( .DIN1(n387), .DIN2(n5502), .Q(n5501) );
  or2s1 U6580 ( .DIN1(n5428), .DIN2(n9477), .Q(n5437) );
  nnd2s1 U6581 ( .DIN1(n5394), .DIN2(\DM_addr[30] ), .Q(n5435) );
  nnd2s1 U6582 ( .DIN1(reg_out_A[30]), .DIN2(n5503), .Q(n5434) );
  nnd4s1 U6583 ( .DIN1(n5504), .DIN2(n5505), .DIN3(n5506), .DIN4(n5507), 
        .Q(n5503) );
  nor2s1 U6584 ( .DIN1(n403), .DIN2(n5508), .Q(n5507) );
  nor2s1 U6585 ( .DIN1(n5290), .DIN2(n5509), .Q(n5508) );
  nnd2s1 U6586 ( .DIN1(n5405), .DIN2(n96), .Q(n5506) );
  nnd2s1 U6587 ( .DIN1(n548), .DIN2(n5424), .Q(n5505) );
  nnd2s1 U6588 ( .DIN1(n791), .DIN2(n5425), .Q(n5504) );
  nnd2s1 U6589 ( .DIN1(n5510), .DIN2(n717), .Q(n5433) );
  nnd3s1 U6590 ( .DIN1(n5511), .DIN2(n5512), .DIN3(n5513), .Q(n5510) );
  nnd2s1 U6591 ( .DIN1(n385), .DIN2(n5509), .Q(n5513) );
  xor2s1 U6592 ( .DIN1(n5418), .DIN2(n5417), .Q(n5509) );
  xnr2s1 U6593 ( .DIN1(n9461), .DIN2(n786), .Q(n5417) );
  and2s1 U6594 ( .DIN1(n5515), .DIN2(n5516), .Q(n5418) );
  nnd2s1 U6595 ( .DIN1(n406), .DIN2(n5517), .Q(n5516) );
  or2s1 U6596 ( .DIN1(n5518), .DIN2(n5519), .Q(n5517) );
  nnd2s1 U6597 ( .DIN1(n5519), .DIN2(n5518), .Q(n5515) );
  nnd2s1 U6598 ( .DIN1(n791), .DIN2(n5424), .Q(n5512) );
  nnd2s1 U6599 ( .DIN1(n549), .DIN2(n5425), .Q(n5511) );
  hi1s1 U6600 ( .DIN(n5424), .Q(n5425) );
  nnd2s1 U6601 ( .DIN1(n5520), .DIN2(n5521), .Q(n5424) );
  nnd2s1 U6602 ( .DIN1(n406), .DIN2(n5522), .Q(n5521) );
  nnd2s1 U6603 ( .DIN1(n5523), .DIN2(n5426), .Q(n5522) );
  nnd2s1 U6604 ( .DIN1(n5423), .DIN2(n5524), .Q(n5520) );
  nnd3s1 U6605 ( .DIN1(n5525), .DIN2(n5526), .DIN3(n5527), .Q(n5431) );
  nnd2s1 U6606 ( .DIN1(n5528), .DIN2(n5529), .Q(n5527) );
  nnd3s1 U6607 ( .DIN1(n5530), .DIN2(n5531), .DIN3(n56), .Q(n5529) );
  nnd2s1 U6608 ( .DIN1(n5532), .DIN2(n735), .Q(n5531) );
  nnd2s1 U6609 ( .DIN1(n5533), .DIN2(n5534), .Q(n5532) );
  nnd2s1 U6610 ( .DIN1(n5535), .DIN2(n792), .Q(n5534) );
  nnd2s1 U6611 ( .DIN1(n29), .DIN2(n5536), .Q(n5533) );
  nnd2s1 U6612 ( .DIN1(n5537), .DIN2(n736), .Q(n5530) );
  nnd2s1 U6613 ( .DIN1(n5538), .DIN2(n5539), .Q(n5537) );
  nnd2s1 U6614 ( .DIN1(n5540), .DIN2(n792), .Q(n5539) );
  nnd2s1 U6615 ( .DIN1(n747), .DIN2(n5541), .Q(n5538) );
  nnd4s1 U6616 ( .DIN1(n5542), .DIN2(n5543), .DIN3(n5544), .DIN4(n5545), 
        .Q(n5541) );
  hi1s1 U6617 ( .DIN(n5546), .Q(n5545) );
  nnd2s1 U6618 ( .DIN1(n5547), .DIN2(n5548), .Q(n5528) );
  nnd2s1 U6619 ( .DIN1(n5301), .DIN2(n5549), .Q(n5548) );
  nnd3s1 U6620 ( .DIN1(n5550), .DIN2(n4831), .DIN3(n5551), .Q(n5526) );
  nnd3s1 U6621 ( .DIN1(n5552), .DIN2(n5553), .DIN3(n5400), .Q(n5525) );
  hi1s1 U6622 ( .DIN(n5554), .Q(n5400) );
  nnd3s1 U6623 ( .DIN1(n5555), .DIN2(n5556), .DIN3(n739), .Q(n5552) );
  nnd2s1 U6624 ( .DIN1(n736), .DIN2(n5557), .Q(n5555) );
  nor2s1 U6625 ( .DIN1(n5558), .DIN2(n5559), .Q(n5430) );
  nor2s1 U6626 ( .DIN1(n5560), .DIN2(n5288), .Q(n5429) );
  or4s1 U6627 ( .DIN1(n5561), .DIN2(n5562), .DIN3(n5563), .DIN4(n5564), 
        .Q(\EXinst/n1461 ) );
  nnd4s1 U6628 ( .DIN1(n5565), .DIN2(n5566), .DIN3(n5567), .DIN4(n5568), 
        .Q(n5564) );
  nnd3s1 U6629 ( .DIN1(n555), .DIN2(n5569), .DIN3(n5570), .Q(n5568) );
  nnd2s1 U6630 ( .DIN1(n5571), .DIN2(n5572), .Q(n5567) );
  nnd2s1 U6631 ( .DIN1(n5573), .DIN2(n5574), .Q(n5572) );
  nnd3s1 U6632 ( .DIN1(n5575), .DIN2(n5553), .DIN3(n554), .Q(n5574) );
  nnd2s1 U6633 ( .DIN1(n5554), .DIN2(n5576), .Q(n5571) );
  nnd2s1 U6634 ( .DIN1(n5577), .DIN2(n5322), .Q(n5576) );
  hi1s1 U6635 ( .DIN(n5578), .Q(n5577) );
  nnd2s1 U6636 ( .DIN1(n5579), .DIN2(n5580), .Q(n5566) );
  nnd3s1 U6637 ( .DIN1(n5581), .DIN2(n5582), .DIN3(n740), .Q(n5580) );
  nnd2s1 U6638 ( .DIN1(n5583), .DIN2(n735), .Q(n5582) );
  nnd2s1 U6639 ( .DIN1(n5584), .DIN2(n5585), .Q(n5583) );
  nnd2s1 U6640 ( .DIN1(n5586), .DIN2(n792), .Q(n5585) );
  nnd2s1 U6641 ( .DIN1(n29), .DIN2(n5587), .Q(n5584) );
  nnd2s1 U6642 ( .DIN1(n5588), .DIN2(n736), .Q(n5581) );
  nnd2s1 U6643 ( .DIN1(n5589), .DIN2(n5590), .Q(n5588) );
  nnd2s1 U6644 ( .DIN1(n5591), .DIN2(n792), .Q(n5590) );
  nnd2s1 U6645 ( .DIN1(n747), .DIN2(n5592), .Q(n5589) );
  nnd4s1 U6646 ( .DIN1(n5593), .DIN2(n5594), .DIN3(n5595), .DIN4(n5596), 
        .Q(n5592) );
  nnd2s1 U6647 ( .DIN1(n5547), .DIN2(n5597), .Q(n5579) );
  nnd2s1 U6648 ( .DIN1(n5301), .DIN2(n5598), .Q(n5597) );
  nnd2s1 U6649 ( .DIN1(n782), .DIN2(n5599), .Q(n5565) );
  nnd4s1 U6650 ( .DIN1(n5600), .DIN2(n5601), .DIN3(n5602), .DIN4(n5603), 
        .Q(n5599) );
  and4s1 U6651 ( .DIN1(n5604), .DIN2(n5605), .DIN3(n5606), .DIN4(n5607), 
        .Q(n5603) );
  nnd2s1 U6652 ( .DIN1(n5608), .DIN2(n5609), .Q(n5607) );
  nnd3s1 U6653 ( .DIN1(n5610), .DIN2(n749), .DIN3(n5611), .Q(n5608) );
  nnd2s1 U6654 ( .DIN1(n705), .DIN2(n5465), .Q(n5611) );
  nnd2s1 U6655 ( .DIN1(n654), .DIN2(n5461), .Q(n5610) );
  hi1s1 U6656 ( .DIN(n5462), .Q(n5461) );
  nnd2s1 U6657 ( .DIN1(n5612), .DIN2(n5613), .Q(n5606) );
  nnd2s1 U6658 ( .DIN1(n5614), .DIN2(n5615), .Q(n5613) );
  nnd2s1 U6659 ( .DIN1(n653), .DIN2(n5462), .Q(n5615) );
  nnd2s1 U6660 ( .DIN1(n5616), .DIN2(n5617), .Q(n5462) );
  nnd2s1 U6661 ( .DIN1(reg_out_B[28]), .DIN2(n5618), .Q(n5617) );
  nnd2s1 U6662 ( .DIN1(n5619), .DIN2(n335), .Q(n5618) );
  nnd2s1 U6663 ( .DIN1(n12), .DIN2(n5620), .Q(n5616) );
  or2s1 U6664 ( .DIN1(n5465), .DIN2(n5375), .Q(n5614) );
  nnd2s1 U6665 ( .DIN1(n5621), .DIN2(n5622), .Q(n5465) );
  nnd2s1 U6666 ( .DIN1(n5623), .DIN2(n5624), .Q(n5622) );
  nnd2s1 U6667 ( .DIN1(reg_out_B[29]), .DIN2(n5625), .Q(n5605) );
  nnd2s1 U6668 ( .DIN1(n723), .DIN2(n5626), .Q(n5625) );
  nnd2s1 U6669 ( .DIN1(n776), .DIN2(n406), .Q(n5626) );
  nnd2s1 U6670 ( .DIN1(n406), .DIN2(n767), .Q(n5604) );
  nnd2s1 U6671 ( .DIN1(n5627), .DIN2(n5628), .Q(n5602) );
  nnd3s1 U6672 ( .DIN1(n5629), .DIN2(n5630), .DIN3(n808), .Q(n5628) );
  nnd2s1 U6673 ( .DIN1(n5631), .DIN2(n337), .Q(n5630) );
  nnd2s1 U6674 ( .DIN1(n5632), .DIN2(n5633), .Q(n5631) );
  nnd2s1 U6675 ( .DIN1(n32), .DIN2(n5634), .Q(n5633) );
  nnd2s1 U6676 ( .DIN1(n5635), .DIN2(n205), .Q(n5632) );
  nnd4s1 U6677 ( .DIN1(n5636), .DIN2(n5637), .DIN3(n5638), .DIN4(n5639), 
        .Q(n5635) );
  nnd2s1 U6678 ( .DIN1(n5640), .DIN2(n438), .Q(n5629) );
  nnd2s1 U6679 ( .DIN1(n5641), .DIN2(n5642), .Q(n5640) );
  nnd2s1 U6680 ( .DIN1(n741), .DIN2(n5643), .Q(n5642) );
  nnd2s1 U6681 ( .DIN1(n5644), .DIN2(n205), .Q(n5641) );
  nnd2s1 U6682 ( .DIN1(n5342), .DIN2(n5645), .Q(n5627) );
  nnd2s1 U6683 ( .DIN1(n387), .DIN2(n5646), .Q(n5645) );
  nnd3s1 U6684 ( .DIN1(n5647), .DIN2(n5648), .DIN3(n5336), .Q(n5601) );
  nnd2s1 U6685 ( .DIN1(n5649), .DIN2(n5650), .Q(n5648) );
  nnd3s1 U6686 ( .DIN1(n5651), .DIN2(n5478), .DIN3(n628), .Q(n5650) );
  nnd2s1 U6687 ( .DIN1(reg_out_B[5]), .DIN2(n5652), .Q(n5647) );
  or2s1 U6688 ( .DIN1(n5653), .DIN2(n753), .Q(n5652) );
  nnd3s1 U6689 ( .DIN1(n628), .DIN2(n5654), .DIN3(n5468), .Q(n5600) );
  nnd3s1 U6690 ( .DIN1(n5655), .DIN2(n5656), .DIN3(n5657), .Q(n5563) );
  nnd2s1 U6691 ( .DIN1(n727), .DIN2(\DM_addr[29] ), .Q(n5657) );
  nnd2s1 U6692 ( .DIN1(n406), .DIN2(n5658), .Q(n5656) );
  or3s1 U6693 ( .DIN1(n404), .DIN2(n5659), .DIN3(n5660), .Q(n5658) );
  nnd4s1 U6694 ( .DIN1(n5661), .DIN2(n5662), .DIN3(n5663), .DIN4(n5664), 
        .Q(n5660) );
  nnd2s1 U6695 ( .DIN1(n548), .DIN2(n5524), .Q(n5664) );
  nnd2s1 U6696 ( .DIN1(n791), .DIN2(n5523), .Q(n5663) );
  nnd2s1 U6697 ( .DIN1(n5405), .DIN2(n14), .Q(n5662) );
  nnd2s1 U6698 ( .DIN1(n5665), .DIN2(n9462), .Q(n5661) );
  nor2s1 U6699 ( .DIN1(n5290), .DIN2(n5666), .Q(n5659) );
  nnd2s1 U6700 ( .DIN1(n5667), .DIN2(n79), .Q(n5655) );
  nnd4s1 U6701 ( .DIN1(n5668), .DIN2(n5669), .DIN3(n5670), .DIN4(n5671), 
        .Q(n5667) );
  nnd2s1 U6702 ( .DIN1(n791), .DIN2(n5524), .Q(n5671) );
  nnd2s1 U6703 ( .DIN1(n549), .DIN2(n5523), .Q(n5670) );
  hi1s1 U6704 ( .DIN(n5524), .Q(n5523) );
  nnd2s1 U6705 ( .DIN1(n5672), .DIN2(n5673), .Q(n5524) );
  nnd2s1 U6706 ( .DIN1(n434), .DIN2(n5674), .Q(n5673) );
  nnd2s1 U6707 ( .DIN1(n5675), .DIN2(n5426), .Q(n5674) );
  nnd2s1 U6708 ( .DIN1(n633), .DIN2(n5676), .Q(n5672) );
  nnd2s1 U6709 ( .DIN1(n385), .DIN2(n5666), .Q(n5669) );
  xor2s1 U6710 ( .DIN1(n5518), .DIN2(n5519), .Q(n5666) );
  xor2s1 U6711 ( .DIN1(n14), .DIN2(n5413), .Q(n5519) );
  nnd2s1 U6712 ( .DIN1(n5677), .DIN2(n5678), .Q(n5518) );
  nnd2s1 U6713 ( .DIN1(n12), .DIN2(n5679), .Q(n5678) );
  nnd2s1 U6714 ( .DIN1(n5680), .DIN2(n5681), .Q(n5679) );
  or2s1 U6715 ( .DIN1(n5681), .DIN2(n5680), .Q(n5677) );
  nnd2s1 U6716 ( .DIN1(n5665), .DIN2(n14), .Q(n5668) );
  nor2s1 U6717 ( .DIN1(n9462), .DIN2(n5427), .Q(n5562) );
  nor2s1 U6718 ( .DIN1(n9478), .DIN2(n5428), .Q(n5561) );
  or4s1 U6719 ( .DIN1(n5682), .DIN2(n5683), .DIN3(n5684), .DIN4(n5685), 
        .Q(\EXinst/n1460 ) );
  nnd4s1 U6720 ( .DIN1(n5686), .DIN2(n5687), .DIN3(n5688), .DIN4(n5689), 
        .Q(n5685) );
  nor2s1 U6721 ( .DIN1(n5690), .DIN2(n5691), .Q(n5689) );
  nor2s1 U6722 ( .DIN1(n9463), .DIN2(n5427), .Q(n5691) );
  nor2s1 U6723 ( .DIN1(n9479), .DIN2(n5428), .Q(n5690) );
  nnd2s1 U6724 ( .DIN1(n5394), .DIN2(\DM_addr[28] ), .Q(n5688) );
  nnd2s1 U6725 ( .DIN1(n434), .DIN2(n5692), .Q(n5687) );
  nnd4s1 U6726 ( .DIN1(n5693), .DIN2(n5694), .DIN3(n5695), .DIN4(n5696), 
        .Q(n5692) );
  nor2s1 U6727 ( .DIN1(n405), .DIN2(n5697), .Q(n5696) );
  nor2s1 U6728 ( .DIN1(n5290), .DIN2(n5698), .Q(n5697) );
  nnd2s1 U6729 ( .DIN1(n5405), .DIN2(n102), .Q(n5695) );
  nnd2s1 U6730 ( .DIN1(n548), .DIN2(n5676), .Q(n5694) );
  nnd2s1 U6731 ( .DIN1(n791), .DIN2(n5675), .Q(n5693) );
  nnd2s1 U6732 ( .DIN1(n5699), .DIN2(n335), .Q(n5686) );
  nnd3s1 U6733 ( .DIN1(n5700), .DIN2(n5701), .DIN3(n5702), .Q(n5699) );
  nnd2s1 U6734 ( .DIN1(n385), .DIN2(n5698), .Q(n5702) );
  xor2s1 U6735 ( .DIN1(n5680), .DIN2(n5681), .Q(n5698) );
  xnr2s1 U6736 ( .DIN1(n9463), .DIN2(n785), .Q(n5681) );
  and2s1 U6737 ( .DIN1(n5703), .DIN2(n5704), .Q(n5680) );
  nnd2s1 U6738 ( .DIN1(n407), .DIN2(n5705), .Q(n5704) );
  or2s1 U6739 ( .DIN1(n5706), .DIN2(n5707), .Q(n5705) );
  nnd2s1 U6740 ( .DIN1(n5707), .DIN2(n5706), .Q(n5703) );
  nnd2s1 U6741 ( .DIN1(n791), .DIN2(n5676), .Q(n5701) );
  nnd2s1 U6742 ( .DIN1(n549), .DIN2(n5675), .Q(n5700) );
  hi1s1 U6743 ( .DIN(n5676), .Q(n5675) );
  nnd2s1 U6744 ( .DIN1(n5708), .DIN2(n5709), .Q(n5676) );
  nnd2s1 U6745 ( .DIN1(n407), .DIN2(n5710), .Q(n5709) );
  nnd2s1 U6746 ( .DIN1(n5711), .DIN2(n5426), .Q(n5710) );
  nnd2s1 U6747 ( .DIN1(n5423), .DIN2(n5712), .Q(n5708) );
  nnd3s1 U6748 ( .DIN1(n5713), .DIN2(n5714), .DIN3(n5715), .Q(n5684) );
  nnd2s1 U6749 ( .DIN1(n5716), .DIN2(n5717), .Q(n5715) );
  nnd3s1 U6750 ( .DIN1(n5718), .DIN2(n5719), .DIN3(n56), .Q(n5717) );
  nnd2s1 U6751 ( .DIN1(n5720), .DIN2(n803), .Q(n5719) );
  nnd2s1 U6752 ( .DIN1(n5721), .DIN2(n5722), .Q(n5720) );
  nnd2s1 U6753 ( .DIN1(n5723), .DIN2(n792), .Q(n5722) );
  nnd2s1 U6754 ( .DIN1(n29), .DIN2(n5724), .Q(n5721) );
  nnd2s1 U6755 ( .DIN1(n5725), .DIN2(n736), .Q(n5718) );
  nnd2s1 U6756 ( .DIN1(n5726), .DIN2(n5727), .Q(n5725) );
  nnd2s1 U6757 ( .DIN1(n5728), .DIN2(n792), .Q(n5727) );
  nnd2s1 U6758 ( .DIN1(n747), .DIN2(n5729), .Q(n5726) );
  nnd4s1 U6759 ( .DIN1(n5730), .DIN2(n5731), .DIN3(n5732), .DIN4(n5733), 
        .Q(n5729) );
  nnd2s1 U6760 ( .DIN1(n5547), .DIN2(n5734), .Q(n5716) );
  nnd2s1 U6761 ( .DIN1(n5301), .DIN2(n5735), .Q(n5734) );
  nnd3s1 U6762 ( .DIN1(n5736), .DIN2(n5737), .DIN3(n5738), .Q(n5714) );
  nnd2s1 U6763 ( .DIN1(n5739), .DIN2(n5740), .Q(n5737) );
  nnd2s1 U6764 ( .DIN1(n5741), .DIN2(n4831), .Q(n5736) );
  nnd3s1 U6765 ( .DIN1(n554), .DIN2(n5742), .DIN3(n5570), .Q(n5713) );
  and2s1 U6766 ( .DIN1(n782), .DIN2(n5743), .Q(n5683) );
  nnd4s1 U6767 ( .DIN1(n5744), .DIN2(n5745), .DIN3(n5746), .DIN4(n5747), 
        .Q(n5743) );
  and4s1 U6768 ( .DIN1(n5748), .DIN2(n5749), .DIN3(n5750), .DIN4(n5751), 
        .Q(n5747) );
  nnd2s1 U6769 ( .DIN1(n5752), .DIN2(n5753), .Q(n5751) );
  nnd3s1 U6770 ( .DIN1(n5754), .DIN2(n5372), .DIN3(n5755), .Q(n5752) );
  nnd2s1 U6771 ( .DIN1(n620), .DIN2(n5624), .Q(n5755) );
  nnd2s1 U6772 ( .DIN1(n656), .DIN2(n5619), .Q(n5754) );
  hi1s1 U6773 ( .DIN(n5620), .Q(n5619) );
  nnd2s1 U6774 ( .DIN1(n5756), .DIN2(n5757), .Q(n5750) );
  nnd2s1 U6775 ( .DIN1(n5758), .DIN2(n5759), .Q(n5757) );
  nnd2s1 U6776 ( .DIN1(n655), .DIN2(n5620), .Q(n5759) );
  nnd2s1 U6777 ( .DIN1(n5760), .DIN2(n5761), .Q(n5620) );
  nnd2s1 U6778 ( .DIN1(reg_out_B[27]), .DIN2(n5762), .Q(n5761) );
  nnd2s1 U6779 ( .DIN1(n5763), .DIN2(n38), .Q(n5762) );
  nnd2s1 U6780 ( .DIN1(n407), .DIN2(n5764), .Q(n5760) );
  or2s1 U6781 ( .DIN1(n5624), .DIN2(n706), .Q(n5758) );
  nnd2s1 U6782 ( .DIN1(n5765), .DIN2(n5766), .Q(n5624) );
  nnd2s1 U6783 ( .DIN1(n5767), .DIN2(n5768), .Q(n5766) );
  nnd2s1 U6784 ( .DIN1(n5769), .DIN2(n5468), .Q(n5749) );
  nnd2s1 U6785 ( .DIN1(n12), .DIN2(n768), .Q(n5748) );
  nnd2s1 U6786 ( .DIN1(reg_out_B[28]), .DIN2(n5770), .Q(n5746) );
  nnd2s1 U6787 ( .DIN1(n723), .DIN2(n5771), .Q(n5770) );
  nnd2s1 U6788 ( .DIN1(n775), .DIN2(n434), .Q(n5771) );
  nnd3s1 U6789 ( .DIN1(n5772), .DIN2(n5773), .DIN3(n769), .Q(n5745) );
  nnd2s1 U6790 ( .DIN1(n5649), .DIN2(n5774), .Q(n5773) );
  nnd2s1 U6791 ( .DIN1(n5769), .DIN2(n5478), .Q(n5774) );
  nnd2s1 U6792 ( .DIN1(n5775), .DIN2(n5776), .Q(n5744) );
  nnd3s1 U6793 ( .DIN1(n5777), .DIN2(n5778), .DIN3(n204), .Q(n5776) );
  nnd2s1 U6794 ( .DIN1(n5779), .DIN2(n801), .Q(n5778) );
  nnd2s1 U6795 ( .DIN1(n5780), .DIN2(n5781), .Q(n5779) );
  nnd2s1 U6796 ( .DIN1(n742), .DIN2(n5782), .Q(n5781) );
  nnd2s1 U6797 ( .DIN1(n5783), .DIN2(n205), .Q(n5780) );
  nnd4s1 U6798 ( .DIN1(n5784), .DIN2(n5785), .DIN3(n5786), .DIN4(n5787), 
        .Q(n5783) );
  nnd2s1 U6799 ( .DIN1(n5788), .DIN2(n438), .Q(n5777) );
  nnd2s1 U6800 ( .DIN1(n5789), .DIN2(n5790), .Q(n5788) );
  nnd2s1 U6801 ( .DIN1(n32), .DIN2(n5791), .Q(n5790) );
  nnd2s1 U6802 ( .DIN1(n5792), .DIN2(n205), .Q(n5789) );
  nnd2s1 U6803 ( .DIN1(n5342), .DIN2(n5793), .Q(n5775) );
  nnd2s1 U6804 ( .DIN1(n387), .DIN2(n5794), .Q(n5793) );
  nor2s1 U6805 ( .DIN1(n5288), .DIN2(n5795), .Q(n5682) );
  or4s1 U6806 ( .DIN1(n5796), .DIN2(n5797), .DIN3(n5798), .DIN4(n5799), 
        .Q(\EXinst/n1459 ) );
  nnd4s1 U6807 ( .DIN1(n5800), .DIN2(n5801), .DIN3(n5802), .DIN4(n5803), 
        .Q(n5799) );
  nnd2s1 U6808 ( .DIN1(n5804), .DIN2(n5805), .Q(n5803) );
  nnd2s1 U6809 ( .DIN1(n5573), .DIN2(n5806), .Q(n5805) );
  nnd3s1 U6810 ( .DIN1(n5807), .DIN2(n5553), .DIN3(n555), .Q(n5806) );
  nor2s1 U6811 ( .DIN1(n5808), .DIN2(n5809), .Q(n5573) );
  nnd2s1 U6812 ( .DIN1(n5554), .DIN2(n5810), .Q(n5804) );
  nnd2s1 U6813 ( .DIN1(n5551), .DIN2(n5811), .Q(n5810) );
  nnd2s1 U6814 ( .DIN1(n5812), .DIN2(n5813), .Q(n5802) );
  nnd4s1 U6815 ( .DIN1(n5814), .DIN2(n5815), .DIN3(n5816), .DIN4(n5817), 
        .Q(n5813) );
  nor2s1 U6816 ( .DIN1(n5818), .DIN2(n805), .Q(n5817) );
  and2s1 U6817 ( .DIN1(n5302), .DIN2(n554), .Q(n5818) );
  nnd4s1 U6818 ( .DIN1(n5819), .DIN2(n5820), .DIN3(n5821), .DIN4(n5822), 
        .Q(n5302) );
  nnd2s1 U6819 ( .DIN1(n545), .DIN2(n5823), .Q(n5816) );
  nnd2s1 U6820 ( .DIN1(n5824), .DIN2(n5825), .Q(n5815) );
  nnd2s1 U6821 ( .DIN1(n726), .DIN2(n5827), .Q(n5814) );
  nnd2s1 U6822 ( .DIN1(n5547), .DIN2(n5828), .Q(n5812) );
  nnd2s1 U6823 ( .DIN1(n5301), .DIN2(n5829), .Q(n5828) );
  nnd2s1 U6824 ( .DIN1(n5323), .DIN2(n5830), .Q(n5801) );
  nnd2s1 U6825 ( .DIN1(n782), .DIN2(n5831), .Q(n5800) );
  nnd4s1 U6826 ( .DIN1(n5832), .DIN2(n5833), .DIN3(n5834), .DIN4(n5835), 
        .Q(n5831) );
  and4s1 U6827 ( .DIN1(n5836), .DIN2(n5837), .DIN3(n5838), .DIN4(n5839), 
        .Q(n5835) );
  nnd2s1 U6828 ( .DIN1(n5840), .DIN2(n5841), .Q(n5839) );
  nnd3s1 U6829 ( .DIN1(n5842), .DIN2(n749), .DIN3(n5843), .Q(n5840) );
  nnd2s1 U6830 ( .DIN1(n705), .DIN2(n5767), .Q(n5843) );
  nnd2s1 U6831 ( .DIN1(n654), .DIN2(n5763), .Q(n5842) );
  hi1s1 U6832 ( .DIN(n5764), .Q(n5763) );
  nnd2s1 U6833 ( .DIN1(n5844), .DIN2(n5845), .Q(n5838) );
  nnd2s1 U6834 ( .DIN1(n5846), .DIN2(n5847), .Q(n5845) );
  nnd2s1 U6835 ( .DIN1(n653), .DIN2(n5764), .Q(n5847) );
  nnd2s1 U6836 ( .DIN1(n5848), .DIN2(n5849), .Q(n5764) );
  nnd2s1 U6837 ( .DIN1(reg_out_B[26]), .DIN2(n5850), .Q(n5849) );
  nnd2s1 U6838 ( .DIN1(n5851), .DIN2(n336), .Q(n5850) );
  nnd2s1 U6839 ( .DIN1(n435), .DIN2(n5852), .Q(n5848) );
  or2s1 U6840 ( .DIN1(n5767), .DIN2(n706), .Q(n5846) );
  nnd2s1 U6841 ( .DIN1(n5853), .DIN2(n5854), .Q(n5767) );
  nnd2s1 U6842 ( .DIN1(n5855), .DIN2(n5856), .Q(n5854) );
  nnd2s1 U6843 ( .DIN1(n5367), .DIN2(n5857), .Q(n5837) );
  nnd2s1 U6844 ( .DIN1(n407), .DIN2(n767), .Q(n5836) );
  nnd2s1 U6845 ( .DIN1(reg_out_B[27]), .DIN2(n5858), .Q(n5834) );
  nnd2s1 U6846 ( .DIN1(n723), .DIN2(n5859), .Q(n5858) );
  nnd2s1 U6847 ( .DIN1(n776), .DIN2(n407), .Q(n5859) );
  nnd3s1 U6848 ( .DIN1(n5860), .DIN2(n5861), .DIN3(n5336), .Q(n5833) );
  nnd2s1 U6849 ( .DIN1(n5649), .DIN2(n5862), .Q(n5861) );
  nnd3s1 U6850 ( .DIN1(n5863), .DIN2(n5478), .DIN3(n628), .Q(n5862) );
  nor2s1 U6851 ( .DIN1(n5864), .DIN2(n5865), .Q(n5649) );
  nnd2s1 U6852 ( .DIN1(reg_out_B[5]), .DIN2(n5866), .Q(n5860) );
  nnd3s1 U6853 ( .DIN1(n801), .DIN2(n204), .DIN3(n5867), .Q(n5866) );
  nnd2s1 U6854 ( .DIN1(n5868), .DIN2(n5869), .Q(n5832) );
  nnd4s1 U6855 ( .DIN1(n5870), .DIN2(n5871), .DIN3(n5872), .DIN4(n5873), 
        .Q(n5869) );
  nnd2s1 U6856 ( .DIN1(n547), .DIN2(n5360), .Q(n5873) );
  nor2s1 U6857 ( .DIN1(n55), .DIN2(n5874), .Q(n5872) );
  and2s1 U6858 ( .DIN1(n5875), .DIN2(n720), .Q(n5874) );
  nnd2s1 U6859 ( .DIN1(n622), .DIN2(n5361), .Q(n5871) );
  nnd2s1 U6860 ( .DIN1(n630), .DIN2(n5358), .Q(n5870) );
  nnd4s1 U6861 ( .DIN1(n5877), .DIN2(n5878), .DIN3(n5879), .DIN4(n5880), 
        .Q(n5358) );
  nnd2s1 U6862 ( .DIN1(n5342), .DIN2(n5881), .Q(n5868) );
  nnd2s1 U6863 ( .DIN1(n387), .DIN2(n5882), .Q(n5881) );
  nnd3s1 U6864 ( .DIN1(n5883), .DIN2(n5884), .DIN3(n5885), .Q(n5798) );
  nnd2s1 U6865 ( .DIN1(n727), .DIN2(\DM_addr[27] ), .Q(n5885) );
  nnd2s1 U6866 ( .DIN1(n407), .DIN2(n5886), .Q(n5884) );
  or3s1 U6867 ( .DIN1(n405), .DIN2(n5887), .DIN3(n5888), .Q(n5886) );
  nnd4s1 U6868 ( .DIN1(n5889), .DIN2(n5890), .DIN3(n5891), .DIN4(n5892), 
        .Q(n5888) );
  nnd2s1 U6869 ( .DIN1(n548), .DIN2(n5712), .Q(n5892) );
  nnd2s1 U6870 ( .DIN1(n791), .DIN2(n5711), .Q(n5891) );
  nnd2s1 U6871 ( .DIN1(n5405), .DIN2(n95), .Q(n5890) );
  nnd2s1 U6872 ( .DIN1(n5665), .DIN2(n9464), .Q(n5889) );
  nor2s1 U6873 ( .DIN1(n5290), .DIN2(n5893), .Q(n5887) );
  nnd2s1 U6874 ( .DIN1(n5894), .DIN2(n38), .Q(n5883) );
  nnd4s1 U6875 ( .DIN1(n5895), .DIN2(n5896), .DIN3(n5897), .DIN4(n5898), 
        .Q(n5894) );
  nnd2s1 U6876 ( .DIN1(n791), .DIN2(n5712), .Q(n5898) );
  nnd2s1 U6877 ( .DIN1(n549), .DIN2(n5711), .Q(n5897) );
  hi1s1 U6878 ( .DIN(n5712), .Q(n5711) );
  nnd2s1 U6879 ( .DIN1(n5899), .DIN2(n5900), .Q(n5712) );
  nnd2s1 U6880 ( .DIN1(n6), .DIN2(n5901), .Q(n5900) );
  nnd2s1 U6881 ( .DIN1(n5902), .DIN2(n5426), .Q(n5901) );
  nnd2s1 U6882 ( .DIN1(n633), .DIN2(n5903), .Q(n5899) );
  nnd2s1 U6883 ( .DIN1(n385), .DIN2(n5893), .Q(n5896) );
  xor2s1 U6884 ( .DIN1(n5706), .DIN2(n5707), .Q(n5893) );
  xor2s1 U6885 ( .DIN1(n95), .DIN2(n745), .Q(n5707) );
  nnd2s1 U6886 ( .DIN1(n5904), .DIN2(n5905), .Q(n5706) );
  nnd2s1 U6887 ( .DIN1(n435), .DIN2(n5906), .Q(n5905) );
  nnd2s1 U6888 ( .DIN1(n5907), .DIN2(n5908), .Q(n5906) );
  or2s1 U6889 ( .DIN1(n5908), .DIN2(n5907), .Q(n5904) );
  nnd2s1 U6890 ( .DIN1(n5665), .DIN2(n95), .Q(n5895) );
  nor2s1 U6891 ( .DIN1(n9464), .DIN2(n5427), .Q(n5797) );
  nor2s1 U6892 ( .DIN1(n9480), .DIN2(n5428), .Q(n5796) );
  or4s1 U6893 ( .DIN1(n5909), .DIN2(n5910), .DIN3(n5911), .DIN4(n5912), 
        .Q(\EXinst/n1458 ) );
  nnd4s1 U6894 ( .DIN1(n5913), .DIN2(n5914), .DIN3(n5915), .DIN4(n5916), 
        .Q(n5912) );
  nor2s1 U6895 ( .DIN1(n5917), .DIN2(n5918), .Q(n5916) );
  nor2s1 U6896 ( .DIN1(n9465), .DIN2(n5427), .Q(n5918) );
  nor2s1 U6897 ( .DIN1(n9481), .DIN2(n5428), .Q(n5917) );
  nnd2s1 U6898 ( .DIN1(n5394), .DIN2(\DM_addr[26] ), .Q(n5915) );
  nnd2s1 U6899 ( .DIN1(n6), .DIN2(n5919), .Q(n5914) );
  nnd4s1 U6900 ( .DIN1(n5920), .DIN2(n5921), .DIN3(n5922), .DIN4(n5923), 
        .Q(n5919) );
  nor2s1 U6901 ( .DIN1(n404), .DIN2(n5924), .Q(n5923) );
  nor2s1 U6902 ( .DIN1(n5290), .DIN2(n5925), .Q(n5924) );
  nnd2s1 U6903 ( .DIN1(n5405), .DIN2(n103), .Q(n5922) );
  nnd2s1 U6904 ( .DIN1(n548), .DIN2(n5903), .Q(n5921) );
  nnd2s1 U6905 ( .DIN1(n791), .DIN2(n5902), .Q(n5920) );
  nnd2s1 U6906 ( .DIN1(n5926), .DIN2(n336), .Q(n5913) );
  nnd3s1 U6907 ( .DIN1(n5927), .DIN2(n5928), .DIN3(n5929), .Q(n5926) );
  nnd2s1 U6908 ( .DIN1(n385), .DIN2(n5925), .Q(n5929) );
  xor2s1 U6909 ( .DIN1(n5907), .DIN2(n5908), .Q(n5925) );
  xnr2s1 U6910 ( .DIN1(n9465), .DIN2(n787), .Q(n5908) );
  and2s1 U6911 ( .DIN1(n5930), .DIN2(n5931), .Q(n5907) );
  nnd2s1 U6912 ( .DIN1(n408), .DIN2(n5932), .Q(n5931) );
  or2s1 U6913 ( .DIN1(n5933), .DIN2(n5934), .Q(n5932) );
  nnd2s1 U6914 ( .DIN1(n5934), .DIN2(n5933), .Q(n5930) );
  nnd2s1 U6915 ( .DIN1(n791), .DIN2(n5903), .Q(n5928) );
  nnd2s1 U6916 ( .DIN1(n549), .DIN2(n5902), .Q(n5927) );
  hi1s1 U6917 ( .DIN(n5903), .Q(n5902) );
  nnd2s1 U6918 ( .DIN1(n5935), .DIN2(n5936), .Q(n5903) );
  nnd2s1 U6919 ( .DIN1(n408), .DIN2(n5937), .Q(n5936) );
  nnd2s1 U6920 ( .DIN1(n5938), .DIN2(n5426), .Q(n5937) );
  nnd2s1 U6921 ( .DIN1(n5423), .DIN2(n5939), .Q(n5935) );
  nnd3s1 U6922 ( .DIN1(n5940), .DIN2(n5941), .DIN3(n5942), .Q(n5911) );
  nnd2s1 U6923 ( .DIN1(n5323), .DIN2(n5943), .Q(n5942) );
  nor2s1 U6924 ( .DIN1(n5558), .DIN2(n803), .Q(n5323) );
  nnd3s1 U6925 ( .DIN1(n5944), .DIN2(n5945), .DIN3(n5738), .Q(n5941) );
  and4s1 U6926 ( .DIN1(n5946), .DIN2(n5947), .DIN3(n5948), .DIN4(n5553), 
        .Q(n5738) );
  nnd2s1 U6927 ( .DIN1(n5949), .DIN2(n5556), .Q(n5948) );
  nnd2s1 U6928 ( .DIN1(n735), .DIN2(n4831), .Q(n5947) );
  nnd3s1 U6929 ( .DIN1(n5741), .DIN2(n4831), .DIN3(n5950), .Q(n5945) );
  nnd2s1 U6930 ( .DIN1(n5951), .DIN2(n5739), .Q(n5944) );
  and3s1 U6931 ( .DIN1(n739), .DIN2(n5556), .DIN3(n9486), .Q(n5739) );
  nnd2s1 U6932 ( .DIN1(n5952), .DIN2(n5953), .Q(n5940) );
  nnd4s1 U6933 ( .DIN1(n740), .DIN2(n5954), .DIN3(n5955), .DIN4(n5956), 
        .Q(n5953) );
  nnd2s1 U6934 ( .DIN1(n726), .DIN2(n5535), .Q(n5956) );
  nor2s1 U6935 ( .DIN1(n5957), .DIN2(n5958), .Q(n5955) );
  and2s1 U6936 ( .DIN1(n5959), .DIN2(n5824), .Q(n5958) );
  and2s1 U6937 ( .DIN1(n5540), .DIN2(n555), .Q(n5957) );
  nnd3s1 U6938 ( .DIN1(n5960), .DIN2(n5961), .DIN3(n5962), .Q(n5540) );
  nnd3s1 U6939 ( .DIN1(n5963), .DIN2(n5964), .DIN3(n707), .Q(n5961) );
  nnd2s1 U6940 ( .DIN1(n9489), .DIN2(n30), .Q(n5964) );
  nnd2s1 U6941 ( .DIN1(n439), .DIN2(n68), .Q(n5963) );
  nnd2s1 U6942 ( .DIN1(n544), .DIN2(n5536), .Q(n5954) );
  nnd2s1 U6943 ( .DIN1(n5547), .DIN2(n5965), .Q(n5952) );
  nnd2s1 U6944 ( .DIN1(n5301), .DIN2(n5966), .Q(n5965) );
  and2s1 U6945 ( .DIN1(n782), .DIN2(n5967), .Q(n5910) );
  nnd4s1 U6946 ( .DIN1(n5968), .DIN2(n5969), .DIN3(n5970), .DIN4(n5971), 
        .Q(n5967) );
  and4s1 U6947 ( .DIN1(n5972), .DIN2(n5973), .DIN3(n5974), .DIN4(n5975), 
        .Q(n5971) );
  nnd2s1 U6948 ( .DIN1(n5976), .DIN2(n5977), .Q(n5975) );
  nnd3s1 U6949 ( .DIN1(n5978), .DIN2(n5372), .DIN3(n5979), .Q(n5976) );
  nnd2s1 U6950 ( .DIN1(n620), .DIN2(n5856), .Q(n5979) );
  nnd2s1 U6951 ( .DIN1(n656), .DIN2(n5851), .Q(n5978) );
  hi1s1 U6952 ( .DIN(n5852), .Q(n5851) );
  nnd2s1 U6953 ( .DIN1(n5980), .DIN2(n5981), .Q(n5974) );
  nnd2s1 U6954 ( .DIN1(n5982), .DIN2(n5983), .Q(n5981) );
  nnd2s1 U6955 ( .DIN1(n655), .DIN2(n5852), .Q(n5983) );
  nnd2s1 U6956 ( .DIN1(n5984), .DIN2(n5985), .Q(n5852) );
  nnd2s1 U6957 ( .DIN1(reg_out_B[25]), .DIN2(n5986), .Q(n5985) );
  nnd2s1 U6958 ( .DIN1(n5987), .DIN2(n83), .Q(n5986) );
  nnd2s1 U6959 ( .DIN1(n408), .DIN2(n5988), .Q(n5984) );
  or2s1 U6960 ( .DIN1(n5856), .DIN2(n706), .Q(n5982) );
  nnd2s1 U6961 ( .DIN1(n5989), .DIN2(n5990), .Q(n5856) );
  nnd2s1 U6962 ( .DIN1(n5991), .DIN2(n5992), .Q(n5990) );
  nnd2s1 U6963 ( .DIN1(n5367), .DIN2(n5993), .Q(n5973) );
  nor2s1 U6964 ( .DIN1(n5994), .DIN2(n438), .Q(n5367) );
  nnd2s1 U6965 ( .DIN1(n435), .DIN2(n768), .Q(n5972) );
  nnd2s1 U6966 ( .DIN1(reg_out_B[26]), .DIN2(n5995), .Q(n5970) );
  nnd2s1 U6967 ( .DIN1(n723), .DIN2(n5996), .Q(n5995) );
  nnd2s1 U6968 ( .DIN1(n775), .DIN2(n435), .Q(n5996) );
  nnd3s1 U6969 ( .DIN1(n5997), .DIN2(n5998), .DIN3(n769), .Q(n5969) );
  nnd2s1 U6970 ( .DIN1(n5475), .DIN2(n5999), .Q(n5998) );
  nnd3s1 U6971 ( .DIN1(n5478), .DIN2(n337), .DIN3(n6000), .Q(n5999) );
  nnd2s1 U6972 ( .DIN1(n6001), .DIN2(n6002), .Q(n5997) );
  nnd2s1 U6973 ( .DIN1(n5366), .DIN2(n714), .Q(n6002) );
  hi1s1 U6974 ( .DIN(n5772), .Q(n6001) );
  nnd2s1 U6975 ( .DIN1(reg_out_B[5]), .DIN2(n6003), .Q(n5772) );
  nnd2s1 U6976 ( .DIN1(n5480), .DIN2(n337), .Q(n6003) );
  nnd2s1 U6977 ( .DIN1(n6004), .DIN2(n6005), .Q(n5968) );
  nnd4s1 U6978 ( .DIN1(n6006), .DIN2(n807), .DIN3(n6007), .DIN4(n6008), 
        .Q(n6005) );
  nor2s1 U6979 ( .DIN1(n6009), .DIN2(n6010), .Q(n6008) );
  and2s1 U6980 ( .DIN1(n5500), .DIN2(n623), .Q(n6010) );
  and2s1 U6981 ( .DIN1(n5499), .DIN2(n547), .Q(n6009) );
  nnd2s1 U6982 ( .DIN1(n720), .DIN2(n6011), .Q(n6007) );
  nnd2s1 U6983 ( .DIN1(n629), .DIN2(n5488), .Q(n6006) );
  nnd3s1 U6984 ( .DIN1(n6012), .DIN2(n6013), .DIN3(n6014), .Q(n5488) );
  nnd3s1 U6985 ( .DIN1(n6015), .DIN2(n6016), .DIN3(reg_out_B[1]), .Q(n6013) );
  nnd2s1 U6986 ( .DIN1(n30), .DIN2(n1), .Q(n6016) );
  nnd2s1 U6987 ( .DIN1(n399), .DIN2(n68), .Q(n6015) );
  nnd2s1 U6988 ( .DIN1(n5342), .DIN2(n6017), .Q(n6004) );
  nnd2s1 U6989 ( .DIN1(n387), .DIN2(n6018), .Q(n6017) );
  nor2s1 U6990 ( .DIN1(n5288), .DIN2(n6019), .Q(n5909) );
  or4s1 U6991 ( .DIN1(n6020), .DIN2(n6021), .DIN3(n6022), .DIN4(n6023), 
        .Q(\EXinst/n1457 ) );
  nnd4s1 U6992 ( .DIN1(n6024), .DIN2(n6025), .DIN3(n6026), .DIN4(n6027), 
        .Q(n6023) );
  nnd2s1 U6993 ( .DIN1(n6028), .DIN2(n6029), .Q(n6027) );
  nnd2s1 U6994 ( .DIN1(n6030), .DIN2(n6031), .Q(n6029) );
  nnd2s1 U6995 ( .DIN1(n6032), .DIN2(n5553), .Q(n6031) );
  nnd2s1 U6996 ( .DIN1(n5554), .DIN2(n6033), .Q(n6028) );
  nnd2s1 U6997 ( .DIN1(n5551), .DIN2(n6034), .Q(n6033) );
  and2s1 U6998 ( .DIN1(n5322), .DIN2(n736), .Q(n5551) );
  nnd2s1 U6999 ( .DIN1(n6035), .DIN2(n6036), .Q(n5554) );
  nnd2s1 U7000 ( .DIN1(n6037), .DIN2(n6038), .Q(n6026) );
  nnd4s1 U7001 ( .DIN1(n56), .DIN2(n6039), .DIN3(n6040), .DIN4(n6041), 
        .Q(n6038) );
  nnd2s1 U7002 ( .DIN1(n726), .DIN2(n5586), .Q(n6041) );
  nor2s1 U7003 ( .DIN1(n6042), .DIN2(n6043), .Q(n6040) );
  and2s1 U7004 ( .DIN1(n6044), .DIN2(n5824), .Q(n6043) );
  and2s1 U7005 ( .DIN1(n5591), .DIN2(n554), .Q(n6042) );
  nnd3s1 U7006 ( .DIN1(n6045), .DIN2(n6046), .DIN3(n6047), .Q(n5591) );
  nnd3s1 U7007 ( .DIN1(n6048), .DIN2(n6049), .DIN3(n707), .Q(n6046) );
  nnd2s1 U7008 ( .DIN1(n9489), .DIN2(n68), .Q(n6049) );
  nnd2s1 U7009 ( .DIN1(n440), .DIN2(n67), .Q(n6048) );
  nnd2s1 U7010 ( .DIN1(n545), .DIN2(n5587), .Q(n6039) );
  nnd2s1 U7011 ( .DIN1(n5547), .DIN2(n6050), .Q(n6037) );
  nnd2s1 U7012 ( .DIN1(n5301), .DIN2(n6051), .Q(n6050) );
  or2s1 U7013 ( .DIN1(n6052), .DIN2(n5558), .Q(n6025) );
  nnd2s1 U7014 ( .DIN1(n782), .DIN2(n6053), .Q(n6024) );
  nnd4s1 U7015 ( .DIN1(n6054), .DIN2(n6055), .DIN3(n6056), .DIN4(n6057), 
        .Q(n6053) );
  and4s1 U7016 ( .DIN1(n6058), .DIN2(n6059), .DIN3(n6060), .DIN4(n6061), 
        .Q(n6057) );
  nnd2s1 U7017 ( .DIN1(n6062), .DIN2(n6063), .Q(n6061) );
  nnd3s1 U7018 ( .DIN1(n6064), .DIN2(n749), .DIN3(n6065), .Q(n6062) );
  nnd2s1 U7019 ( .DIN1(n705), .DIN2(n5991), .Q(n6065) );
  nnd2s1 U7020 ( .DIN1(n654), .DIN2(n5987), .Q(n6064) );
  hi1s1 U7021 ( .DIN(n5988), .Q(n5987) );
  nnd2s1 U7022 ( .DIN1(n6066), .DIN2(n6067), .Q(n6060) );
  nnd2s1 U7023 ( .DIN1(n6068), .DIN2(n6069), .Q(n6067) );
  nnd2s1 U7024 ( .DIN1(n653), .DIN2(n5988), .Q(n6069) );
  nnd2s1 U7025 ( .DIN1(n6070), .DIN2(n6071), .Q(n5988) );
  nnd2s1 U7026 ( .DIN1(reg_out_B[24]), .DIN2(n6072), .Q(n6071) );
  nnd2s1 U7027 ( .DIN1(n6073), .DIN2(n30), .Q(n6072) );
  nnd2s1 U7028 ( .DIN1(n409), .DIN2(n6074), .Q(n6070) );
  or2s1 U7029 ( .DIN1(n5991), .DIN2(n5375), .Q(n6068) );
  nnd2s1 U7030 ( .DIN1(n6075), .DIN2(n6076), .Q(n5991) );
  nnd2s1 U7031 ( .DIN1(n6077), .DIN2(n6078), .Q(n6076) );
  nnd2s1 U7032 ( .DIN1(n6079), .DIN2(n5468), .Q(n6059) );
  nnd2s1 U7033 ( .DIN1(n408), .DIN2(n767), .Q(n6058) );
  nnd2s1 U7034 ( .DIN1(reg_out_B[25]), .DIN2(n6080), .Q(n6056) );
  nnd2s1 U7035 ( .DIN1(n723), .DIN2(n6081), .Q(n6080) );
  nnd2s1 U7036 ( .DIN1(n776), .DIN2(n408), .Q(n6081) );
  nnd3s1 U7037 ( .DIN1(n6082), .DIN2(n6083), .DIN3(n5336), .Q(n6055) );
  nnd2s1 U7038 ( .DIN1(n5475), .DIN2(n6084), .Q(n6083) );
  nnd2s1 U7039 ( .DIN1(n6085), .DIN2(n5478), .Q(n6084) );
  nnd2s1 U7040 ( .DIN1(reg_out_B[5]), .DIN2(n6086), .Q(n6082) );
  nnd3s1 U7041 ( .DIN1(n337), .DIN2(n808), .DIN3(n6087), .Q(n6086) );
  nnd2s1 U7042 ( .DIN1(n6088), .DIN2(n6089), .Q(n6054) );
  nnd4s1 U7043 ( .DIN1(n6090), .DIN2(n807), .DIN3(n6091), .DIN4(n6092), 
        .Q(n6089) );
  nor2s1 U7044 ( .DIN1(n6093), .DIN2(n6094), .Q(n6092) );
  and2s1 U7045 ( .DIN1(n5644), .DIN2(n622), .Q(n6094) );
  and2s1 U7046 ( .DIN1(n5643), .DIN2(n546), .Q(n6093) );
  nnd2s1 U7047 ( .DIN1(n720), .DIN2(n6095), .Q(n6091) );
  nnd2s1 U7048 ( .DIN1(n630), .DIN2(n5634), .Q(n6090) );
  nnd3s1 U7049 ( .DIN1(n6096), .DIN2(n6097), .DIN3(n6098), .Q(n5634) );
  nnd3s1 U7050 ( .DIN1(n6099), .DIN2(n6100), .DIN3(reg_out_B[1]), .Q(n6097) );
  nnd2s1 U7051 ( .DIN1(n68), .DIN2(n1), .Q(n6100) );
  nnd2s1 U7052 ( .DIN1(n399), .DIN2(n67), .Q(n6099) );
  nnd2s1 U7053 ( .DIN1(n5342), .DIN2(n6101), .Q(n6088) );
  nnd2s1 U7054 ( .DIN1(n387), .DIN2(n6102), .Q(n6101) );
  nnd3s1 U7055 ( .DIN1(n6103), .DIN2(n6104), .DIN3(n6105), .Q(n6022) );
  nnd2s1 U7056 ( .DIN1(n727), .DIN2(\DM_addr[25] ), .Q(n6105) );
  nnd2s1 U7057 ( .DIN1(n408), .DIN2(n6106), .Q(n6104) );
  or3s1 U7058 ( .DIN1(n403), .DIN2(n6107), .DIN3(n6108), .Q(n6106) );
  nnd4s1 U7059 ( .DIN1(n6109), .DIN2(n6110), .DIN3(n6111), .DIN4(n6112), 
        .Q(n6108) );
  nnd2s1 U7060 ( .DIN1(n548), .DIN2(n5939), .Q(n6112) );
  nnd2s1 U7061 ( .DIN1(n791), .DIN2(n5938), .Q(n6111) );
  nnd2s1 U7062 ( .DIN1(n5405), .DIN2(n15), .Q(n6110) );
  nnd2s1 U7063 ( .DIN1(n5665), .DIN2(n9466), .Q(n6109) );
  nor2s1 U7064 ( .DIN1(n5290), .DIN2(n6113), .Q(n6107) );
  nnd2s1 U7065 ( .DIN1(n6114), .DIN2(n83), .Q(n6103) );
  nnd4s1 U7066 ( .DIN1(n6115), .DIN2(n6116), .DIN3(n6117), .DIN4(n6118), 
        .Q(n6114) );
  nnd2s1 U7067 ( .DIN1(n791), .DIN2(n5939), .Q(n6118) );
  nnd2s1 U7068 ( .DIN1(n549), .DIN2(n5938), .Q(n6117) );
  hi1s1 U7069 ( .DIN(n5939), .Q(n5938) );
  nnd2s1 U7070 ( .DIN1(n6119), .DIN2(n6120), .Q(n5939) );
  nnd2s1 U7071 ( .DIN1(n409), .DIN2(n6121), .Q(n6120) );
  nnd2s1 U7072 ( .DIN1(n6122), .DIN2(n5426), .Q(n6121) );
  nnd2s1 U7073 ( .DIN1(n633), .DIN2(n6123), .Q(n6119) );
  nnd2s1 U7074 ( .DIN1(n385), .DIN2(n6113), .Q(n6116) );
  xor2s1 U7075 ( .DIN1(n5933), .DIN2(n5934), .Q(n6113) );
  xor2s1 U7076 ( .DIN1(n15), .DIN2(n5413), .Q(n5934) );
  nnd2s1 U7077 ( .DIN1(n6124), .DIN2(n6125), .Q(n5933) );
  nnd2s1 U7078 ( .DIN1(n409), .DIN2(n6126), .Q(n6125) );
  nnd2s1 U7079 ( .DIN1(n6127), .DIN2(n6128), .Q(n6126) );
  or2s1 U7080 ( .DIN1(n6128), .DIN2(n6127), .Q(n6124) );
  nnd2s1 U7081 ( .DIN1(n5665), .DIN2(n15), .Q(n6115) );
  nor2s1 U7082 ( .DIN1(n9466), .DIN2(n5427), .Q(n6021) );
  nor2s1 U7083 ( .DIN1(n9482), .DIN2(n5428), .Q(n6020) );
  or4s1 U7084 ( .DIN1(n6129), .DIN2(n6130), .DIN3(n6131), .DIN4(n6132), 
        .Q(\EXinst/n1456 ) );
  nnd4s1 U7085 ( .DIN1(n6133), .DIN2(n6134), .DIN3(n6135), .DIN4(n6136), 
        .Q(n6132) );
  nor2s1 U7086 ( .DIN1(n6137), .DIN2(n6138), .Q(n6136) );
  nor2s1 U7087 ( .DIN1(n9467), .DIN2(n5427), .Q(n6138) );
  nor2s1 U7088 ( .DIN1(n9483), .DIN2(n5428), .Q(n6137) );
  nnd2s1 U7089 ( .DIN1(n5394), .DIN2(\DM_addr[24] ), .Q(n6135) );
  nnd2s1 U7090 ( .DIN1(n409), .DIN2(n6139), .Q(n6134) );
  nnd4s1 U7091 ( .DIN1(n6140), .DIN2(n6141), .DIN3(n6142), .DIN4(n6143), 
        .Q(n6139) );
  nor2s1 U7092 ( .DIN1(n403), .DIN2(n6144), .Q(n6143) );
  nor2s1 U7093 ( .DIN1(n5290), .DIN2(n6145), .Q(n6144) );
  nnd2s1 U7094 ( .DIN1(n5405), .DIN2(n120), .Q(n6142) );
  nnd2s1 U7095 ( .DIN1(n548), .DIN2(n6123), .Q(n6141) );
  nnd2s1 U7096 ( .DIN1(n791), .DIN2(n6122), .Q(n6140) );
  nnd2s1 U7097 ( .DIN1(n6146), .DIN2(n30), .Q(n6133) );
  nnd3s1 U7098 ( .DIN1(n6147), .DIN2(n6148), .DIN3(n6149), .Q(n6146) );
  nnd2s1 U7099 ( .DIN1(n385), .DIN2(n6145), .Q(n6149) );
  xor2s1 U7100 ( .DIN1(n6127), .DIN2(n6128), .Q(n6145) );
  xnr2s1 U7101 ( .DIN1(n9467), .DIN2(n786), .Q(n6128) );
  and2s1 U7102 ( .DIN1(n6150), .DIN2(n6151), .Q(n6127) );
  nnd2s1 U7103 ( .DIN1(n410), .DIN2(n6152), .Q(n6151) );
  or2s1 U7104 ( .DIN1(n6153), .DIN2(n6154), .Q(n6152) );
  nnd2s1 U7105 ( .DIN1(n6154), .DIN2(n6153), .Q(n6150) );
  nnd2s1 U7106 ( .DIN1(n5406), .DIN2(n6123), .Q(n6148) );
  nnd2s1 U7107 ( .DIN1(n549), .DIN2(n6122), .Q(n6147) );
  hi1s1 U7108 ( .DIN(n6123), .Q(n6122) );
  nnd2s1 U7109 ( .DIN1(n6155), .DIN2(n6156), .Q(n6123) );
  nnd2s1 U7110 ( .DIN1(n410), .DIN2(n6157), .Q(n6156) );
  nnd2s1 U7111 ( .DIN1(n6158), .DIN2(n5426), .Q(n6157) );
  nnd2s1 U7112 ( .DIN1(n5423), .DIN2(n6159), .Q(n6155) );
  nnd3s1 U7113 ( .DIN1(n6160), .DIN2(n6161), .DIN3(n6162), .Q(n6131) );
  or2s1 U7114 ( .DIN1(n6163), .DIN2(n5288), .Q(n6162) );
  nnd2s1 U7115 ( .DIN1(n6164), .DIN2(n6165), .Q(n6161) );
  nnd2s1 U7116 ( .DIN1(n6030), .DIN2(n6166), .Q(n6165) );
  nnd2s1 U7117 ( .DIN1(n6167), .DIN2(n5553), .Q(n6166) );
  hi1s1 U7118 ( .DIN(n6168), .Q(n6164) );
  nnd2s1 U7119 ( .DIN1(n6169), .DIN2(n6170), .Q(n6160) );
  nnd4s1 U7120 ( .DIN1(n739), .DIN2(n6171), .DIN3(n6172), .DIN4(n6173), 
        .Q(n6170) );
  nnd2s1 U7121 ( .DIN1(n726), .DIN2(n5723), .Q(n6173) );
  nor2s1 U7122 ( .DIN1(n6174), .DIN2(n6175), .Q(n6172) );
  and2s1 U7123 ( .DIN1(n6176), .DIN2(n5824), .Q(n6175) );
  and2s1 U7124 ( .DIN1(n5728), .DIN2(n555), .Q(n6174) );
  nnd3s1 U7125 ( .DIN1(n6177), .DIN2(n6178), .DIN3(n6179), .Q(n5728) );
  nnd3s1 U7126 ( .DIN1(n6180), .DIN2(n6181), .DIN3(n707), .Q(n6178) );
  nnd2s1 U7127 ( .DIN1(n9489), .DIN2(n67), .Q(n6181) );
  nnd2s1 U7128 ( .DIN1(n439), .DIN2(n78), .Q(n6180) );
  nnd2s1 U7129 ( .DIN1(n544), .DIN2(n5724), .Q(n6171) );
  nnd2s1 U7130 ( .DIN1(n5547), .DIN2(n6182), .Q(n6169) );
  nnd2s1 U7131 ( .DIN1(n5301), .DIN2(n6183), .Q(n6182) );
  and2s1 U7132 ( .DIN1(n782), .DIN2(n6184), .Q(n6130) );
  nnd4s1 U7133 ( .DIN1(n6185), .DIN2(n6186), .DIN3(n6187), .DIN4(n6188), 
        .Q(n6184) );
  and4s1 U7134 ( .DIN1(n6189), .DIN2(n6190), .DIN3(n6191), .DIN4(n6192), 
        .Q(n6188) );
  nnd2s1 U7135 ( .DIN1(n6193), .DIN2(n6194), .Q(n6192) );
  nnd3s1 U7136 ( .DIN1(n6195), .DIN2(n5372), .DIN3(n6196), .Q(n6193) );
  nnd2s1 U7137 ( .DIN1(n620), .DIN2(n6078), .Q(n6196) );
  nnd2s1 U7138 ( .DIN1(n656), .DIN2(n6073), .Q(n6195) );
  hi1s1 U7139 ( .DIN(n6074), .Q(n6073) );
  nnd2s1 U7140 ( .DIN1(n6197), .DIN2(n6198), .Q(n6191) );
  nnd2s1 U7141 ( .DIN1(n6199), .DIN2(n6200), .Q(n6198) );
  nnd2s1 U7142 ( .DIN1(n655), .DIN2(n6074), .Q(n6200) );
  nnd2s1 U7143 ( .DIN1(n6201), .DIN2(n6202), .Q(n6074) );
  nnd2s1 U7144 ( .DIN1(reg_out_B[23]), .DIN2(n6203), .Q(n6202) );
  nnd2s1 U7145 ( .DIN1(n6204), .DIN2(n68), .Q(n6203) );
  nnd2s1 U7146 ( .DIN1(n410), .DIN2(n6205), .Q(n6201) );
  or2s1 U7147 ( .DIN1(n6078), .DIN2(n706), .Q(n6199) );
  nnd2s1 U7148 ( .DIN1(n6206), .DIN2(n6207), .Q(n6078) );
  nnd2s1 U7149 ( .DIN1(n6208), .DIN2(n6209), .Q(n6207) );
  nnd2s1 U7150 ( .DIN1(n6210), .DIN2(n5468), .Q(n6190) );
  nnd2s1 U7151 ( .DIN1(n409), .DIN2(n768), .Q(n6189) );
  nnd2s1 U7152 ( .DIN1(reg_out_B[24]), .DIN2(n6211), .Q(n6187) );
  nnd2s1 U7153 ( .DIN1(n723), .DIN2(n6212), .Q(n6211) );
  nnd2s1 U7154 ( .DIN1(n775), .DIN2(n409), .Q(n6212) );
  nnd3s1 U7155 ( .DIN1(n6213), .DIN2(n6214), .DIN3(n769), .Q(n6186) );
  nnd2s1 U7156 ( .DIN1(n5475), .DIN2(n6215), .Q(n6214) );
  nnd2s1 U7157 ( .DIN1(n6210), .DIN2(n5478), .Q(n6215) );
  nor2s1 U7158 ( .DIN1(n5865), .DIN2(n6216), .Q(n5475) );
  nnd2s1 U7159 ( .DIN1(n6217), .DIN2(n6218), .Q(n6185) );
  nnd4s1 U7160 ( .DIN1(n6219), .DIN2(n807), .DIN3(n6220), .DIN4(n6221), 
        .Q(n6218) );
  nor2s1 U7161 ( .DIN1(n6222), .DIN2(n6223), .Q(n6221) );
  and2s1 U7162 ( .DIN1(n5792), .DIN2(n621), .Q(n6223) );
  and2s1 U7163 ( .DIN1(n5791), .DIN2(n547), .Q(n6222) );
  nnd2s1 U7164 ( .DIN1(n720), .DIN2(n6224), .Q(n6220) );
  nnd2s1 U7165 ( .DIN1(n629), .DIN2(n5782), .Q(n6219) );
  nnd3s1 U7166 ( .DIN1(n6225), .DIN2(n6226), .DIN3(n6227), .Q(n5782) );
  nnd3s1 U7167 ( .DIN1(n6228), .DIN2(n6229), .DIN3(reg_out_B[1]), .Q(n6226) );
  nnd2s1 U7168 ( .DIN1(n67), .DIN2(n1), .Q(n6229) );
  nnd2s1 U7169 ( .DIN1(n399), .DIN2(n78), .Q(n6228) );
  nnd2s1 U7170 ( .DIN1(n5342), .DIN2(n6230), .Q(n6217) );
  nnd2s1 U7171 ( .DIN1(n387), .DIN2(n6231), .Q(n6230) );
  nor2s1 U7172 ( .DIN1(n5558), .DIN2(n6232), .Q(n6129) );
  or4s1 U7173 ( .DIN1(n6233), .DIN2(n6234), .DIN3(n6235), .DIN4(n6236), 
        .Q(\EXinst/n1455 ) );
  nnd4s1 U7174 ( .DIN1(n6237), .DIN2(n6238), .DIN3(n6239), .DIN4(n6240), 
        .Q(n6236) );
  nnd2s1 U7175 ( .DIN1(n6241), .DIN2(n6242), .Q(n6240) );
  nnd2s1 U7176 ( .DIN1(n6030), .DIN2(n6243), .Q(n6242) );
  nnd2s1 U7177 ( .DIN1(n6244), .DIN2(n5553), .Q(n6243) );
  nnd2s1 U7178 ( .DIN1(n6168), .DIN2(n6245), .Q(n6241) );
  nnd2s1 U7179 ( .DIN1(n5317), .DIN2(n5322), .Q(n6245) );
  nnd2s1 U7180 ( .DIN1(n6246), .DIN2(n6247), .Q(n6239) );
  nnd4s1 U7181 ( .DIN1(n6248), .DIN2(n6249), .DIN3(n6250), .DIN4(n6251), 
        .Q(n6247) );
  nor2s1 U7182 ( .DIN1(n6252), .DIN2(n806), .Q(n6251) );
  nor2s1 U7183 ( .DIN1(n5316), .DIN2(n6253), .Q(n6252) );
  hi1s1 U7184 ( .DIN(n5823), .Q(n5316) );
  nnd4s1 U7185 ( .DIN1(n6254), .DIN2(n6255), .DIN3(n6256), .DIN4(n6257), 
        .Q(n5823) );
  nnd2s1 U7186 ( .DIN1(n545), .DIN2(n5827), .Q(n6250) );
  nnd2s1 U7187 ( .DIN1(n5824), .DIN2(n6258), .Q(n6249) );
  nnd2s1 U7188 ( .DIN1(n726), .DIN2(n5825), .Q(n6248) );
  nnd2s1 U7189 ( .DIN1(n5547), .DIN2(n6259), .Q(n6246) );
  nnd2s1 U7190 ( .DIN1(n6260), .DIN2(n5301), .Q(n6259) );
  nnd2s1 U7191 ( .DIN1(n5570), .DIN2(n6261), .Q(n6238) );
  nnd2s1 U7192 ( .DIN1(n782), .DIN2(n6262), .Q(n6237) );
  nnd4s1 U7193 ( .DIN1(n6263), .DIN2(n6264), .DIN3(n6265), .DIN4(n6266), 
        .Q(n6262) );
  and4s1 U7194 ( .DIN1(n6267), .DIN2(n6268), .DIN3(n6269), .DIN4(n6270), 
        .Q(n6266) );
  nnd2s1 U7195 ( .DIN1(n6271), .DIN2(n6272), .Q(n6270) );
  nnd3s1 U7196 ( .DIN1(n6273), .DIN2(n749), .DIN3(n6274), .Q(n6271) );
  nnd2s1 U7197 ( .DIN1(n705), .DIN2(n6208), .Q(n6274) );
  nnd2s1 U7198 ( .DIN1(n654), .DIN2(n6204), .Q(n6273) );
  hi1s1 U7199 ( .DIN(n6205), .Q(n6204) );
  nnd2s1 U7200 ( .DIN1(n6275), .DIN2(n6276), .Q(n6269) );
  nnd2s1 U7201 ( .DIN1(n6277), .DIN2(n6278), .Q(n6276) );
  nnd2s1 U7202 ( .DIN1(n653), .DIN2(n6205), .Q(n6278) );
  nnd2s1 U7203 ( .DIN1(n6279), .DIN2(n6280), .Q(n6205) );
  nnd2s1 U7204 ( .DIN1(reg_out_B[22]), .DIN2(n6281), .Q(n6280) );
  nnd2s1 U7205 ( .DIN1(n6282), .DIN2(n67), .Q(n6281) );
  nnd2s1 U7206 ( .DIN1(n411), .DIN2(n6283), .Q(n6279) );
  or2s1 U7207 ( .DIN1(n6208), .DIN2(n706), .Q(n6277) );
  nnd2s1 U7208 ( .DIN1(n6284), .DIN2(n6285), .Q(n6208) );
  nnd2s1 U7209 ( .DIN1(n6286), .DIN2(n6287), .Q(n6285) );
  nnd2s1 U7210 ( .DIN1(n5468), .DIN2(n6288), .Q(n6268) );
  nnd2s1 U7211 ( .DIN1(n410), .DIN2(n767), .Q(n6267) );
  nnd2s1 U7212 ( .DIN1(reg_out_B[23]), .DIN2(n6289), .Q(n6265) );
  nnd2s1 U7213 ( .DIN1(n723), .DIN2(n6290), .Q(n6289) );
  nnd2s1 U7214 ( .DIN1(n776), .DIN2(n410), .Q(n6290) );
  nnd3s1 U7215 ( .DIN1(n6291), .DIN2(n6292), .DIN3(n6293), .Q(n6264) );
  nnd4s1 U7216 ( .DIN1(n6294), .DIN2(n807), .DIN3(n6295), .DIN4(n5337), 
        .Q(n6292) );
  nnd3s1 U7217 ( .DIN1(n6296), .DIN2(n6297), .DIN3(n801), .Q(n6295) );
  nnd2s1 U7218 ( .DIN1(n6298), .DIN2(n205), .Q(n6297) );
  nnd2s1 U7219 ( .DIN1(n6299), .DIN2(n32), .Q(n6296) );
  nnd3s1 U7220 ( .DIN1(n6300), .DIN2(n6301), .DIN3(reg_out_B[5]), .Q(n6291) );
  nnd2s1 U7221 ( .DIN1(n6302), .DIN2(n6303), .Q(n6263) );
  nnd4s1 U7222 ( .DIN1(n6304), .DIN2(n6305), .DIN3(n6306), .DIN4(n6307), 
        .Q(n6303) );
  nnd2s1 U7223 ( .DIN1(n546), .DIN2(n5875), .Q(n6307) );
  nor2s1 U7224 ( .DIN1(n752), .DIN2(n6308), .Q(n6306) );
  and2s1 U7225 ( .DIN1(n6309), .DIN2(n720), .Q(n6308) );
  nnd2s1 U7226 ( .DIN1(n621), .DIN2(n5360), .Q(n6305) );
  nnd2s1 U7227 ( .DIN1(n630), .DIN2(n5361), .Q(n6304) );
  nnd4s1 U7228 ( .DIN1(n6310), .DIN2(n6311), .DIN3(n6312), .DIN4(n6313), 
        .Q(n5361) );
  nnd2s1 U7229 ( .DIN1(n5342), .DIN2(n6314), .Q(n6302) );
  nnd2s1 U7230 ( .DIN1(n6315), .DIN2(n387), .Q(n6314) );
  nnd3s1 U7231 ( .DIN1(n6316), .DIN2(n6317), .DIN3(n6318), .Q(n6235) );
  nnd2s1 U7232 ( .DIN1(n727), .DIN2(\DM_addr[23] ), .Q(n6318) );
  nnd2s1 U7233 ( .DIN1(n410), .DIN2(n6319), .Q(n6317) );
  or3s1 U7234 ( .DIN1(n404), .DIN2(n6320), .DIN3(n6321), .Q(n6319) );
  nnd4s1 U7235 ( .DIN1(n6322), .DIN2(n6323), .DIN3(n6324), .DIN4(n6325), 
        .Q(n6321) );
  nnd2s1 U7236 ( .DIN1(n548), .DIN2(n6159), .Q(n6325) );
  nnd2s1 U7237 ( .DIN1(n5406), .DIN2(n6158), .Q(n6324) );
  nnd2s1 U7238 ( .DIN1(n5405), .DIN2(n93), .Q(n6323) );
  nnd2s1 U7239 ( .DIN1(n5665), .DIN2(n9468), .Q(n6322) );
  nor2s1 U7240 ( .DIN1(n5290), .DIN2(n6326), .Q(n6320) );
  nnd2s1 U7241 ( .DIN1(n6327), .DIN2(n68), .Q(n6316) );
  nnd4s1 U7242 ( .DIN1(n6328), .DIN2(n6329), .DIN3(n6330), .DIN4(n6331), 
        .Q(n6327) );
  nnd2s1 U7243 ( .DIN1(n5406), .DIN2(n6159), .Q(n6331) );
  nnd2s1 U7244 ( .DIN1(n549), .DIN2(n6158), .Q(n6330) );
  hi1s1 U7245 ( .DIN(n6159), .Q(n6158) );
  nnd2s1 U7246 ( .DIN1(n6332), .DIN2(n6333), .Q(n6159) );
  nnd2s1 U7247 ( .DIN1(n411), .DIN2(n6334), .Q(n6333) );
  nnd2s1 U7248 ( .DIN1(n6335), .DIN2(n5426), .Q(n6334) );
  nnd2s1 U7249 ( .DIN1(n633), .DIN2(n6336), .Q(n6332) );
  nnd2s1 U7250 ( .DIN1(n385), .DIN2(n6326), .Q(n6329) );
  xor2s1 U7251 ( .DIN1(n6153), .DIN2(n6154), .Q(n6326) );
  xor2s1 U7252 ( .DIN1(n93), .DIN2(n745), .Q(n6154) );
  nnd2s1 U7253 ( .DIN1(n6337), .DIN2(n6338), .Q(n6153) );
  nnd2s1 U7254 ( .DIN1(n411), .DIN2(n6339), .Q(n6338) );
  nnd2s1 U7255 ( .DIN1(n6340), .DIN2(n6341), .Q(n6339) );
  or2s1 U7256 ( .DIN1(n6341), .DIN2(n6340), .Q(n6337) );
  nnd2s1 U7257 ( .DIN1(n5665), .DIN2(n93), .Q(n6328) );
  nor2s1 U7258 ( .DIN1(n9468), .DIN2(n5427), .Q(n6234) );
  nor2s1 U7259 ( .DIN1(n9484), .DIN2(n5428), .Q(n6233) );
  or4s1 U7260 ( .DIN1(n6342), .DIN2(n6343), .DIN3(n6344), .DIN4(n6345), 
        .Q(\EXinst/n1454 ) );
  nnd4s1 U7261 ( .DIN1(n6346), .DIN2(n6347), .DIN3(n6348), .DIN4(n6349), 
        .Q(n6345) );
  nor2s1 U7262 ( .DIN1(n6350), .DIN2(n6351), .Q(n6349) );
  nor2s1 U7263 ( .DIN1(n9469), .DIN2(n5427), .Q(n6351) );
  nor2s1 U7264 ( .DIN1(n9485), .DIN2(n5428), .Q(n6350) );
  nnd2s1 U7265 ( .DIN1(n5394), .DIN2(\DM_addr[22] ), .Q(n6348) );
  nnd2s1 U7266 ( .DIN1(n411), .DIN2(n6352), .Q(n6347) );
  nnd4s1 U7267 ( .DIN1(n6353), .DIN2(n6354), .DIN3(n6355), .DIN4(n6356), 
        .Q(n6352) );
  nor2s1 U7268 ( .DIN1(n405), .DIN2(n6357), .Q(n6356) );
  nor2s1 U7269 ( .DIN1(n5290), .DIN2(n6358), .Q(n6357) );
  nnd2s1 U7270 ( .DIN1(n5405), .DIN2(n121), .Q(n6355) );
  nnd2s1 U7271 ( .DIN1(n548), .DIN2(n6336), .Q(n6354) );
  nnd2s1 U7272 ( .DIN1(n5406), .DIN2(n6335), .Q(n6353) );
  nnd2s1 U7273 ( .DIN1(n6359), .DIN2(n67), .Q(n6346) );
  nnd3s1 U7274 ( .DIN1(n6360), .DIN2(n6361), .DIN3(n6362), .Q(n6359) );
  nnd2s1 U7275 ( .DIN1(n385), .DIN2(n6358), .Q(n6362) );
  xor2s1 U7276 ( .DIN1(n6340), .DIN2(n6341), .Q(n6358) );
  xnr2s1 U7277 ( .DIN1(n9469), .DIN2(n785), .Q(n6341) );
  and2s1 U7278 ( .DIN1(n6363), .DIN2(n6364), .Q(n6340) );
  nnd2s1 U7279 ( .DIN1(n412), .DIN2(n6365), .Q(n6364) );
  or2s1 U7280 ( .DIN1(n6366), .DIN2(n6367), .Q(n6365) );
  nnd2s1 U7281 ( .DIN1(n6367), .DIN2(n6366), .Q(n6363) );
  nnd2s1 U7282 ( .DIN1(n5406), .DIN2(n6336), .Q(n6361) );
  nnd2s1 U7283 ( .DIN1(n549), .DIN2(n6335), .Q(n6360) );
  hi1s1 U7284 ( .DIN(n6336), .Q(n6335) );
  nnd2s1 U7285 ( .DIN1(n6368), .DIN2(n6369), .Q(n6336) );
  nnd2s1 U7286 ( .DIN1(n412), .DIN2(n6370), .Q(n6369) );
  nnd2s1 U7287 ( .DIN1(n6371), .DIN2(n5426), .Q(n6370) );
  nnd2s1 U7288 ( .DIN1(n5423), .DIN2(n6372), .Q(n6368) );
  nnd3s1 U7289 ( .DIN1(n6373), .DIN2(n6374), .DIN3(n6375), .Q(n6344) );
  nnd2s1 U7290 ( .DIN1(n6376), .DIN2(n5665), .Q(n6375) );
  nnd3s1 U7291 ( .DIN1(n6377), .DIN2(n6378), .DIN3(n5946), .Q(n6374) );
  and3s1 U7292 ( .DIN1(n6379), .DIN2(n6380), .DIN3(n6035), .Q(n5946) );
  nnd2s1 U7293 ( .DIN1(n9486), .DIN2(n6381), .Q(n6378) );
  nnd4s1 U7294 ( .DIN1(n6382), .DIN2(n6383), .DIN3(n6384), .DIN4(n5553), 
        .Q(n6381) );
  nnd2s1 U7295 ( .DIN1(n6385), .DIN2(n398), .Q(n6384) );
  nnd2s1 U7296 ( .DIN1(n6386), .DIN2(n700), .Q(n6383) );
  nnd2s1 U7297 ( .DIN1(n6387), .DIN2(n5949), .Q(n6382) );
  or3s1 U7298 ( .DIN1(n5550), .DIN2(n5321), .DIN3(n9486), .Q(n6377) );
  nor2s1 U7299 ( .DIN1(n5741), .DIN2(n711), .Q(n5550) );
  nnd2s1 U7300 ( .DIN1(n6388), .DIN2(n6389), .Q(n6373) );
  nnd4s1 U7301 ( .DIN1(n6390), .DIN2(n6391), .DIN3(n6392), .DIN4(n6393), 
        .Q(n6389) );
  nor2s1 U7302 ( .DIN1(n6394), .DIN2(n805), .Q(n6393) );
  and2s1 U7303 ( .DIN1(n5536), .DIN2(n554), .Q(n6394) );
  nnd4s1 U7304 ( .DIN1(n6395), .DIN2(n6396), .DIN3(n6397), .DIN4(n6398), 
        .Q(n5536) );
  nnd2s1 U7305 ( .DIN1(n544), .DIN2(n5535), .Q(n6392) );
  nnd2s1 U7306 ( .DIN1(n5824), .DIN2(n6399), .Q(n6391) );
  nnd2s1 U7307 ( .DIN1(n726), .DIN2(n5959), .Q(n6390) );
  nnd2s1 U7308 ( .DIN1(n5547), .DIN2(n6400), .Q(n6388) );
  nnd2s1 U7309 ( .DIN1(n6401), .DIN2(n5301), .Q(n6400) );
  and2s1 U7310 ( .DIN1(n782), .DIN2(n6402), .Q(n6343) );
  nnd4s1 U7311 ( .DIN1(n6403), .DIN2(n6404), .DIN3(n6405), .DIN4(n6406), 
        .Q(n6402) );
  and4s1 U7312 ( .DIN1(n6407), .DIN2(n6408), .DIN3(n6409), .DIN4(n6410), 
        .Q(n6406) );
  nnd2s1 U7313 ( .DIN1(n6411), .DIN2(n6412), .Q(n6410) );
  nnd3s1 U7314 ( .DIN1(n6413), .DIN2(n5372), .DIN3(n6414), .Q(n6411) );
  nnd2s1 U7315 ( .DIN1(n620), .DIN2(n6287), .Q(n6414) );
  nnd2s1 U7316 ( .DIN1(n656), .DIN2(n6282), .Q(n6413) );
  hi1s1 U7317 ( .DIN(n6283), .Q(n6282) );
  nnd2s1 U7318 ( .DIN1(n6415), .DIN2(n6416), .Q(n6409) );
  nnd2s1 U7319 ( .DIN1(n6417), .DIN2(n6418), .Q(n6416) );
  nnd2s1 U7320 ( .DIN1(n655), .DIN2(n6283), .Q(n6418) );
  nnd2s1 U7321 ( .DIN1(n6419), .DIN2(n6420), .Q(n6283) );
  nnd2s1 U7322 ( .DIN1(reg_out_B[21]), .DIN2(n6421), .Q(n6420) );
  nnd2s1 U7323 ( .DIN1(n6422), .DIN2(n78), .Q(n6421) );
  nnd2s1 U7324 ( .DIN1(n412), .DIN2(n6423), .Q(n6419) );
  or2s1 U7325 ( .DIN1(n6287), .DIN2(n706), .Q(n6417) );
  nnd2s1 U7326 ( .DIN1(n6424), .DIN2(n6425), .Q(n6287) );
  nnd2s1 U7327 ( .DIN1(n6426), .DIN2(n6427), .Q(n6425) );
  nnd2s1 U7328 ( .DIN1(n5468), .DIN2(n6428), .Q(n6408) );
  nnd2s1 U7329 ( .DIN1(n411), .DIN2(n768), .Q(n6407) );
  nnd2s1 U7330 ( .DIN1(reg_out_B[22]), .DIN2(n6429), .Q(n6405) );
  nnd2s1 U7331 ( .DIN1(n723), .DIN2(n6430), .Q(n6429) );
  nnd2s1 U7332 ( .DIN1(n775), .DIN2(n411), .Q(n6430) );
  nnd3s1 U7333 ( .DIN1(n6431), .DIN2(n6432), .DIN3(n5336), .Q(n6404) );
  nnd2s1 U7334 ( .DIN1(n6433), .DIN2(n6434), .Q(n6432) );
  nnd2s1 U7335 ( .DIN1(n6435), .DIN2(n5478), .Q(n6434) );
  nnd2s1 U7336 ( .DIN1(n6436), .DIN2(n6437), .Q(n6431) );
  nnd2s1 U7337 ( .DIN1(n5480), .DIN2(n714), .Q(n6437) );
  nnd2s1 U7338 ( .DIN1(n6438), .DIN2(n6439), .Q(n6403) );
  nnd4s1 U7339 ( .DIN1(n6440), .DIN2(n6441), .DIN3(n6442), .DIN4(n6443), 
        .Q(n6439) );
  nnd2s1 U7340 ( .DIN1(n547), .DIN2(n6011), .Q(n6443) );
  nor2s1 U7341 ( .DIN1(n753), .DIN2(n6444), .Q(n6442) );
  and2s1 U7342 ( .DIN1(n6445), .DIN2(n720), .Q(n6444) );
  nnd2s1 U7343 ( .DIN1(n623), .DIN2(n5499), .Q(n6441) );
  nnd2s1 U7344 ( .DIN1(n629), .DIN2(n5500), .Q(n6440) );
  nnd4s1 U7345 ( .DIN1(n6446), .DIN2(n6447), .DIN3(n6448), .DIN4(n6449), 
        .Q(n5500) );
  nnd2s1 U7346 ( .DIN1(n5342), .DIN2(n6450), .Q(n6438) );
  nnd2s1 U7347 ( .DIN1(n6451), .DIN2(n387), .Q(n6450) );
  nor2s1 U7348 ( .DIN1(n6452), .DIN2(n5558), .Q(n6342) );
  or4s1 U7349 ( .DIN1(n6453), .DIN2(n6454), .DIN3(n6455), .DIN4(n6456), 
        .Q(\EXinst/n1453 ) );
  nnd4s1 U7350 ( .DIN1(n6457), .DIN2(n6458), .DIN3(n6459), .DIN4(n6460), 
        .Q(n6456) );
  nnd4s1 U7351 ( .DIN1(n6035), .DIN2(n6379), .DIN3(n6461), .DIN4(n6462), 
        .Q(n6460) );
  nnd2s1 U7352 ( .DIN1(n6463), .DIN2(n6464), .Q(n6462) );
  nnd3s1 U7353 ( .DIN1(n739), .DIN2(n5313), .DIN3(n6465), .Q(n6464) );
  nnd2s1 U7354 ( .DIN1(n6030), .DIN2(n6466), .Q(n6461) );
  nnd2s1 U7355 ( .DIN1(n6467), .DIN2(n5553), .Q(n6466) );
  nnd2s1 U7356 ( .DIN1(n6468), .DIN2(n6469), .Q(n6459) );
  nnd4s1 U7357 ( .DIN1(n6470), .DIN2(n6471), .DIN3(n6472), .DIN4(n6473), 
        .Q(n6469) );
  nor2s1 U7358 ( .DIN1(n6474), .DIN2(n806), .Q(n6473) );
  and2s1 U7359 ( .DIN1(n5587), .DIN2(n555), .Q(n6474) );
  nnd4s1 U7360 ( .DIN1(n6475), .DIN2(n6476), .DIN3(n6477), .DIN4(n6478), 
        .Q(n5587) );
  nnd2s1 U7361 ( .DIN1(n545), .DIN2(n5586), .Q(n6472) );
  nnd2s1 U7362 ( .DIN1(n5824), .DIN2(n6479), .Q(n6471) );
  nnd2s1 U7363 ( .DIN1(n726), .DIN2(n6044), .Q(n6470) );
  nnd2s1 U7364 ( .DIN1(n5547), .DIN2(n6480), .Q(n6468) );
  nnd3s1 U7365 ( .DIN1(n9487), .DIN2(n6481), .DIN3(n5301), .Q(n6480) );
  nnd2s1 U7366 ( .DIN1(n5570), .DIN2(n6482), .Q(n6458) );
  nnd2s1 U7367 ( .DIN1(n782), .DIN2(n6483), .Q(n6457) );
  nnd4s1 U7368 ( .DIN1(n6484), .DIN2(n6485), .DIN3(n6486), .DIN4(n6487), 
        .Q(n6483) );
  and4s1 U7369 ( .DIN1(n6488), .DIN2(n6489), .DIN3(n6490), .DIN4(n6491), 
        .Q(n6487) );
  nnd2s1 U7370 ( .DIN1(n6492), .DIN2(n6493), .Q(n6491) );
  nnd3s1 U7371 ( .DIN1(n6494), .DIN2(n749), .DIN3(n6495), .Q(n6492) );
  nnd2s1 U7372 ( .DIN1(n705), .DIN2(n6426), .Q(n6495) );
  nnd2s1 U7373 ( .DIN1(n654), .DIN2(n6422), .Q(n6494) );
  hi1s1 U7374 ( .DIN(n6423), .Q(n6422) );
  nnd2s1 U7375 ( .DIN1(n6496), .DIN2(n6497), .Q(n6490) );
  nnd2s1 U7376 ( .DIN1(n6498), .DIN2(n6499), .Q(n6497) );
  nnd2s1 U7377 ( .DIN1(n653), .DIN2(n6423), .Q(n6499) );
  nnd2s1 U7378 ( .DIN1(n6500), .DIN2(n6501), .Q(n6423) );
  nnd2s1 U7379 ( .DIN1(reg_out_B[20]), .DIN2(n6502), .Q(n6501) );
  nnd2s1 U7380 ( .DIN1(n6503), .DIN2(n69), .Q(n6502) );
  nnd2s1 U7381 ( .DIN1(n413), .DIN2(n6504), .Q(n6500) );
  or2s1 U7382 ( .DIN1(n6426), .DIN2(n5375), .Q(n6498) );
  nnd2s1 U7383 ( .DIN1(n6505), .DIN2(n6506), .Q(n6426) );
  nnd2s1 U7384 ( .DIN1(n6507), .DIN2(n6508), .Q(n6506) );
  nnd2s1 U7385 ( .DIN1(n5468), .DIN2(n6509), .Q(n6489) );
  nnd2s1 U7386 ( .DIN1(n412), .DIN2(n767), .Q(n6488) );
  nnd2s1 U7387 ( .DIN1(reg_out_B[21]), .DIN2(n6510), .Q(n6486) );
  nnd2s1 U7388 ( .DIN1(n723), .DIN2(n6511), .Q(n6510) );
  nnd2s1 U7389 ( .DIN1(n776), .DIN2(n412), .Q(n6511) );
  nnd3s1 U7390 ( .DIN1(n6512), .DIN2(n6513), .DIN3(n769), .Q(n6485) );
  nnd2s1 U7391 ( .DIN1(n6436), .DIN2(n6514), .Q(n6513) );
  nnd2s1 U7392 ( .DIN1(n5480), .DIN2(n211), .Q(n6514) );
  nnd2s1 U7393 ( .DIN1(n6433), .DIN2(n6515), .Q(n6512) );
  nnd2s1 U7394 ( .DIN1(n6516), .DIN2(n5478), .Q(n6515) );
  nnd2s1 U7395 ( .DIN1(n6517), .DIN2(n6518), .Q(n6484) );
  nnd4s1 U7396 ( .DIN1(n6519), .DIN2(n6520), .DIN3(n6521), .DIN4(n6522), 
        .Q(n6518) );
  nnd2s1 U7397 ( .DIN1(n546), .DIN2(n6095), .Q(n6522) );
  nor2s1 U7398 ( .DIN1(n55), .DIN2(n6523), .Q(n6521) );
  and2s1 U7399 ( .DIN1(n6524), .DIN2(n720), .Q(n6523) );
  nnd2s1 U7400 ( .DIN1(n622), .DIN2(n5643), .Q(n6520) );
  nnd2s1 U7401 ( .DIN1(n630), .DIN2(n5644), .Q(n6519) );
  nnd4s1 U7402 ( .DIN1(n6525), .DIN2(n6526), .DIN3(n6527), .DIN4(n6528), 
        .Q(n5644) );
  nnd2s1 U7403 ( .DIN1(n5342), .DIN2(n6529), .Q(n6517) );
  nnd3s1 U7404 ( .DIN1(n6530), .DIN2(n801), .DIN3(n387), .Q(n6529) );
  nnd3s1 U7405 ( .DIN1(n6531), .DIN2(n6532), .DIN3(n6533), .Q(n6455) );
  nnd2s1 U7406 ( .DIN1(n727), .DIN2(\DM_addr[21] ), .Q(n6533) );
  nnd2s1 U7407 ( .DIN1(n412), .DIN2(n6534), .Q(n6532) );
  or3s1 U7408 ( .DIN1(n402), .DIN2(n6535), .DIN3(n6536), .Q(n6534) );
  nnd4s1 U7409 ( .DIN1(n6537), .DIN2(n6538), .DIN3(n6539), .DIN4(n6540), 
        .Q(n6536) );
  nnd2s1 U7410 ( .DIN1(n548), .DIN2(n6372), .Q(n6540) );
  nnd2s1 U7411 ( .DIN1(n5406), .DIN2(n6371), .Q(n6539) );
  nnd2s1 U7412 ( .DIN1(n5405), .DIN2(n16), .Q(n6538) );
  nnd2s1 U7413 ( .DIN1(n5665), .DIN2(n9470), .Q(n6537) );
  nor2s1 U7414 ( .DIN1(n5290), .DIN2(n6541), .Q(n6535) );
  nnd2s1 U7415 ( .DIN1(n6542), .DIN2(n78), .Q(n6531) );
  nnd4s1 U7416 ( .DIN1(n6543), .DIN2(n6544), .DIN3(n6545), .DIN4(n6546), 
        .Q(n6542) );
  nnd2s1 U7417 ( .DIN1(n5406), .DIN2(n6372), .Q(n6546) );
  nnd2s1 U7418 ( .DIN1(n549), .DIN2(n6371), .Q(n6545) );
  hi1s1 U7419 ( .DIN(n6372), .Q(n6371) );
  nnd2s1 U7420 ( .DIN1(n6547), .DIN2(n6548), .Q(n6372) );
  nnd2s1 U7421 ( .DIN1(n413), .DIN2(n6549), .Q(n6548) );
  nnd2s1 U7422 ( .DIN1(n6550), .DIN2(n5426), .Q(n6549) );
  nnd2s1 U7423 ( .DIN1(n633), .DIN2(n6551), .Q(n6547) );
  nnd2s1 U7424 ( .DIN1(n385), .DIN2(n6541), .Q(n6544) );
  xor2s1 U7425 ( .DIN1(n6366), .DIN2(n6367), .Q(n6541) );
  xor2s1 U7426 ( .DIN1(n16), .DIN2(n5413), .Q(n6367) );
  nnd2s1 U7427 ( .DIN1(n6552), .DIN2(n6553), .Q(n6366) );
  nnd2s1 U7428 ( .DIN1(n413), .DIN2(n6554), .Q(n6553) );
  nnd2s1 U7429 ( .DIN1(n6555), .DIN2(n6556), .Q(n6554) );
  or2s1 U7430 ( .DIN1(n6556), .DIN2(n6555), .Q(n6552) );
  nnd2s1 U7431 ( .DIN1(n5665), .DIN2(n16), .Q(n6543) );
  nor2s1 U7432 ( .DIN1(n9470), .DIN2(n5427), .Q(n6454) );
  nor2s1 U7433 ( .DIN1(n9486), .DIN2(n5428), .Q(n6453) );
  or4s1 U7434 ( .DIN1(n6557), .DIN2(n6558), .DIN3(n6559), .DIN4(n6560), 
        .Q(\EXinst/n1452 ) );
  nnd4s1 U7435 ( .DIN1(n6561), .DIN2(n6562), .DIN3(n6563), .DIN4(n6564), 
        .Q(n6560) );
  nor2s1 U7436 ( .DIN1(n6565), .DIN2(n6566), .Q(n6564) );
  nor2s1 U7437 ( .DIN1(n9471), .DIN2(n5427), .Q(n6566) );
  nor2s1 U7438 ( .DIN1(n740), .DIN2(n5428), .Q(n6565) );
  nnd2s1 U7439 ( .DIN1(n5394), .DIN2(\DM_addr[20] ), .Q(n6563) );
  nnd2s1 U7440 ( .DIN1(n413), .DIN2(n6567), .Q(n6562) );
  nnd4s1 U7441 ( .DIN1(n6568), .DIN2(n6569), .DIN3(n6570), .DIN4(n6571), 
        .Q(n6567) );
  nor2s1 U7442 ( .DIN1(n404), .DIN2(n6572), .Q(n6571) );
  nor2s1 U7443 ( .DIN1(n5290), .DIN2(n6573), .Q(n6572) );
  nnd2s1 U7444 ( .DIN1(n5405), .DIN2(n123), .Q(n6570) );
  nnd2s1 U7445 ( .DIN1(n548), .DIN2(n6551), .Q(n6569) );
  nnd2s1 U7446 ( .DIN1(n5406), .DIN2(n6550), .Q(n6568) );
  nnd2s1 U7447 ( .DIN1(n6574), .DIN2(n69), .Q(n6561) );
  nnd3s1 U7448 ( .DIN1(n6575), .DIN2(n6576), .DIN3(n6577), .Q(n6574) );
  nnd2s1 U7449 ( .DIN1(n385), .DIN2(n6573), .Q(n6577) );
  xor2s1 U7450 ( .DIN1(n6555), .DIN2(n6556), .Q(n6573) );
  xnr2s1 U7451 ( .DIN1(n9471), .DIN2(n5514), .Q(n6556) );
  and2s1 U7452 ( .DIN1(n6578), .DIN2(n6579), .Q(n6555) );
  nnd2s1 U7453 ( .DIN1(n414), .DIN2(n6580), .Q(n6579) );
  or2s1 U7454 ( .DIN1(n6581), .DIN2(n6582), .Q(n6580) );
  nnd2s1 U7455 ( .DIN1(n6582), .DIN2(n6581), .Q(n6578) );
  nnd2s1 U7456 ( .DIN1(n5406), .DIN2(n6551), .Q(n6576) );
  nnd2s1 U7457 ( .DIN1(n549), .DIN2(n6550), .Q(n6575) );
  hi1s1 U7458 ( .DIN(n6551), .Q(n6550) );
  nnd2s1 U7459 ( .DIN1(n6583), .DIN2(n6584), .Q(n6551) );
  nnd2s1 U7460 ( .DIN1(n414), .DIN2(n6585), .Q(n6584) );
  nnd2s1 U7461 ( .DIN1(n6586), .DIN2(n5426), .Q(n6585) );
  nnd2s1 U7462 ( .DIN1(n5423), .DIN2(n6587), .Q(n6583) );
  nnd3s1 U7463 ( .DIN1(n6588), .DIN2(n6589), .DIN3(n6590), .Q(n6559) );
  nnd2s1 U7464 ( .DIN1(n6591), .DIN2(n5665), .Q(n6590) );
  nnd2s1 U7465 ( .DIN1(n6592), .DIN2(n6593), .Q(n6589) );
  nnd2s1 U7466 ( .DIN1(n6030), .DIN2(n6594), .Q(n6593) );
  nnd2s1 U7467 ( .DIN1(n6595), .DIN2(n5553), .Q(n6594) );
  nnd2s1 U7468 ( .DIN1(n6168), .DIN2(n6596), .Q(n6592) );
  nnd2s1 U7469 ( .DIN1(n5322), .DIN2(n6465), .Q(n6596) );
  nnd2s1 U7470 ( .DIN1(n6597), .DIN2(n6598), .Q(n6588) );
  nnd4s1 U7471 ( .DIN1(n6599), .DIN2(n6600), .DIN3(n6601), .DIN4(n6602), 
        .Q(n6598) );
  nor2s1 U7472 ( .DIN1(n6603), .DIN2(n806), .Q(n6602) );
  and2s1 U7473 ( .DIN1(n5724), .DIN2(n554), .Q(n6603) );
  nnd4s1 U7474 ( .DIN1(n6604), .DIN2(n6605), .DIN3(n6606), .DIN4(n6607), 
        .Q(n5724) );
  nnd2s1 U7475 ( .DIN1(n544), .DIN2(n5723), .Q(n6601) );
  nnd2s1 U7476 ( .DIN1(n5824), .DIN2(n6608), .Q(n6600) );
  nnd2s1 U7477 ( .DIN1(n5826), .DIN2(n6176), .Q(n6599) );
  nnd2s1 U7478 ( .DIN1(n5547), .DIN2(n6609), .Q(n6597) );
  nnd3s1 U7479 ( .DIN1(n9487), .DIN2(n6610), .DIN3(n5301), .Q(n6609) );
  and2s1 U7480 ( .DIN1(n782), .DIN2(n6611), .Q(n6558) );
  nnd4s1 U7481 ( .DIN1(n6612), .DIN2(n6613), .DIN3(n6614), .DIN4(n6615), 
        .Q(n6611) );
  and4s1 U7482 ( .DIN1(n6616), .DIN2(n6617), .DIN3(n6618), .DIN4(n6619), 
        .Q(n6615) );
  nnd2s1 U7483 ( .DIN1(n6620), .DIN2(n6621), .Q(n6619) );
  nnd3s1 U7484 ( .DIN1(n6622), .DIN2(n5372), .DIN3(n6623), .Q(n6620) );
  nnd2s1 U7485 ( .DIN1(n620), .DIN2(n6508), .Q(n6623) );
  nnd2s1 U7486 ( .DIN1(n656), .DIN2(n6503), .Q(n6622) );
  hi1s1 U7487 ( .DIN(n6504), .Q(n6503) );
  nnd2s1 U7488 ( .DIN1(n6624), .DIN2(n6625), .Q(n6618) );
  nnd2s1 U7489 ( .DIN1(n6626), .DIN2(n6627), .Q(n6625) );
  nnd2s1 U7490 ( .DIN1(n655), .DIN2(n6504), .Q(n6627) );
  nnd2s1 U7491 ( .DIN1(n6628), .DIN2(n6629), .Q(n6504) );
  nnd2s1 U7492 ( .DIN1(reg_out_B[19]), .DIN2(n6630), .Q(n6629) );
  nnd2s1 U7493 ( .DIN1(n6631), .DIN2(n37), .Q(n6630) );
  nnd2s1 U7494 ( .DIN1(n414), .DIN2(n6632), .Q(n6628) );
  or2s1 U7495 ( .DIN1(n6508), .DIN2(n706), .Q(n6626) );
  nnd2s1 U7496 ( .DIN1(n6633), .DIN2(n6634), .Q(n6508) );
  nnd2s1 U7497 ( .DIN1(n6635), .DIN2(n6636), .Q(n6634) );
  nnd2s1 U7498 ( .DIN1(n5468), .DIN2(n6637), .Q(n6617) );
  nnd2s1 U7499 ( .DIN1(n413), .DIN2(n768), .Q(n6616) );
  nnd2s1 U7500 ( .DIN1(reg_out_B[20]), .DIN2(n6638), .Q(n6614) );
  nnd2s1 U7501 ( .DIN1(n723), .DIN2(n6639), .Q(n6638) );
  nnd2s1 U7502 ( .DIN1(n775), .DIN2(n413), .Q(n6639) );
  nnd3s1 U7503 ( .DIN1(n6640), .DIN2(n6641), .DIN3(n5336), .Q(n6613) );
  nnd2s1 U7504 ( .DIN1(n6433), .DIN2(n6642), .Q(n6641) );
  nnd2s1 U7505 ( .DIN1(n6643), .DIN2(n5478), .Q(n6642) );
  hi1s1 U7506 ( .DIN(n6644), .Q(n6640) );
  nnd2s1 U7507 ( .DIN1(n6645), .DIN2(n6646), .Q(n6612) );
  nnd4s1 U7508 ( .DIN1(n6647), .DIN2(n6648), .DIN3(n6649), .DIN4(n6650), 
        .Q(n6646) );
  nnd2s1 U7509 ( .DIN1(n547), .DIN2(n6224), .Q(n6650) );
  nor2s1 U7510 ( .DIN1(n752), .DIN2(n6651), .Q(n6649) );
  and2s1 U7511 ( .DIN1(n6652), .DIN2(n720), .Q(n6651) );
  nnd2s1 U7512 ( .DIN1(n621), .DIN2(n5791), .Q(n6648) );
  nnd2s1 U7513 ( .DIN1(n629), .DIN2(n5792), .Q(n6647) );
  nnd4s1 U7514 ( .DIN1(n6653), .DIN2(n6654), .DIN3(n6655), .DIN4(n6656), 
        .Q(n5792) );
  nnd2s1 U7515 ( .DIN1(n5342), .DIN2(n6657), .Q(n6645) );
  nnd3s1 U7516 ( .DIN1(n6658), .DIN2(n337), .DIN3(n387), .Q(n6657) );
  nor2s1 U7517 ( .DIN1(n6659), .DIN2(n5558), .Q(n6557) );
  or4s1 U7518 ( .DIN1(n6660), .DIN2(n6661), .DIN3(n6662), .DIN4(n6663), 
        .Q(\EXinst/n1451 ) );
  nnd4s1 U7519 ( .DIN1(n6664), .DIN2(n6665), .DIN3(n6666), .DIN4(n6667), 
        .Q(n6663) );
  nnd2s1 U7520 ( .DIN1(n6668), .DIN2(n6669), .Q(n6667) );
  nnd2s1 U7521 ( .DIN1(n6030), .DIN2(n6670), .Q(n6669) );
  nnd2s1 U7522 ( .DIN1(n6671), .DIN2(n5553), .Q(n6670) );
  nnd2s1 U7523 ( .DIN1(n6672), .DIN2(n6673), .Q(n6671) );
  nnd2s1 U7524 ( .DIN1(n6168), .DIN2(n6674), .Q(n6668) );
  nnd2s1 U7525 ( .DIN1(n5322), .DIN2(n5811), .Q(n6674) );
  nnd2s1 U7526 ( .DIN1(n6675), .DIN2(n6676), .Q(n6666) );
  nnd4s1 U7527 ( .DIN1(n6677), .DIN2(n6678), .DIN3(n6679), .DIN4(n6680), 
        .Q(n6676) );
  nor2s1 U7528 ( .DIN1(n6681), .DIN2(n805), .Q(n6680) );
  nor2s1 U7529 ( .DIN1(n5305), .DIN2(n6253), .Q(n6681) );
  hi1s1 U7530 ( .DIN(n5827), .Q(n5305) );
  nnd4s1 U7531 ( .DIN1(n6682), .DIN2(n6683), .DIN3(n6684), .DIN4(n6685), 
        .Q(n5827) );
  nnd2s1 U7532 ( .DIN1(n545), .DIN2(n5825), .Q(n6679) );
  nnd2s1 U7533 ( .DIN1(n5824), .DIN2(n6686), .Q(n6678) );
  nnd2s1 U7534 ( .DIN1(n5826), .DIN2(n6258), .Q(n6677) );
  nnd2s1 U7535 ( .DIN1(n5547), .DIN2(n6687), .Q(n6675) );
  nnd2s1 U7536 ( .DIN1(n6688), .DIN2(n6689), .Q(n6687) );
  nnd2s1 U7537 ( .DIN1(n5570), .DIN2(n6690), .Q(n6665) );
  nnd2s1 U7538 ( .DIN1(n782), .DIN2(n6691), .Q(n6664) );
  nnd4s1 U7539 ( .DIN1(n6692), .DIN2(n6693), .DIN3(n6694), .DIN4(n6695), 
        .Q(n6691) );
  and4s1 U7540 ( .DIN1(n6696), .DIN2(n6697), .DIN3(n6698), .DIN4(n6699), 
        .Q(n6695) );
  nnd2s1 U7541 ( .DIN1(n6700), .DIN2(n6701), .Q(n6699) );
  nnd3s1 U7542 ( .DIN1(n6702), .DIN2(n749), .DIN3(n6703), .Q(n6700) );
  nnd2s1 U7543 ( .DIN1(n705), .DIN2(n6635), .Q(n6703) );
  nnd2s1 U7544 ( .DIN1(n654), .DIN2(n6631), .Q(n6702) );
  hi1s1 U7545 ( .DIN(n6632), .Q(n6631) );
  nnd2s1 U7546 ( .DIN1(n6704), .DIN2(n6705), .Q(n6698) );
  nnd2s1 U7547 ( .DIN1(n6706), .DIN2(n6707), .Q(n6705) );
  nnd2s1 U7548 ( .DIN1(n653), .DIN2(n6632), .Q(n6707) );
  nnd2s1 U7549 ( .DIN1(n6708), .DIN2(n6709), .Q(n6632) );
  nnd2s1 U7550 ( .DIN1(reg_out_B[18]), .DIN2(n6710), .Q(n6709) );
  nnd2s1 U7551 ( .DIN1(n6711), .DIN2(n70), .Q(n6710) );
  nnd2s1 U7552 ( .DIN1(n415), .DIN2(n6712), .Q(n6708) );
  or2s1 U7553 ( .DIN1(n6635), .DIN2(n706), .Q(n6706) );
  nnd2s1 U7554 ( .DIN1(n6713), .DIN2(n6714), .Q(n6635) );
  nnd2s1 U7555 ( .DIN1(n6715), .DIN2(n6716), .Q(n6714) );
  nnd2s1 U7556 ( .DIN1(n5468), .DIN2(n6717), .Q(n6697) );
  nnd2s1 U7557 ( .DIN1(n414), .DIN2(n767), .Q(n6696) );
  nnd2s1 U7558 ( .DIN1(reg_out_B[19]), .DIN2(n6718), .Q(n6694) );
  nnd2s1 U7559 ( .DIN1(n5471), .DIN2(n6719), .Q(n6718) );
  nnd2s1 U7560 ( .DIN1(n776), .DIN2(n414), .Q(n6719) );
  nnd3s1 U7561 ( .DIN1(n6720), .DIN2(n6721), .DIN3(n6293), .Q(n6693) );
  and3s1 U7562 ( .DIN1(n5478), .DIN2(n6722), .DIN3(n5336), .Q(n6293) );
  hi1s1 U7563 ( .DIN(n6723), .Q(n6722) );
  nnd4s1 U7564 ( .DIN1(n6724), .DIN2(n807), .DIN3(n6725), .DIN4(n5337), 
        .Q(n6721) );
  nnd3s1 U7565 ( .DIN1(n6726), .DIN2(n6727), .DIN3(n337), .Q(n6725) );
  or2s1 U7566 ( .DIN1(n6728), .DIN2(n742), .Q(n6727) );
  nnd2s1 U7567 ( .DIN1(n6298), .DIN2(n741), .Q(n6726) );
  hi1s1 U7568 ( .DIN(n6729), .Q(n6298) );
  nnd3s1 U7569 ( .DIN1(n6730), .DIN2(n6301), .DIN3(reg_out_B[5]), .Q(n6720) );
  nnd2s1 U7570 ( .DIN1(n6731), .DIN2(n6732), .Q(n6692) );
  nnd4s1 U7571 ( .DIN1(n6733), .DIN2(n6734), .DIN3(n6735), .DIN4(n6736), 
        .Q(n6732) );
  nnd2s1 U7572 ( .DIN1(n546), .DIN2(n6309), .Q(n6736) );
  nor2s1 U7573 ( .DIN1(n753), .DIN2(n6737), .Q(n6735) );
  nor2s1 U7574 ( .DIN1(n6738), .DIN2(n5359), .Q(n6737) );
  nnd2s1 U7575 ( .DIN1(n623), .DIN2(n5875), .Q(n6734) );
  nnd2s1 U7576 ( .DIN1(n630), .DIN2(n5360), .Q(n6733) );
  nnd4s1 U7577 ( .DIN1(n6739), .DIN2(n6740), .DIN3(n6741), .DIN4(n6742), 
        .Q(n5360) );
  nnd2s1 U7578 ( .DIN1(n5342), .DIN2(n6743), .Q(n6731) );
  nnd2s1 U7579 ( .DIN1(n6744), .DIN2(n6745), .Q(n6743) );
  nnd3s1 U7580 ( .DIN1(n6746), .DIN2(n6747), .DIN3(n6748), .Q(n6662) );
  nnd2s1 U7581 ( .DIN1(n727), .DIN2(\DM_addr[19] ), .Q(n6748) );
  nnd2s1 U7582 ( .DIN1(n414), .DIN2(n6749), .Q(n6747) );
  or3s1 U7583 ( .DIN1(n402), .DIN2(n6750), .DIN3(n6751), .Q(n6749) );
  nnd4s1 U7584 ( .DIN1(n6752), .DIN2(n6753), .DIN3(n6754), .DIN4(n6755), 
        .Q(n6751) );
  nnd2s1 U7585 ( .DIN1(n548), .DIN2(n6587), .Q(n6755) );
  nnd2s1 U7586 ( .DIN1(n5406), .DIN2(n6586), .Q(n6754) );
  nnd2s1 U7587 ( .DIN1(n5405), .DIN2(n94), .Q(n6753) );
  nnd2s1 U7588 ( .DIN1(n5665), .DIN2(n9472), .Q(n6752) );
  nor2s1 U7589 ( .DIN1(n5290), .DIN2(n6756), .Q(n6750) );
  nnd2s1 U7590 ( .DIN1(n6757), .DIN2(n37), .Q(n6746) );
  nnd4s1 U7591 ( .DIN1(n6758), .DIN2(n6759), .DIN3(n6760), .DIN4(n6761), 
        .Q(n6757) );
  nnd2s1 U7592 ( .DIN1(n5406), .DIN2(n6587), .Q(n6761) );
  nnd2s1 U7593 ( .DIN1(n549), .DIN2(n6586), .Q(n6760) );
  hi1s1 U7594 ( .DIN(n6587), .Q(n6586) );
  nnd2s1 U7595 ( .DIN1(n6762), .DIN2(n6763), .Q(n6587) );
  nnd2s1 U7596 ( .DIN1(n415), .DIN2(n6764), .Q(n6763) );
  nnd2s1 U7597 ( .DIN1(n6765), .DIN2(n5426), .Q(n6764) );
  nnd2s1 U7598 ( .DIN1(n633), .DIN2(n6766), .Q(n6762) );
  nnd2s1 U7599 ( .DIN1(n385), .DIN2(n6756), .Q(n6759) );
  xor2s1 U7600 ( .DIN1(n6581), .DIN2(n6582), .Q(n6756) );
  xor2s1 U7601 ( .DIN1(n94), .DIN2(n745), .Q(n6582) );
  nnd2s1 U7602 ( .DIN1(n6767), .DIN2(n6768), .Q(n6581) );
  nnd2s1 U7603 ( .DIN1(n415), .DIN2(n6769), .Q(n6768) );
  nnd2s1 U7604 ( .DIN1(n6770), .DIN2(n6771), .Q(n6769) );
  or2s1 U7605 ( .DIN1(n6771), .DIN2(n6770), .Q(n6767) );
  nnd2s1 U7606 ( .DIN1(n5665), .DIN2(n94), .Q(n6758) );
  nor2s1 U7607 ( .DIN1(n9472), .DIN2(n5427), .Q(n6661) );
  nor2s1 U7608 ( .DIN1(n9487), .DIN2(n5428), .Q(n6660) );
  or4s1 U7609 ( .DIN1(n6772), .DIN2(n6773), .DIN3(n6774), .DIN4(n6775), 
        .Q(\EXinst/n1450 ) );
  nnd4s1 U7610 ( .DIN1(n6776), .DIN2(n6777), .DIN3(n6778), .DIN4(n6779), 
        .Q(n6775) );
  nor2s1 U7611 ( .DIN1(n6780), .DIN2(n6781), .Q(n6779) );
  nor2s1 U7612 ( .DIN1(n9473), .DIN2(n5427), .Q(n6781) );
  nor2s1 U7613 ( .DIN1(n29), .DIN2(n5428), .Q(n6780) );
  nnd2s1 U7614 ( .DIN1(n5394), .DIN2(\DM_addr[18] ), .Q(n6778) );
  nnd2s1 U7615 ( .DIN1(n415), .DIN2(n6782), .Q(n6777) );
  nnd4s1 U7616 ( .DIN1(n6783), .DIN2(n6784), .DIN3(n6785), .DIN4(n6786), 
        .Q(n6782) );
  nor2s1 U7617 ( .DIN1(n403), .DIN2(n6787), .Q(n6786) );
  nor2s1 U7618 ( .DIN1(n5290), .DIN2(n6788), .Q(n6787) );
  nnd2s1 U7619 ( .DIN1(n5405), .DIN2(n122), .Q(n6785) );
  nnd2s1 U7620 ( .DIN1(n548), .DIN2(n6766), .Q(n6784) );
  nnd2s1 U7621 ( .DIN1(n5406), .DIN2(n6765), .Q(n6783) );
  nnd2s1 U7622 ( .DIN1(n6789), .DIN2(n70), .Q(n6776) );
  nnd3s1 U7623 ( .DIN1(n6790), .DIN2(n6791), .DIN3(n6792), .Q(n6789) );
  nnd2s1 U7624 ( .DIN1(n385), .DIN2(n6788), .Q(n6792) );
  xor2s1 U7625 ( .DIN1(n6770), .DIN2(n6771), .Q(n6788) );
  xnr2s1 U7626 ( .DIN1(n9473), .DIN2(n786), .Q(n6771) );
  and2s1 U7627 ( .DIN1(n6793), .DIN2(n6794), .Q(n6770) );
  nnd2s1 U7628 ( .DIN1(n416), .DIN2(n6795), .Q(n6794) );
  or2s1 U7629 ( .DIN1(n6796), .DIN2(n6797), .Q(n6795) );
  nnd2s1 U7630 ( .DIN1(n6797), .DIN2(n6796), .Q(n6793) );
  nnd2s1 U7631 ( .DIN1(n5406), .DIN2(n6766), .Q(n6791) );
  nnd2s1 U7632 ( .DIN1(n549), .DIN2(n6765), .Q(n6790) );
  hi1s1 U7633 ( .DIN(n6766), .Q(n6765) );
  nnd2s1 U7634 ( .DIN1(n6798), .DIN2(n6799), .Q(n6766) );
  nnd2s1 U7635 ( .DIN1(n416), .DIN2(n6800), .Q(n6799) );
  nnd2s1 U7636 ( .DIN1(n6801), .DIN2(n5426), .Q(n6800) );
  nnd2s1 U7637 ( .DIN1(n5423), .DIN2(n6802), .Q(n6798) );
  nnd3s1 U7638 ( .DIN1(n6803), .DIN2(n6804), .DIN3(n6805), .Q(n6774) );
  nnd2s1 U7639 ( .DIN1(n6806), .DIN2(n5665), .Q(n6805) );
  nnd4s1 U7640 ( .DIN1(n6035), .DIN2(n6379), .DIN3(n6807), .DIN4(n6808), 
        .Q(n6804) );
  nnd2s1 U7641 ( .DIN1(n6463), .DIN2(n6809), .Q(n6808) );
  nnd2s1 U7642 ( .DIN1(n739), .DIN2(n6810), .Q(n6809) );
  nnd2s1 U7643 ( .DIN1(n5741), .DIN2(n5950), .Q(n6810) );
  nnd2s1 U7644 ( .DIN1(n712), .DIN2(reg_out_A[31]), .Q(n5950) );
  and2s1 U7645 ( .DIN1(n4831), .DIN2(n6811), .Q(n6463) );
  nnd2s1 U7646 ( .DIN1(n5321), .DIN2(n56), .Q(n6811) );
  nnd2s1 U7647 ( .DIN1(n6030), .DIN2(n6812), .Q(n6807) );
  nnd2s1 U7648 ( .DIN1(n6813), .DIN2(n5553), .Q(n6812) );
  nnd2s1 U7649 ( .DIN1(n6814), .DIN2(n6815), .Q(n6813) );
  nnd2s1 U7650 ( .DIN1(n6816), .DIN2(n4840), .Q(n6815) );
  nnd2s1 U7651 ( .DIN1(n6817), .DIN2(n6818), .Q(n6803) );
  nnd4s1 U7652 ( .DIN1(n6819), .DIN2(n6820), .DIN3(n6821), .DIN4(n6822), 
        .Q(n6818) );
  nor2s1 U7653 ( .DIN1(n6823), .DIN2(n806), .Q(n6822) );
  and2s1 U7654 ( .DIN1(n5535), .DIN2(n555), .Q(n6823) );
  nnd4s1 U7655 ( .DIN1(n6824), .DIN2(n6825), .DIN3(n6826), .DIN4(n6827), 
        .Q(n5535) );
  nnd2s1 U7656 ( .DIN1(n544), .DIN2(n5959), .Q(n6821) );
  nnd2s1 U7657 ( .DIN1(n5824), .DIN2(n6828), .Q(n6820) );
  nnd2s1 U7658 ( .DIN1(n5826), .DIN2(n6399), .Q(n6819) );
  nnd2s1 U7659 ( .DIN1(n5547), .DIN2(n6829), .Q(n6817) );
  nnd2s1 U7660 ( .DIN1(n6688), .DIN2(n6830), .Q(n6829) );
  and2s1 U7661 ( .DIN1(n782), .DIN2(n6831), .Q(n6773) );
  nnd4s1 U7662 ( .DIN1(n6832), .DIN2(n6833), .DIN3(n6834), .DIN4(n6835), 
        .Q(n6831) );
  and4s1 U7663 ( .DIN1(n6836), .DIN2(n6837), .DIN3(n6838), .DIN4(n6839), 
        .Q(n6835) );
  nnd2s1 U7664 ( .DIN1(n6840), .DIN2(n6841), .Q(n6839) );
  nnd3s1 U7665 ( .DIN1(n6842), .DIN2(n5372), .DIN3(n6843), .Q(n6840) );
  nnd2s1 U7666 ( .DIN1(n620), .DIN2(n6716), .Q(n6843) );
  nnd2s1 U7667 ( .DIN1(n656), .DIN2(n6711), .Q(n6842) );
  hi1s1 U7668 ( .DIN(n6712), .Q(n6711) );
  nnd2s1 U7669 ( .DIN1(n6844), .DIN2(n6845), .Q(n6838) );
  nnd2s1 U7670 ( .DIN1(n6846), .DIN2(n6847), .Q(n6845) );
  nnd2s1 U7671 ( .DIN1(n655), .DIN2(n6712), .Q(n6847) );
  nnd2s1 U7672 ( .DIN1(n6848), .DIN2(n6849), .Q(n6712) );
  nnd2s1 U7673 ( .DIN1(reg_out_B[17]), .DIN2(n6850), .Q(n6849) );
  nnd2s1 U7674 ( .DIN1(n6851), .DIN2(n82), .Q(n6850) );
  nnd2s1 U7675 ( .DIN1(n416), .DIN2(n6852), .Q(n6848) );
  or2s1 U7676 ( .DIN1(n6716), .DIN2(n706), .Q(n6846) );
  nnd2s1 U7677 ( .DIN1(n6853), .DIN2(n6854), .Q(n6716) );
  nnd2s1 U7678 ( .DIN1(n6855), .DIN2(n6856), .Q(n6854) );
  nnd2s1 U7679 ( .DIN1(n5468), .DIN2(n6857), .Q(n6837) );
  nnd2s1 U7680 ( .DIN1(n415), .DIN2(n768), .Q(n6836) );
  nnd2s1 U7681 ( .DIN1(reg_out_B[18]), .DIN2(n6858), .Q(n6834) );
  nnd2s1 U7682 ( .DIN1(n5471), .DIN2(n6859), .Q(n6858) );
  nnd2s1 U7683 ( .DIN1(n775), .DIN2(n415), .Q(n6859) );
  nnd3s1 U7684 ( .DIN1(n6860), .DIN2(n6861), .DIN3(n769), .Q(n6833) );
  nnd2s1 U7685 ( .DIN1(n6644), .DIN2(n6862), .Q(n6861) );
  nnd3s1 U7686 ( .DIN1(n714), .DIN2(n808), .DIN3(n734), .Q(n6862) );
  nor2s1 U7687 ( .DIN1(n6213), .DIN2(n5480), .Q(n6644) );
  nor2s1 U7688 ( .DIN1(n6863), .DIN2(n752), .Q(n5480) );
  hi1s1 U7689 ( .DIN(n6436), .Q(n6213) );
  nnd2s1 U7690 ( .DIN1(n6433), .DIN2(n6864), .Q(n6860) );
  nnd2s1 U7691 ( .DIN1(n6865), .DIN2(n5478), .Q(n6864) );
  nnd2s1 U7692 ( .DIN1(n6866), .DIN2(n6867), .Q(n6832) );
  nnd4s1 U7693 ( .DIN1(n6868), .DIN2(n6869), .DIN3(n6870), .DIN4(n6871), 
        .Q(n6867) );
  nnd2s1 U7694 ( .DIN1(n547), .DIN2(n6445), .Q(n6871) );
  nor2s1 U7695 ( .DIN1(n55), .DIN2(n6872), .Q(n6870) );
  nor2s1 U7696 ( .DIN1(n6873), .DIN2(n5359), .Q(n6872) );
  nnd2s1 U7697 ( .DIN1(n622), .DIN2(n6011), .Q(n6869) );
  nnd2s1 U7698 ( .DIN1(n629), .DIN2(n5499), .Q(n6868) );
  nnd4s1 U7699 ( .DIN1(n6874), .DIN2(n6875), .DIN3(n6876), .DIN4(n6877), 
        .Q(n5499) );
  nnd2s1 U7700 ( .DIN1(n5342), .DIN2(n6878), .Q(n6866) );
  nnd2s1 U7701 ( .DIN1(n6744), .DIN2(n6879), .Q(n6878) );
  nor2s1 U7702 ( .DIN1(n6880), .DIN2(n5558), .Q(n6772) );
  or4s1 U7703 ( .DIN1(n6881), .DIN2(n6882), .DIN3(n6883), .DIN4(n6884), 
        .Q(\EXinst/n1449 ) );
  nnd4s1 U7704 ( .DIN1(n6885), .DIN2(n6886), .DIN3(n6887), .DIN4(n6888), 
        .Q(n6884) );
  nnd2s1 U7705 ( .DIN1(n6889), .DIN2(n6890), .Q(n6888) );
  nnd2s1 U7706 ( .DIN1(n6030), .DIN2(n6891), .Q(n6890) );
  nnd2s1 U7707 ( .DIN1(n6892), .DIN2(n5553), .Q(n6891) );
  nnd2s1 U7708 ( .DIN1(n6893), .DIN2(n6894), .Q(n6892) );
  nnd2s1 U7709 ( .DIN1(n6168), .DIN2(n6895), .Q(n6889) );
  nnd2s1 U7710 ( .DIN1(n5322), .DIN2(n6034), .Q(n6895) );
  and2s1 U7711 ( .DIN1(n6035), .DIN2(n6896), .Q(n5322) );
  nnd2s1 U7712 ( .DIN1(n6035), .DIN2(n6897), .Q(n6168) );
  nnd2s1 U7713 ( .DIN1(n6898), .DIN2(n6899), .Q(n6897) );
  nnd2s1 U7714 ( .DIN1(n5321), .DIN2(n6896), .Q(n6899) );
  nnd2s1 U7715 ( .DIN1(n6900), .DIN2(n6901), .Q(n6887) );
  nnd4s1 U7716 ( .DIN1(n6902), .DIN2(n6903), .DIN3(n6904), .DIN4(n6905), 
        .Q(n6901) );
  nor2s1 U7717 ( .DIN1(n6906), .DIN2(n805), .Q(n6905) );
  and2s1 U7718 ( .DIN1(n5586), .DIN2(n554), .Q(n6906) );
  nnd4s1 U7719 ( .DIN1(n6907), .DIN2(n6908), .DIN3(n6909), .DIN4(n6910), 
        .Q(n5586) );
  nnd2s1 U7720 ( .DIN1(n545), .DIN2(n6044), .Q(n6904) );
  nnd2s1 U7721 ( .DIN1(n5824), .DIN2(n6911), .Q(n6903) );
  nnd2s1 U7722 ( .DIN1(n5826), .DIN2(n6479), .Q(n6902) );
  nnd2s1 U7723 ( .DIN1(n5547), .DIN2(n6912), .Q(n6900) );
  nnd2s1 U7724 ( .DIN1(n6913), .DIN2(n5301), .Q(n6912) );
  hi1s1 U7725 ( .DIN(n6914), .Q(n5301) );
  nnd2s1 U7726 ( .DIN1(n5570), .DIN2(n6915), .Q(n6886) );
  hi1s1 U7727 ( .DIN(n5558), .Q(n5570) );
  nnd2s1 U7728 ( .DIN1(n782), .DIN2(n6916), .Q(n6885) );
  nnd4s1 U7729 ( .DIN1(n6917), .DIN2(n6918), .DIN3(n6919), .DIN4(n6920), 
        .Q(n6916) );
  and4s1 U7730 ( .DIN1(n6921), .DIN2(n6922), .DIN3(n6923), .DIN4(n6924), 
        .Q(n6920) );
  nnd2s1 U7731 ( .DIN1(n6925), .DIN2(n6926), .Q(n6924) );
  nnd3s1 U7732 ( .DIN1(n6927), .DIN2(n749), .DIN3(n6928), .Q(n6925) );
  nnd2s1 U7733 ( .DIN1(n705), .DIN2(n6855), .Q(n6928) );
  nnd2s1 U7734 ( .DIN1(n654), .DIN2(n6851), .Q(n6927) );
  hi1s1 U7735 ( .DIN(n6852), .Q(n6851) );
  nnd2s1 U7736 ( .DIN1(n6929), .DIN2(n6930), .Q(n6923) );
  nnd2s1 U7737 ( .DIN1(n6931), .DIN2(n6932), .Q(n6930) );
  nnd2s1 U7738 ( .DIN1(n653), .DIN2(n6852), .Q(n6932) );
  nnd2s1 U7739 ( .DIN1(n6933), .DIN2(n6934), .Q(n6852) );
  nnd2s1 U7740 ( .DIN1(reg_out_B[16]), .DIN2(n6935), .Q(n6934) );
  nnd2s1 U7741 ( .DIN1(n6936), .DIN2(n71), .Q(n6935) );
  nnd2s1 U7742 ( .DIN1(n417), .DIN2(n6937), .Q(n6933) );
  or2s1 U7743 ( .DIN1(n6855), .DIN2(n706), .Q(n6931) );
  nnd2s1 U7744 ( .DIN1(n6938), .DIN2(n6939), .Q(n6855) );
  nnd2s1 U7745 ( .DIN1(n6940), .DIN2(n6941), .Q(n6939) );
  nnd2s1 U7746 ( .DIN1(n5468), .DIN2(n6942), .Q(n6922) );
  nnd2s1 U7747 ( .DIN1(n416), .DIN2(n767), .Q(n6921) );
  nnd2s1 U7748 ( .DIN1(reg_out_B[17]), .DIN2(n6943), .Q(n6919) );
  nnd2s1 U7749 ( .DIN1(n5471), .DIN2(n6944), .Q(n6943) );
  nnd2s1 U7750 ( .DIN1(n776), .DIN2(n416), .Q(n6944) );
  nnd3s1 U7751 ( .DIN1(n6945), .DIN2(n6946), .DIN3(n5336), .Q(n6918) );
  nnd2s1 U7752 ( .DIN1(n6433), .DIN2(n6947), .Q(n6946) );
  nnd2s1 U7753 ( .DIN1(n6948), .DIN2(n5478), .Q(n6947) );
  nnd2s1 U7754 ( .DIN1(n6436), .DIN2(n6949), .Q(n6945) );
  nnd2s1 U7755 ( .DIN1(n6087), .DIN2(n204), .Q(n6949) );
  nor2s1 U7756 ( .DIN1(n5337), .DIN2(n5366), .Q(n6436) );
  nor2s1 U7757 ( .DIN1(n6301), .DIN2(n753), .Q(n5366) );
  nnd2s1 U7758 ( .DIN1(n6950), .DIN2(n6951), .Q(n6917) );
  nnd4s1 U7759 ( .DIN1(n6952), .DIN2(n6953), .DIN3(n6954), .DIN4(n6955), 
        .Q(n6951) );
  nnd2s1 U7760 ( .DIN1(n546), .DIN2(n6524), .Q(n6955) );
  nor2s1 U7761 ( .DIN1(n752), .DIN2(n6956), .Q(n6954) );
  and2s1 U7762 ( .DIN1(n6957), .DIN2(n720), .Q(n6956) );
  nnd2s1 U7763 ( .DIN1(n621), .DIN2(n6095), .Q(n6953) );
  nnd2s1 U7764 ( .DIN1(n630), .DIN2(n5643), .Q(n6952) );
  nnd4s1 U7765 ( .DIN1(n6958), .DIN2(n6959), .DIN3(n6960), .DIN4(n6961), 
        .Q(n5643) );
  nnd2s1 U7766 ( .DIN1(n5342), .DIN2(n6962), .Q(n6950) );
  nnd2s1 U7767 ( .DIN1(n6963), .DIN2(n387), .Q(n6962) );
  nnd3s1 U7768 ( .DIN1(n6964), .DIN2(n6965), .DIN3(n6966), .Q(n6883) );
  nnd2s1 U7769 ( .DIN1(n727), .DIN2(\DM_addr[17] ), .Q(n6966) );
  nnd2s1 U7770 ( .DIN1(n416), .DIN2(n6967), .Q(n6965) );
  or3s1 U7771 ( .DIN1(n402), .DIN2(n6968), .DIN3(n6969), .Q(n6967) );
  nnd4s1 U7772 ( .DIN1(n6970), .DIN2(n6971), .DIN3(n6972), .DIN4(n6973), 
        .Q(n6969) );
  nnd2s1 U7773 ( .DIN1(n548), .DIN2(n6802), .Q(n6973) );
  nnd2s1 U7774 ( .DIN1(n5406), .DIN2(n6801), .Q(n6972) );
  nnd2s1 U7775 ( .DIN1(n5405), .DIN2(n13), .Q(n6971) );
  nnd2s1 U7776 ( .DIN1(n5665), .DIN2(n9474), .Q(n6970) );
  nor2s1 U7777 ( .DIN1(n5290), .DIN2(n6974), .Q(n6968) );
  nnd2s1 U7778 ( .DIN1(n6975), .DIN2(n82), .Q(n6964) );
  nnd4s1 U7779 ( .DIN1(n6976), .DIN2(n6977), .DIN3(n6978), .DIN4(n6979), 
        .Q(n6975) );
  nnd2s1 U7780 ( .DIN1(n5406), .DIN2(n6802), .Q(n6979) );
  nnd2s1 U7781 ( .DIN1(n549), .DIN2(n6801), .Q(n6978) );
  hi1s1 U7782 ( .DIN(n6802), .Q(n6801) );
  nnd2s1 U7783 ( .DIN1(n6980), .DIN2(n6981), .Q(n6802) );
  nnd2s1 U7784 ( .DIN1(n417), .DIN2(n6982), .Q(n6981) );
  nnd2s1 U7785 ( .DIN1(n6983), .DIN2(n5426), .Q(n6982) );
  nnd2s1 U7786 ( .DIN1(n633), .DIN2(n6984), .Q(n6980) );
  nnd2s1 U7787 ( .DIN1(n385), .DIN2(n6974), .Q(n6977) );
  xor2s1 U7788 ( .DIN1(n6796), .DIN2(n6797), .Q(n6974) );
  xor2s1 U7789 ( .DIN1(n13), .DIN2(n5413), .Q(n6797) );
  nnd2s1 U7790 ( .DIN1(n6985), .DIN2(n6986), .Q(n6796) );
  nnd2s1 U7791 ( .DIN1(n417), .DIN2(n6987), .Q(n6986) );
  nnd2s1 U7792 ( .DIN1(n6988), .DIN2(n6989), .Q(n6987) );
  or2s1 U7793 ( .DIN1(n6989), .DIN2(n6988), .Q(n6985) );
  nnd2s1 U7794 ( .DIN1(n5665), .DIN2(n13), .Q(n6976) );
  nor2s1 U7795 ( .DIN1(n9474), .DIN2(n5427), .Q(n6882) );
  nor2s1 U7796 ( .DIN1(n712), .DIN2(n5428), .Q(n6881) );
  nnd4s1 U7797 ( .DIN1(n6990), .DIN2(n6991), .DIN3(n6992), .DIN4(n6993), 
        .Q(\EXinst/n1448 ) );
  and4s1 U7798 ( .DIN1(n6994), .DIN2(n6995), .DIN3(n6996), .DIN4(n6997), 
        .Q(n6993) );
  nor2s1 U7799 ( .DIN1(n6998), .DIN2(n6999), .Q(n6997) );
  nor2s1 U7800 ( .DIN1(n9489), .DIN2(n5428), .Q(n6999) );
  nnd3s1 U7801 ( .DIN1(n7000), .DIN2(n9453), .DIN3(n7001), .Q(n5428) );
  nor2s1 U7802 ( .DIN1(n7002), .DIN2(n5558), .Q(n6998) );
  nnd2s1 U7803 ( .DIN1(n7003), .DIN2(n7004), .Q(n5558) );
  or2s1 U7804 ( .DIN1(n7005), .DIN2(n5288), .Q(n6996) );
  hi1s1 U7805 ( .DIN(n5665), .Q(n5288) );
  nor2s1 U7806 ( .DIN1(n7006), .DIN2(n48), .Q(n5665) );
  nnd3s1 U7807 ( .DIN1(n7007), .DIN2(n7008), .DIN3(n6035), .Q(n6995) );
  nnd2s1 U7808 ( .DIN1(n6030), .DIN2(n7009), .Q(n7008) );
  nnd2s1 U7809 ( .DIN1(n7010), .DIN2(n5553), .Q(n7009) );
  hi1s1 U7810 ( .DIN(n5808), .Q(n6030) );
  nnd2s1 U7811 ( .DIN1(n733), .DIN2(n7011), .Q(n5808) );
  nnd2s1 U7812 ( .DIN1(n5553), .DIN2(n805), .Q(n7011) );
  hi1s1 U7813 ( .DIN(n7012), .Q(n5553) );
  nnd2s1 U7814 ( .DIN1(n7013), .DIN2(n7014), .Q(n6994) );
  nnd4s1 U7815 ( .DIN1(n7015), .DIN2(n7016), .DIN3(n7017), .DIN4(n7018), 
        .Q(n7014) );
  nor2s1 U7816 ( .DIN1(n7019), .DIN2(n206), .Q(n7018) );
  and2s1 U7817 ( .DIN1(n5723), .DIN2(n555), .Q(n7019) );
  nnd4s1 U7818 ( .DIN1(n7020), .DIN2(n7021), .DIN3(n7022), .DIN4(n7023), 
        .Q(n5723) );
  nnd2s1 U7819 ( .DIN1(n544), .DIN2(n6176), .Q(n7017) );
  nnd2s1 U7820 ( .DIN1(n5824), .DIN2(n7024), .Q(n7016) );
  nnd2s1 U7821 ( .DIN1(n5826), .DIN2(n6608), .Q(n7015) );
  nnd2s1 U7822 ( .DIN1(n5547), .DIN2(n7025), .Q(n7013) );
  nnd2s1 U7823 ( .DIN1(n6688), .DIN2(n7026), .Q(n7025) );
  nor2s1 U7824 ( .DIN1(n6914), .DIN2(n6253), .Q(n6688) );
  nnd2s1 U7825 ( .DIN1(n7027), .DIN2(n6036), .Q(n6914) );
  and3s1 U7826 ( .DIN1(n7028), .DIN2(n7029), .DIN3(n7030), .Q(n6992) );
  nnd2s1 U7827 ( .DIN1(n5394), .DIN2(\DM_addr[16] ), .Q(n7030) );
  nnd2s1 U7828 ( .DIN1(n417), .DIN2(n7031), .Q(n7029) );
  nnd4s1 U7829 ( .DIN1(n7032), .DIN2(n7033), .DIN3(n7034), .DIN4(n5427), 
        .Q(n7031) );
  hi1s1 U7830 ( .DIN(n403), .Q(n5427) );
  nnd2s1 U7831 ( .DIN1(n7035), .DIN2(n385), .Q(n7034) );
  xnr2s1 U7832 ( .DIN1(n6989), .DIN2(n6988), .Q(n7035) );
  hi1s1 U7833 ( .DIN(n7036), .Q(n6988) );
  nnd2s1 U7834 ( .DIN1(n5405), .DIN2(n109), .Q(n7033) );
  nor2s1 U7835 ( .DIN1(n7037), .DIN2(n48), .Q(n5405) );
  nor2s1 U7836 ( .DIN1(n7038), .DIN2(n7039), .Q(n7032) );
  nor2s1 U7837 ( .DIN1(n6984), .DIN2(n7040), .Q(n7039) );
  nor2s1 U7838 ( .DIN1(n6983), .DIN2(n7041), .Q(n7038) );
  nnd2s1 U7839 ( .DIN1(n7042), .DIN2(n71), .Q(n7028) );
  nnd3s1 U7840 ( .DIN1(n7043), .DIN2(n7044), .DIN3(n7045), .Q(n7042) );
  nnd2s1 U7841 ( .DIN1(n385), .DIN2(n7046), .Q(n7045) );
  xnr2s1 U7842 ( .DIN1(n7036), .DIN2(n6989), .Q(n7046) );
  xor2s1 U7843 ( .DIN1(n9475), .DIN2(n745), .Q(n6989) );
  nnd2s1 U7844 ( .DIN1(n7047), .DIN2(n7048), .Q(n7036) );
  nnd2s1 U7845 ( .DIN1(n418), .DIN2(n7049), .Q(n7048) );
  or2s1 U7846 ( .DIN1(n7050), .DIN2(n7051), .Q(n7049) );
  nnd2s1 U7847 ( .DIN1(n7051), .DIN2(n7050), .Q(n7047) );
  nnd2s1 U7848 ( .DIN1(n5406), .DIN2(n6984), .Q(n7044) );
  hi1s1 U7849 ( .DIN(n7040), .Q(n5406) );
  nnd2s1 U7850 ( .DIN1(n7052), .DIN2(n5426), .Q(n7040) );
  nnd2s1 U7851 ( .DIN1(n548), .DIN2(n6983), .Q(n7043) );
  hi1s1 U7852 ( .DIN(n6984), .Q(n6983) );
  nnd2s1 U7853 ( .DIN1(n7053), .DIN2(n7054), .Q(n6984) );
  nnd2s1 U7854 ( .DIN1(n418), .DIN2(n7055), .Q(n7054) );
  or2s1 U7855 ( .DIN1(n7056), .DIN2(n7057), .Q(n7055) );
  nnd2s1 U7856 ( .DIN1(n7057), .DIN2(n7056), .Q(n7053) );
  nnd2s1 U7857 ( .DIN1(n5423), .DIN2(n7052), .Q(n7041) );
  and2s1 U7858 ( .DIN1(n550), .DIN2(n7058), .Q(n7052) );
  nnd2s1 U7859 ( .DIN1(n404), .DIN2(n109), .Q(n6991) );
  nnd2s1 U7860 ( .DIN1(n782), .DIN2(n7060), .Q(n6990) );
  nnd4s1 U7861 ( .DIN1(n7061), .DIN2(n7062), .DIN3(n7063), .DIN4(n7064), 
        .Q(n7060) );
  and4s1 U7862 ( .DIN1(n7065), .DIN2(n7066), .DIN3(n7067), .DIN4(n7068), 
        .Q(n7064) );
  nnd2s1 U7863 ( .DIN1(n7069), .DIN2(n7070), .Q(n7068) );
  nnd3s1 U7864 ( .DIN1(n7071), .DIN2(n5372), .DIN3(n7072), .Q(n7069) );
  nnd2s1 U7865 ( .DIN1(n620), .DIN2(n6941), .Q(n7072) );
  nnd2s1 U7866 ( .DIN1(n656), .DIN2(n6936), .Q(n7071) );
  hi1s1 U7867 ( .DIN(n6937), .Q(n6936) );
  nnd2s1 U7868 ( .DIN1(n7073), .DIN2(n7074), .Q(n7067) );
  nnd2s1 U7869 ( .DIN1(n7075), .DIN2(n7076), .Q(n7074) );
  nnd2s1 U7870 ( .DIN1(n655), .DIN2(n6937), .Q(n7076) );
  nnd2s1 U7871 ( .DIN1(n7077), .DIN2(n7078), .Q(n6937) );
  nnd2s1 U7872 ( .DIN1(reg_out_B[15]), .DIN2(n7079), .Q(n7078) );
  nnd2s1 U7873 ( .DIN1(n7080), .DIN2(n85), .Q(n7079) );
  nnd2s1 U7874 ( .DIN1(n418), .DIN2(n7081), .Q(n7077) );
  or2s1 U7875 ( .DIN1(n6941), .DIN2(n706), .Q(n7075) );
  nnd2s1 U7876 ( .DIN1(n7082), .DIN2(n7083), .Q(n6941) );
  nnd2s1 U7877 ( .DIN1(n7084), .DIN2(n7085), .Q(n7083) );
  nnd2s1 U7878 ( .DIN1(n5468), .DIN2(n7086), .Q(n7066) );
  hi1s1 U7879 ( .DIN(n5994), .Q(n5468) );
  nnd2s1 U7880 ( .DIN1(n417), .DIN2(n768), .Q(n7065) );
  nnd2s1 U7881 ( .DIN1(reg_out_B[16]), .DIN2(n7087), .Q(n7063) );
  nnd2s1 U7882 ( .DIN1(n5471), .DIN2(n7088), .Q(n7087) );
  nnd2s1 U7883 ( .DIN1(n775), .DIN2(n417), .Q(n7088) );
  nnd3s1 U7884 ( .DIN1(n7089), .DIN2(n7090), .DIN3(n769), .Q(n7062) );
  nnd2s1 U7885 ( .DIN1(n6433), .DIN2(n7091), .Q(n7090) );
  nnd2s1 U7886 ( .DIN1(n7086), .DIN2(n5478), .Q(n7091) );
  hi1s1 U7887 ( .DIN(n5865), .Q(n6433) );
  nnd2s1 U7888 ( .DIN1(n5337), .DIN2(n7092), .Q(n5865) );
  nnd2s1 U7889 ( .DIN1(n753), .DIN2(n5478), .Q(n7092) );
  nnd2s1 U7890 ( .DIN1(n7093), .DIN2(n7094), .Q(n7061) );
  nnd4s1 U7891 ( .DIN1(n7095), .DIN2(n7096), .DIN3(n7097), .DIN4(n7098), 
        .Q(n7094) );
  nnd2s1 U7892 ( .DIN1(n547), .DIN2(n6652), .Q(n7098) );
  nor2s1 U7893 ( .DIN1(n753), .DIN2(n7099), .Q(n7097) );
  and2s1 U7894 ( .DIN1(n7100), .DIN2(n720), .Q(n7099) );
  nnd2s1 U7895 ( .DIN1(n623), .DIN2(n6224), .Q(n7096) );
  nnd2s1 U7896 ( .DIN1(n629), .DIN2(n5791), .Q(n7095) );
  nnd4s1 U7897 ( .DIN1(n7101), .DIN2(n7102), .DIN3(n7103), .DIN4(n7104), 
        .Q(n5791) );
  nnd2s1 U7898 ( .DIN1(n5342), .DIN2(n7105), .Q(n7093) );
  nnd2s1 U7899 ( .DIN1(n6744), .DIN2(n7106), .Q(n7105) );
  and2s1 U7900 ( .DIN1(n387), .DIN2(n630), .Q(n6744) );
  nnd3s1 U7901 ( .DIN1(n7109), .DIN2(n7110), .DIN3(n7111), .Q(\EXinst/n1447 )
         );
  nnd2s1 U7902 ( .DIN1(n727), .DIN2(\DM_addr[15] ), .Q(n7111) );
  nnd2s1 U7903 ( .DIN1(n782), .DIN2(n7112), .Q(n7110) );
  nnd4s1 U7904 ( .DIN1(n7113), .DIN2(n7114), .DIN3(n7115), .DIN4(n7116), 
        .Q(n7112) );
  and4s1 U7905 ( .DIN1(n7117), .DIN2(n7118), .DIN3(n7119), .DIN4(n7120), 
        .Q(n7116) );
  nnd2s1 U7906 ( .DIN1(n7121), .DIN2(n7122), .Q(n7120) );
  nnd3s1 U7907 ( .DIN1(n7123), .DIN2(n749), .DIN3(n7124), .Q(n7121) );
  nnd2s1 U7908 ( .DIN1(n705), .DIN2(n7084), .Q(n7124) );
  nnd2s1 U7909 ( .DIN1(n654), .DIN2(n7080), .Q(n7123) );
  hi1s1 U7910 ( .DIN(n7081), .Q(n7080) );
  nnd2s1 U7911 ( .DIN1(n7125), .DIN2(n7126), .Q(n7119) );
  nnd2s1 U7912 ( .DIN1(n7127), .DIN2(n7128), .Q(n7126) );
  nnd2s1 U7913 ( .DIN1(n653), .DIN2(n7081), .Q(n7128) );
  nnd2s1 U7914 ( .DIN1(n7129), .DIN2(n7130), .Q(n7081) );
  nnd2s1 U7915 ( .DIN1(reg_out_B[14]), .DIN2(n7131), .Q(n7130) );
  nnd2s1 U7916 ( .DIN1(n7132), .DIN2(n31), .Q(n7131) );
  nnd2s1 U7917 ( .DIN1(n419), .DIN2(n7133), .Q(n7129) );
  or2s1 U7918 ( .DIN1(n7084), .DIN2(n5375), .Q(n7127) );
  nnd2s1 U7919 ( .DIN1(n7134), .DIN2(n7135), .Q(n7084) );
  nnd2s1 U7920 ( .DIN1(n7136), .DIN2(n7137), .Q(n7135) );
  nnd2s1 U7921 ( .DIN1(n7138), .DIN2(n5344), .Q(n7118) );
  nnd4s1 U7922 ( .DIN1(n7139), .DIN2(n7140), .DIN3(n7141), .DIN4(n7142), 
        .Q(n5344) );
  nnd2s1 U7923 ( .DIN1(n720), .DIN2(n6745), .Q(n7142) );
  nnd2s1 U7924 ( .DIN1(n546), .DIN2(n7143), .Q(n7141) );
  nnd2s1 U7925 ( .DIN1(n622), .DIN2(n6309), .Q(n7140) );
  nnd2s1 U7926 ( .DIN1(n630), .DIN2(n5875), .Q(n7139) );
  nnd4s1 U7927 ( .DIN1(n7144), .DIN2(n7145), .DIN3(n7146), .DIN4(n7147), 
        .Q(n5875) );
  nnd2s1 U7928 ( .DIN1(n418), .DIN2(n767), .Q(n7117) );
  nnd2s1 U7929 ( .DIN1(reg_out_B[15]), .DIN2(n7148), .Q(n7115) );
  nnd2s1 U7930 ( .DIN1(n5471), .DIN2(n7149), .Q(n7148) );
  nnd2s1 U7931 ( .DIN1(n776), .DIN2(n418), .Q(n7149) );
  nnd3s1 U7932 ( .DIN1(n7150), .DIN2(n7151), .DIN3(n5336), .Q(n7114) );
  nnd2s1 U7933 ( .DIN1(n5337), .DIN2(n7152), .Q(n7151) );
  nnd2s1 U7934 ( .DIN1(n7153), .DIN2(n5478), .Q(n7152) );
  nnd2s1 U7935 ( .DIN1(n55), .DIN2(n401), .Q(n5478) );
  nnd2s1 U7936 ( .DIN1(n7154), .DIN2(n7155), .Q(n7150) );
  nnd2s1 U7937 ( .DIN1(n5362), .DIN2(n7156), .Q(n7155) );
  nnd2s1 U7938 ( .DIN1(n7157), .DIN2(n7153), .Q(n7113) );
  nnd4s1 U7939 ( .DIN1(n7158), .DIN2(n7159), .DIN3(n7160), .DIN4(n7161), 
        .Q(n7153) );
  nnd2s1 U7940 ( .DIN1(n547), .DIN2(n6729), .Q(n7161) );
  nor2s1 U7941 ( .DIN1(n55), .DIN2(n7162), .Q(n7160) );
  nor2s1 U7942 ( .DIN1(n6299), .DIN2(n5359), .Q(n7162) );
  nnd2s1 U7943 ( .DIN1(n621), .DIN2(n6728), .Q(n7159) );
  nnd2s1 U7944 ( .DIN1(n629), .DIN2(n7163), .Q(n7158) );
  nnd2s1 U7945 ( .DIN1(n5994), .DIN2(n7164), .Q(n7157) );
  nnd2s1 U7946 ( .DIN1(n7165), .DIN2(n5362), .Q(n7164) );
  nnd2s1 U7947 ( .DIN1(n550), .DIN2(n7166), .Q(n7109) );
  nnd4s1 U7948 ( .DIN1(n7167), .DIN2(n7168), .DIN3(n7169), .DIN4(n7170), 
        .Q(n7166) );
  and3s1 U7949 ( .DIN1(n7171), .DIN2(n7172), .DIN3(n7173), .Q(n7170) );
  nnd2s1 U7950 ( .DIN1(n400), .DIN2(n5300), .Q(n7173) );
  nnd4s1 U7951 ( .DIN1(n7174), .DIN2(n7175), .DIN3(n7176), .DIN4(n7177), 
        .Q(n5300) );
  nnd2s1 U7952 ( .DIN1(n5824), .DIN2(n6689), .Q(n7177) );
  nnd2s1 U7953 ( .DIN1(n5826), .DIN2(n6686), .Q(n7176) );
  nnd2s1 U7954 ( .DIN1(n545), .DIN2(n6258), .Q(n7175) );
  nnd2s1 U7955 ( .DIN1(n554), .DIN2(n5825), .Q(n7174) );
  nnd4s1 U7956 ( .DIN1(n7178), .DIN2(n7179), .DIN3(n7180), .DIN4(n7181), 
        .Q(n5825) );
  nnd4s1 U7957 ( .DIN1(n7182), .DIN2(n7183), .DIN3(n7184), .DIN4(n7185), 
        .Q(n7172) );
  and3s1 U7958 ( .DIN1(n7186), .DIN2(n7187), .DIN3(n7188), .Q(n7185) );
  nnd2s1 U7959 ( .DIN1(n7189), .DIN2(n544), .Q(n7187) );
  nnd2s1 U7960 ( .DIN1(n7190), .DIN2(n806), .Q(n7186) );
  nnd2s1 U7961 ( .DIN1(n7191), .DIN2(n5824), .Q(n7183) );
  nnd2s1 U7962 ( .DIN1(n7192), .DIN2(n726), .Q(n7182) );
  nnd4s1 U7963 ( .DIN1(n7193), .DIN2(n7194), .DIN3(n7195), .DIN4(n7196), 
        .Q(n7171) );
  nnd2s1 U7964 ( .DIN1(n9486), .DIN2(n7197), .Q(n7195) );
  nnd4s1 U7965 ( .DIN1(n7184), .DIN2(n7198), .DIN3(n7199), .DIN4(n7200), 
        .Q(n7197) );
  nnd2s1 U7966 ( .DIN1(n7191), .DIN2(n719), .Q(n7200) );
  nor2s1 U7967 ( .DIN1(n7012), .DIN2(n7201), .Q(n7199) );
  nor2s1 U7968 ( .DIN1(n7202), .DIN2(n7203), .Q(n7201) );
  nor2s1 U7969 ( .DIN1(n734), .DIN2(n56), .Q(n7012) );
  nnd2s1 U7970 ( .DIN1(n7189), .DIN2(n397), .Q(n7198) );
  nnd2s1 U7971 ( .DIN1(n7204), .DIN2(n700), .Q(n7184) );
  nnd2s1 U7972 ( .DIN1(n7205), .DIN2(n7190), .Q(n7194) );
  nnd2s1 U7973 ( .DIN1(n7206), .DIN2(n7), .Q(n7169) );
  nnd2s1 U7974 ( .DIN1(n418), .DIN2(n7207), .Q(n7168) );
  nnd4s1 U7975 ( .DIN1(n7208), .DIN2(n7209), .DIN3(n7210), .DIN4(n7059), 
        .Q(n7207) );
  nnd2s1 U7976 ( .DIN1(n7211), .DIN2(n7212), .Q(n7210) );
  xnr2s1 U7977 ( .DIN1(n7050), .DIN2(n7051), .Q(n7211) );
  hi1s1 U7978 ( .DIN(n7213), .Q(n7051) );
  nnd2s1 U7979 ( .DIN1(n7214), .DIN2(n743), .Q(n7209) );
  xnr2s1 U7980 ( .DIN1(n7056), .DIN2(n7057), .Q(n7214) );
  hi1s1 U7981 ( .DIN(n7215), .Q(n7057) );
  nor2s1 U7982 ( .DIN1(n7216), .DIN2(n7217), .Q(n7208) );
  nor2s1 U7983 ( .DIN1(n7), .DIN2(n7006), .Q(n7217) );
  nor2s1 U7984 ( .DIN1(n9476), .DIN2(n7037), .Q(n7216) );
  nnd2s1 U7985 ( .DIN1(n7218), .DIN2(n85), .Q(n7167) );
  nnd3s1 U7986 ( .DIN1(n7219), .DIN2(n7220), .DIN3(n7221), .Q(n7218) );
  nnd2s1 U7987 ( .DIN1(n7222), .DIN2(n7), .Q(n7221) );
  nnd2s1 U7988 ( .DIN1(n7223), .DIN2(n722), .Q(n7220) );
  xnr2s1 U7989 ( .DIN1(n7050), .DIN2(n7213), .Q(n7223) );
  xnr2s1 U7990 ( .DIN1(n9476), .DIN2(n785), .Q(n7213) );
  nnd2s1 U7991 ( .DIN1(n7224), .DIN2(n7225), .Q(n7050) );
  nnd2s1 U7992 ( .DIN1(n419), .DIN2(n7226), .Q(n7225) );
  nnd2s1 U7993 ( .DIN1(n7227), .DIN2(n7228), .Q(n7226) );
  or2s1 U7994 ( .DIN1(n7228), .DIN2(n7227), .Q(n7224) );
  nnd2s1 U7995 ( .DIN1(n7229), .DIN2(n7058), .Q(n7219) );
  xnr2s1 U7996 ( .DIN1(n7056), .DIN2(n7215), .Q(n7229) );
  xnr2s1 U7997 ( .DIN1(n633), .DIN2(n7), .Q(n7215) );
  nnd2s1 U7998 ( .DIN1(n7230), .DIN2(n7231), .Q(n7056) );
  nnd2s1 U7999 ( .DIN1(n419), .DIN2(n7232), .Q(n7231) );
  nnd2s1 U8000 ( .DIN1(n7233), .DIN2(n388), .Q(n7232) );
  or2s1 U8001 ( .DIN1(n388), .DIN2(n7233), .Q(n7230) );
  nnd3s1 U8002 ( .DIN1(n7234), .DIN2(n7235), .DIN3(n7236), .Q(\EXinst/n1446 )
         );
  nnd2s1 U8003 ( .DIN1(n5394), .DIN2(\DM_addr[14] ), .Q(n7236) );
  nnd2s1 U8004 ( .DIN1(n5324), .DIN2(n7237), .Q(n7235) );
  nnd4s1 U8005 ( .DIN1(n7238), .DIN2(n7239), .DIN3(n7240), .DIN4(n7241), 
        .Q(n7237) );
  and4s1 U8006 ( .DIN1(n7242), .DIN2(n7243), .DIN3(n7244), .DIN4(n7245), 
        .Q(n7241) );
  nnd2s1 U8007 ( .DIN1(n7246), .DIN2(n7247), .Q(n7245) );
  nnd3s1 U8008 ( .DIN1(n7248), .DIN2(n5372), .DIN3(n7249), .Q(n7246) );
  nnd2s1 U8009 ( .DIN1(n620), .DIN2(n7137), .Q(n7249) );
  nnd2s1 U8010 ( .DIN1(n656), .DIN2(n7132), .Q(n7248) );
  hi1s1 U8011 ( .DIN(n7133), .Q(n7132) );
  nnd2s1 U8012 ( .DIN1(n7250), .DIN2(n7251), .Q(n7244) );
  nnd2s1 U8013 ( .DIN1(n7252), .DIN2(n7253), .Q(n7251) );
  nnd2s1 U8014 ( .DIN1(n655), .DIN2(n7133), .Q(n7253) );
  nnd2s1 U8015 ( .DIN1(n7254), .DIN2(n7255), .Q(n7133) );
  nnd2s1 U8016 ( .DIN1(reg_out_B[13]), .DIN2(n7256), .Q(n7255) );
  nnd2s1 U8017 ( .DIN1(n7257), .DIN2(n86), .Q(n7256) );
  nnd2s1 U8018 ( .DIN1(n420), .DIN2(n7258), .Q(n7254) );
  or2s1 U8019 ( .DIN1(n7137), .DIN2(n706), .Q(n7252) );
  nnd2s1 U8020 ( .DIN1(n7259), .DIN2(n7260), .Q(n7137) );
  nnd2s1 U8021 ( .DIN1(n7261), .DIN2(n7262), .Q(n7260) );
  nnd2s1 U8022 ( .DIN1(n7138), .DIN2(n5502), .Q(n7243) );
  nnd4s1 U8023 ( .DIN1(n7263), .DIN2(n7264), .DIN3(n7265), .DIN4(n7266), 
        .Q(n5502) );
  nnd2s1 U8024 ( .DIN1(n720), .DIN2(n6879), .Q(n7266) );
  nnd2s1 U8025 ( .DIN1(n546), .DIN2(n7267), .Q(n7265) );
  nnd2s1 U8026 ( .DIN1(n623), .DIN2(n6445), .Q(n7264) );
  nnd2s1 U8027 ( .DIN1(n630), .DIN2(n6011), .Q(n7263) );
  nnd4s1 U8028 ( .DIN1(n7268), .DIN2(n7269), .DIN3(n7270), .DIN4(n7271), 
        .Q(n6011) );
  nnd2s1 U8029 ( .DIN1(n419), .DIN2(n768), .Q(n7242) );
  nnd2s1 U8030 ( .DIN1(reg_out_B[14]), .DIN2(n7272), .Q(n7240) );
  nnd2s1 U8031 ( .DIN1(n5471), .DIN2(n7273), .Q(n7272) );
  nnd2s1 U8032 ( .DIN1(n775), .DIN2(n419), .Q(n7273) );
  nnd3s1 U8033 ( .DIN1(n7274), .DIN2(n7275), .DIN3(n769), .Q(n7239) );
  nnd4s1 U8034 ( .DIN1(n7276), .DIN2(n7277), .DIN3(n7278), .DIN4(n7279), 
        .Q(n7275) );
  nnd2s1 U8035 ( .DIN1(n7280), .DIN2(n808), .Q(n7279) );
  nnd3s1 U8036 ( .DIN1(n5477), .DIN2(n801), .DIN3(n752), .Q(n7278) );
  nnd2s1 U8037 ( .DIN1(n5345), .DIN2(n7281), .Q(n7277) );
  nnd2s1 U8038 ( .DIN1(n7154), .DIN2(n7282), .Q(n7274) );
  nnd3s1 U8039 ( .DIN1(n714), .DIN2(n337), .DIN3(n7283), .Q(n7282) );
  nnd2s1 U8040 ( .DIN1(n7284), .DIN2(n7285), .Q(n7238) );
  nnd3s1 U8041 ( .DIN1(n7286), .DIN2(n808), .DIN3(n7287), .Q(n7285) );
  hi1s1 U8042 ( .DIN(n7280), .Q(n7287) );
  nnd3s1 U8043 ( .DIN1(n7288), .DIN2(n7289), .DIN3(n7290), .Q(n7280) );
  nnd2s1 U8044 ( .DIN1(n622), .DIN2(n7291), .Q(n7290) );
  nnd2s1 U8045 ( .DIN1(n720), .DIN2(n7292), .Q(n7289) );
  nnd2s1 U8046 ( .DIN1(n547), .DIN2(n7293), .Q(n7288) );
  nnd2s1 U8047 ( .DIN1(n629), .DIN2(n7281), .Q(n7286) );
  nnd2s1 U8048 ( .DIN1(n5994), .DIN2(n7294), .Q(n7284) );
  nnd2s1 U8049 ( .DIN1(n386), .DIN2(n5467), .Q(n7294) );
  and4s1 U8050 ( .DIN1(n630), .DIN2(n714), .DIN3(n7295), .DIN4(n7296), 
        .Q(n5467) );
  nnd2s1 U8051 ( .DIN1(n399), .DIN2(n62), .Q(n7296) );
  nnd2s1 U8052 ( .DIN1(n717), .DIN2(n1), .Q(n7295) );
  nnd2s1 U8053 ( .DIN1(n9453), .DIN2(n7297), .Q(n7234) );
  nnd4s1 U8054 ( .DIN1(n7298), .DIN2(n7299), .DIN3(n7300), .DIN4(n7301), 
        .Q(n7297) );
  and4s1 U8055 ( .DIN1(n7302), .DIN2(n7303), .DIN3(n7304), .DIN4(n7305), 
        .Q(n7301) );
  nnd2s1 U8056 ( .DIN1(n419), .DIN2(n7306), .Q(n7305) );
  nnd4s1 U8057 ( .DIN1(n7307), .DIN2(n7308), .DIN3(n7309), .DIN4(n7059), 
        .Q(n7306) );
  nnd2s1 U8058 ( .DIN1(n7310), .DIN2(n7212), .Q(n7309) );
  xnr2s1 U8059 ( .DIN1(n7228), .DIN2(n7227), .Q(n7310) );
  hi1s1 U8060 ( .DIN(n7311), .Q(n7227) );
  nnd2s1 U8061 ( .DIN1(n7312), .DIN2(n743), .Q(n7308) );
  xnr2s1 U8062 ( .DIN1(n388), .DIN2(n7233), .Q(n7312) );
  hi1s1 U8063 ( .DIN(n7313), .Q(n7233) );
  nnd2s1 U8064 ( .DIN1(n7314), .DIN2(n108), .Q(n7307) );
  nnd2s1 U8065 ( .DIN1(n7315), .DIN2(n31), .Q(n7304) );
  nnd2s1 U8066 ( .DIN1(n7316), .DIN2(n7317), .Q(n7315) );
  nnd2s1 U8067 ( .DIN1(n7318), .DIN2(n722), .Q(n7317) );
  xnr2s1 U8068 ( .DIN1(n7311), .DIN2(n7228), .Q(n7318) );
  xor2s1 U8069 ( .DIN1(n9477), .DIN2(n5413), .Q(n7228) );
  nnd2s1 U8070 ( .DIN1(n7319), .DIN2(n7320), .Q(n7311) );
  nnd2s1 U8071 ( .DIN1(n420), .DIN2(n7321), .Q(n7320) );
  or2s1 U8072 ( .DIN1(n7322), .DIN2(n7323), .Q(n7321) );
  nnd2s1 U8073 ( .DIN1(n7323), .DIN2(n7322), .Q(n7319) );
  nnd2s1 U8074 ( .DIN1(n7324), .DIN2(n7058), .Q(n7316) );
  xnr2s1 U8075 ( .DIN1(n7313), .DIN2(n388), .Q(n7324) );
  nnd2s1 U8076 ( .DIN1(n7325), .DIN2(n7326), .Q(n7313) );
  nnd2s1 U8077 ( .DIN1(n420), .DIN2(n7327), .Q(n7326) );
  or2s1 U8078 ( .DIN1(n7328), .DIN2(n7329), .Q(n7327) );
  nnd2s1 U8079 ( .DIN1(n7329), .DIN2(n7328), .Q(n7325) );
  nnd2s1 U8080 ( .DIN1(n400), .DIN2(n5549), .Q(n7303) );
  nnd4s1 U8081 ( .DIN1(n7330), .DIN2(n7331), .DIN3(n7332), .DIN4(n7333), 
        .Q(n5549) );
  nnd2s1 U8082 ( .DIN1(n5824), .DIN2(n6830), .Q(n7333) );
  nnd2s1 U8083 ( .DIN1(n5826), .DIN2(n6828), .Q(n7332) );
  nnd2s1 U8084 ( .DIN1(n544), .DIN2(n6399), .Q(n7331) );
  nnd2s1 U8085 ( .DIN1(n555), .DIN2(n5959), .Q(n7330) );
  nnd4s1 U8086 ( .DIN1(n7334), .DIN2(n7335), .DIN3(n7336), .DIN4(n7337), 
        .Q(n5959) );
  nnd2s1 U8087 ( .DIN1(n7206), .DIN2(n108), .Q(n7302) );
  or2s1 U8088 ( .DIN1(n7338), .DIN2(n7006), .Q(n7300) );
  nnd3s1 U8089 ( .DIN1(n730), .DIN2(n7340), .DIN3(n7341), .Q(n7299) );
  hi1s1 U8090 ( .DIN(n7342), .Q(n7341) );
  nnd2s1 U8091 ( .DIN1(n5559), .DIN2(n805), .Q(n7340) );
  nnd3s1 U8092 ( .DIN1(n7343), .DIN2(n7344), .DIN3(n7345), .Q(n5559) );
  nnd2s1 U8093 ( .DIN1(n9489), .DIN2(n717), .Q(n7344) );
  nnd2s1 U8094 ( .DIN1(n440), .DIN2(n401), .Q(n7343) );
  nnd4s1 U8095 ( .DIN1(n7346), .DIN2(n7347), .DIN3(n7348), .DIN4(n7349), 
        .Q(n7298) );
  nnd2s1 U8096 ( .DIN1(n7350), .DIN2(n6387), .Q(n7349) );
  hi1s1 U8097 ( .DIN(n5557), .Q(n6387) );
  or2s1 U8098 ( .DIN1(n6380), .DIN2(n7345), .Q(n7348) );
  nnd2s1 U8099 ( .DIN1(n9486), .DIN2(n7342), .Q(n7347) );
  nnd4s1 U8100 ( .DIN1(n7351), .DIN2(n7352), .DIN3(n7353), .DIN4(n7354), 
        .Q(n7342) );
  nnd2s1 U8101 ( .DIN1(n6386), .DIN2(n763), .Q(n7354) );
  nnd2s1 U8102 ( .DIN1(n6385), .DIN2(n5304), .Q(n7353) );
  hi1s1 U8103 ( .DIN(n7355), .Q(n6385) );
  nnd2s1 U8104 ( .DIN1(n7356), .DIN2(n398), .Q(n7352) );
  nnd2s1 U8105 ( .DIN1(n7357), .DIN2(n700), .Q(n7351) );
  nnd3s1 U8106 ( .DIN1(n7358), .DIN2(n7359), .DIN3(n7360), .Q(\EXinst/n1445 )
         );
  nnd2s1 U8107 ( .DIN1(n727), .DIN2(\DM_addr[13] ), .Q(n7360) );
  nnd2s1 U8108 ( .DIN1(n5324), .DIN2(n7361), .Q(n7359) );
  nnd4s1 U8109 ( .DIN1(n7362), .DIN2(n7363), .DIN3(n7364), .DIN4(n7365), 
        .Q(n7361) );
  and4s1 U8110 ( .DIN1(n7366), .DIN2(n7367), .DIN3(n7368), .DIN4(n7369), 
        .Q(n7365) );
  nnd2s1 U8111 ( .DIN1(n7370), .DIN2(n7371), .Q(n7369) );
  nnd3s1 U8112 ( .DIN1(n7372), .DIN2(n749), .DIN3(n7373), .Q(n7370) );
  nnd2s1 U8113 ( .DIN1(n705), .DIN2(n7261), .Q(n7373) );
  nnd2s1 U8114 ( .DIN1(n654), .DIN2(n7257), .Q(n7372) );
  hi1s1 U8115 ( .DIN(n7258), .Q(n7257) );
  nnd2s1 U8116 ( .DIN1(n7374), .DIN2(n7375), .Q(n7368) );
  nnd2s1 U8117 ( .DIN1(n7376), .DIN2(n7377), .Q(n7375) );
  nnd2s1 U8118 ( .DIN1(n653), .DIN2(n7258), .Q(n7377) );
  nnd2s1 U8119 ( .DIN1(n7378), .DIN2(n7379), .Q(n7258) );
  nnd2s1 U8120 ( .DIN1(reg_out_B[12]), .DIN2(n7380), .Q(n7379) );
  nnd2s1 U8121 ( .DIN1(n7381), .DIN2(n64), .Q(n7380) );
  nnd2s1 U8122 ( .DIN1(n421), .DIN2(n7382), .Q(n7378) );
  or2s1 U8123 ( .DIN1(n7261), .DIN2(n706), .Q(n7376) );
  nnd2s1 U8124 ( .DIN1(n7383), .DIN2(n7384), .Q(n7261) );
  nnd2s1 U8125 ( .DIN1(n7385), .DIN2(n7386), .Q(n7384) );
  nnd2s1 U8126 ( .DIN1(n7138), .DIN2(n5646), .Q(n7367) );
  nnd3s1 U8127 ( .DIN1(n7387), .DIN2(n7388), .DIN3(n7389), .Q(n5646) );
  nnd2s1 U8128 ( .DIN1(n438), .DIN2(n6530), .Q(n7389) );
  nnd2s1 U8129 ( .DIN1(n621), .DIN2(n6524), .Q(n7388) );
  nnd2s1 U8130 ( .DIN1(n630), .DIN2(n6095), .Q(n7387) );
  nnd4s1 U8131 ( .DIN1(n7390), .DIN2(n7391), .DIN3(n7392), .DIN4(n7393), 
        .Q(n6095) );
  nnd2s1 U8132 ( .DIN1(n532), .DIN2(n423), .Q(n7392) );
  nnd2s1 U8133 ( .DIN1(n420), .DIN2(n767), .Q(n7366) );
  nnd2s1 U8134 ( .DIN1(reg_out_B[13]), .DIN2(n7394), .Q(n7364) );
  nnd2s1 U8135 ( .DIN1(n5471), .DIN2(n7395), .Q(n7394) );
  nnd2s1 U8136 ( .DIN1(n776), .DIN2(n420), .Q(n7395) );
  nnd3s1 U8137 ( .DIN1(n7396), .DIN2(n7397), .DIN3(n7398), .Q(n7363) );
  nnd4s1 U8138 ( .DIN1(n7399), .DIN2(n7400), .DIN3(n7401), .DIN4(n7402), 
        .Q(n7397) );
  nnd2s1 U8139 ( .DIN1(n7403), .DIN2(n204), .Q(n7402) );
  nnd3s1 U8140 ( .DIN1(n628), .DIN2(n5651), .DIN3(n753), .Q(n7401) );
  nnd2s1 U8141 ( .DIN1(n5345), .DIN2(n7404), .Q(n7400) );
  nnd2s1 U8142 ( .DIN1(n6723), .DIN2(n5653), .Q(n7396) );
  nnd3s1 U8143 ( .DIN1(n211), .DIN2(n801), .DIN3(n7283), .Q(n5653) );
  nnd2s1 U8144 ( .DIN1(n7405), .DIN2(n7406), .Q(n7362) );
  nnd3s1 U8145 ( .DIN1(n7407), .DIN2(n808), .DIN3(n7408), .Q(n7406) );
  hi1s1 U8146 ( .DIN(n7403), .Q(n7408) );
  nnd3s1 U8147 ( .DIN1(n7409), .DIN2(n7410), .DIN3(n7411), .Q(n7403) );
  nnd2s1 U8148 ( .DIN1(n623), .DIN2(n7412), .Q(n7411) );
  nnd2s1 U8149 ( .DIN1(n720), .DIN2(n7413), .Q(n7410) );
  nnd2s1 U8150 ( .DIN1(n546), .DIN2(n7414), .Q(n7409) );
  nnd2s1 U8151 ( .DIN1(n629), .DIN2(n7404), .Q(n7407) );
  nnd2s1 U8152 ( .DIN1(n5994), .DIN2(n7415), .Q(n7405) );
  nnd3s1 U8153 ( .DIN1(n628), .DIN2(n5654), .DIN3(n386), .Q(n7415) );
  nnd2s1 U8154 ( .DIN1(n551), .DIN2(n7416), .Q(n7358) );
  nnd4s1 U8155 ( .DIN1(n7417), .DIN2(n7418), .DIN3(n7419), .DIN4(n7420), 
        .Q(n7416) );
  and3s1 U8156 ( .DIN1(n7421), .DIN2(n7422), .DIN3(n7423), .Q(n7420) );
  nnd2s1 U8157 ( .DIN1(n400), .DIN2(n5598), .Q(n7423) );
  nnd3s1 U8158 ( .DIN1(n7424), .DIN2(n7425), .DIN3(n7426), .Q(n5598) );
  nnd2s1 U8159 ( .DIN1(n6481), .DIN2(n4840), .Q(n7426) );
  nnd2s1 U8160 ( .DIN1(n545), .DIN2(n6479), .Q(n7425) );
  nnd2s1 U8161 ( .DIN1(n554), .DIN2(n6044), .Q(n7424) );
  nnd4s1 U8162 ( .DIN1(n7427), .DIN2(n7428), .DIN3(n7429), .DIN4(n7430), 
        .Q(n6044) );
  nnd2s1 U8163 ( .DIN1(n759), .DIN2(n423), .Q(n7429) );
  nnd4s1 U8164 ( .DIN1(n7431), .DIN2(n7432), .DIN3(n7433), .DIN4(n7434), 
        .Q(n7422) );
  and3s1 U8165 ( .DIN1(n7435), .DIN2(n7436), .DIN3(n7437), .Q(n7434) );
  nnd2s1 U8166 ( .DIN1(n7438), .DIN2(n700), .Q(n7437) );
  nnd2s1 U8167 ( .DIN1(n7439), .DIN2(n5824), .Q(n7436) );
  nnd2s1 U8168 ( .DIN1(n7440), .DIN2(n726), .Q(n7435) );
  nnd2s1 U8169 ( .DIN1(n7441), .DIN2(n545), .Q(n7432) );
  nnd2s1 U8170 ( .DIN1(n7442), .DIN2(n806), .Q(n7431) );
  nnd3s1 U8171 ( .DIN1(n7443), .DIN2(n7444), .DIN3(n7193), .Q(n7421) );
  nnd4s1 U8172 ( .DIN1(n7445), .DIN2(n7446), .DIN3(n7447), .DIN4(n7448), 
        .Q(n7444) );
  and3s1 U8173 ( .DIN1(n7449), .DIN2(n7450), .DIN3(n7451), .Q(n7448) );
  nnd2s1 U8174 ( .DIN1(n5304), .DIN2(n7452), .Q(n7451) );
  nnd2s1 U8175 ( .DIN1(n7453), .DIN2(n5575), .Q(n7450) );
  nnd2s1 U8176 ( .DIN1(n5315), .DIN2(n7454), .Q(n7449) );
  nnd2s1 U8177 ( .DIN1(n397), .DIN2(n7455), .Q(n7446) );
  nnd2s1 U8178 ( .DIN1(n5306), .DIN2(n7456), .Q(n7445) );
  nnd2s1 U8179 ( .DIN1(n7205), .DIN2(n5578), .Q(n7443) );
  nnd3s1 U8180 ( .DIN1(n9487), .DIN2(n5313), .DIN3(n6465), .Q(n5578) );
  nnd2s1 U8181 ( .DIN1(n7206), .DIN2(n9), .Q(n7419) );
  nnd2s1 U8182 ( .DIN1(n420), .DIN2(n7457), .Q(n7418) );
  nnd4s1 U8183 ( .DIN1(n7458), .DIN2(n7459), .DIN3(n7460), .DIN4(n7059), 
        .Q(n7457) );
  nnd2s1 U8184 ( .DIN1(n7461), .DIN2(n7212), .Q(n7460) );
  xnr2s1 U8185 ( .DIN1(n7322), .DIN2(n7323), .Q(n7461) );
  hi1s1 U8186 ( .DIN(n7462), .Q(n7323) );
  nnd2s1 U8187 ( .DIN1(n7463), .DIN2(n743), .Q(n7459) );
  xnr2s1 U8188 ( .DIN1(n7328), .DIN2(n7329), .Q(n7463) );
  hi1s1 U8189 ( .DIN(n7464), .Q(n7329) );
  nor2s1 U8190 ( .DIN1(n7465), .DIN2(n7466), .Q(n7458) );
  nor2s1 U8191 ( .DIN1(n9), .DIN2(n7006), .Q(n7466) );
  nor2s1 U8192 ( .DIN1(n9478), .DIN2(n7037), .Q(n7465) );
  nnd2s1 U8193 ( .DIN1(n7467), .DIN2(n86), .Q(n7417) );
  nnd3s1 U8194 ( .DIN1(n7468), .DIN2(n7469), .DIN3(n7470), .Q(n7467) );
  nnd2s1 U8195 ( .DIN1(n7222), .DIN2(n9), .Q(n7470) );
  nnd2s1 U8196 ( .DIN1(n7471), .DIN2(n722), .Q(n7469) );
  xnr2s1 U8197 ( .DIN1(n7322), .DIN2(n7462), .Q(n7471) );
  xnr2s1 U8198 ( .DIN1(n9478), .DIN2(n788), .Q(n7462) );
  nnd2s1 U8199 ( .DIN1(n7472), .DIN2(n7473), .Q(n7322) );
  nnd2s1 U8200 ( .DIN1(n421), .DIN2(n7474), .Q(n7473) );
  nnd2s1 U8201 ( .DIN1(n7475), .DIN2(n7476), .Q(n7474) );
  or2s1 U8202 ( .DIN1(n7476), .DIN2(n7475), .Q(n7472) );
  nnd2s1 U8203 ( .DIN1(n7477), .DIN2(n7058), .Q(n7468) );
  xnr2s1 U8204 ( .DIN1(n7328), .DIN2(n7464), .Q(n7477) );
  xnr2s1 U8205 ( .DIN1(n5423), .DIN2(n9), .Q(n7464) );
  nnd2s1 U8206 ( .DIN1(n7478), .DIN2(n7479), .Q(n7328) );
  nnd2s1 U8207 ( .DIN1(n421), .DIN2(n7480), .Q(n7479) );
  nnd2s1 U8208 ( .DIN1(n7481), .DIN2(n389), .Q(n7480) );
  or2s1 U8209 ( .DIN1(n389), .DIN2(n7481), .Q(n7478) );
  nnd3s1 U8210 ( .DIN1(n7482), .DIN2(n7483), .DIN3(n7484), .Q(\EXinst/n1444 )
         );
  nnd2s1 U8211 ( .DIN1(n5394), .DIN2(\DM_addr[12] ), .Q(n7484) );
  nnd2s1 U8212 ( .DIN1(n5324), .DIN2(n7485), .Q(n7483) );
  nnd4s1 U8213 ( .DIN1(n7486), .DIN2(n7487), .DIN3(n7488), .DIN4(n7489), 
        .Q(n7485) );
  and4s1 U8214 ( .DIN1(n7490), .DIN2(n7491), .DIN3(n7492), .DIN4(n7493), 
        .Q(n7489) );
  nnd2s1 U8215 ( .DIN1(n7494), .DIN2(n7495), .Q(n7493) );
  nnd3s1 U8216 ( .DIN1(n7496), .DIN2(n5372), .DIN3(n7497), .Q(n7494) );
  nnd2s1 U8217 ( .DIN1(n620), .DIN2(n7386), .Q(n7497) );
  nnd2s1 U8218 ( .DIN1(n656), .DIN2(n7381), .Q(n7496) );
  hi1s1 U8219 ( .DIN(n7382), .Q(n7381) );
  nnd2s1 U8220 ( .DIN1(n7498), .DIN2(n7499), .Q(n7492) );
  nnd2s1 U8221 ( .DIN1(n7500), .DIN2(n7501), .Q(n7499) );
  nnd2s1 U8222 ( .DIN1(n655), .DIN2(n7382), .Q(n7501) );
  nnd2s1 U8223 ( .DIN1(n7502), .DIN2(n7503), .Q(n7382) );
  nnd2s1 U8224 ( .DIN1(reg_out_B[11]), .DIN2(n7504), .Q(n7503) );
  nnd2s1 U8225 ( .DIN1(n7505), .DIN2(n84), .Q(n7504) );
  nnd2s1 U8226 ( .DIN1(n422), .DIN2(n7506), .Q(n7502) );
  or2s1 U8227 ( .DIN1(n7386), .DIN2(n706), .Q(n7500) );
  nnd2s1 U8228 ( .DIN1(n7507), .DIN2(n7508), .Q(n7386) );
  nnd2s1 U8229 ( .DIN1(n7509), .DIN2(n7510), .Q(n7508) );
  nnd2s1 U8230 ( .DIN1(n7138), .DIN2(n5794), .Q(n7491) );
  nnd3s1 U8231 ( .DIN1(n7511), .DIN2(n7512), .DIN3(n7513), .Q(n5794) );
  nnd2s1 U8232 ( .DIN1(n61), .DIN2(n6658), .Q(n7513) );
  nnd2s1 U8233 ( .DIN1(n622), .DIN2(n6652), .Q(n7512) );
  nnd2s1 U8234 ( .DIN1(n630), .DIN2(n6224), .Q(n7511) );
  nnd4s1 U8235 ( .DIN1(n7514), .DIN2(n7515), .DIN3(n7516), .DIN4(n7517), 
        .Q(n6224) );
  nnd2s1 U8236 ( .DIN1(n531), .DIN2(n424), .Q(n7516) );
  nnd2s1 U8237 ( .DIN1(n421), .DIN2(n768), .Q(n7490) );
  nnd2s1 U8238 ( .DIN1(reg_out_B[12]), .DIN2(n7518), .Q(n7488) );
  nnd2s1 U8239 ( .DIN1(n5471), .DIN2(n7519), .Q(n7518) );
  nnd2s1 U8240 ( .DIN1(n775), .DIN2(n421), .Q(n7519) );
  nnd3s1 U8241 ( .DIN1(n7520), .DIN2(n7521), .DIN3(n5336), .Q(n7487) );
  nnd4s1 U8242 ( .DIN1(n7399), .DIN2(n7522), .DIN3(n7523), .DIN4(n7524), 
        .Q(n7521) );
  nnd2s1 U8243 ( .DIN1(n5769), .DIN2(n752), .Q(n7524) );
  nnd2s1 U8244 ( .DIN1(n7525), .DIN2(n808), .Q(n7523) );
  nnd2s1 U8245 ( .DIN1(n5345), .DIN2(n7526), .Q(n7522) );
  nnd2s1 U8246 ( .DIN1(n7154), .DIN2(n7527), .Q(n7520) );
  nnd2s1 U8247 ( .DIN1(n7283), .DIN2(n801), .Q(n7527) );
  nnd2s1 U8248 ( .DIN1(n7528), .DIN2(n7529), .Q(n7486) );
  nnd3s1 U8249 ( .DIN1(n7530), .DIN2(n807), .DIN3(n7531), .Q(n7529) );
  hi1s1 U8250 ( .DIN(n7525), .Q(n7531) );
  nnd3s1 U8251 ( .DIN1(n7532), .DIN2(n7533), .DIN3(n7534), .Q(n7525) );
  nnd2s1 U8252 ( .DIN1(n621), .DIN2(n7535), .Q(n7534) );
  nnd2s1 U8253 ( .DIN1(n720), .DIN2(n7536), .Q(n7533) );
  nnd2s1 U8254 ( .DIN1(n547), .DIN2(n7537), .Q(n7532) );
  nnd2s1 U8255 ( .DIN1(n629), .DIN2(n7526), .Q(n7530) );
  nnd2s1 U8256 ( .DIN1(n5994), .DIN2(n7538), .Q(n7528) );
  nnd2s1 U8257 ( .DIN1(n386), .DIN2(n5769), .Q(n7538) );
  and2s1 U8258 ( .DIN1(n630), .DIN2(n7539), .Q(n5769) );
  nnd2s1 U8259 ( .DIN1(n550), .DIN2(n7540), .Q(n7482) );
  nnd4s1 U8260 ( .DIN1(n7541), .DIN2(n7542), .DIN3(n7543), .DIN4(n7544), 
        .Q(n7540) );
  and4s1 U8261 ( .DIN1(n7545), .DIN2(n7546), .DIN3(n7547), .DIN4(n7548), 
        .Q(n7544) );
  nnd2s1 U8262 ( .DIN1(n421), .DIN2(n7549), .Q(n7548) );
  nnd4s1 U8263 ( .DIN1(n7550), .DIN2(n7551), .DIN3(n7552), .DIN4(n7059), 
        .Q(n7549) );
  nnd2s1 U8264 ( .DIN1(n7553), .DIN2(n7212), .Q(n7552) );
  xnr2s1 U8265 ( .DIN1(n7476), .DIN2(n7475), .Q(n7553) );
  hi1s1 U8266 ( .DIN(n7554), .Q(n7475) );
  nnd2s1 U8267 ( .DIN1(n7555), .DIN2(n743), .Q(n7551) );
  xnr2s1 U8268 ( .DIN1(n389), .DIN2(n7481), .Q(n7555) );
  hi1s1 U8269 ( .DIN(n7556), .Q(n7481) );
  nnd2s1 U8270 ( .DIN1(n7314), .DIN2(n106), .Q(n7550) );
  nnd2s1 U8271 ( .DIN1(n7557), .DIN2(n64), .Q(n7547) );
  nnd2s1 U8272 ( .DIN1(n7558), .DIN2(n7559), .Q(n7557) );
  nnd2s1 U8273 ( .DIN1(n7560), .DIN2(n722), .Q(n7559) );
  xnr2s1 U8274 ( .DIN1(n7554), .DIN2(n7476), .Q(n7560) );
  xor2s1 U8275 ( .DIN1(n9479), .DIN2(n745), .Q(n7476) );
  nnd2s1 U8276 ( .DIN1(n7561), .DIN2(n7562), .Q(n7554) );
  nnd2s1 U8277 ( .DIN1(n422), .DIN2(n7563), .Q(n7562) );
  or2s1 U8278 ( .DIN1(n7564), .DIN2(n7565), .Q(n7563) );
  nnd2s1 U8279 ( .DIN1(n7565), .DIN2(n7564), .Q(n7561) );
  nnd2s1 U8280 ( .DIN1(n7566), .DIN2(n7058), .Q(n7558) );
  xnr2s1 U8281 ( .DIN1(n7556), .DIN2(n389), .Q(n7566) );
  nnd2s1 U8282 ( .DIN1(n7567), .DIN2(n7568), .Q(n7556) );
  nnd2s1 U8283 ( .DIN1(n422), .DIN2(n7569), .Q(n7568) );
  or2s1 U8284 ( .DIN1(n7570), .DIN2(n7571), .Q(n7569) );
  nnd2s1 U8285 ( .DIN1(n7571), .DIN2(n7570), .Q(n7567) );
  nnd2s1 U8286 ( .DIN1(n400), .DIN2(n5735), .Q(n7546) );
  nnd3s1 U8287 ( .DIN1(n7572), .DIN2(n7573), .DIN3(n7574), .Q(n5735) );
  nnd2s1 U8288 ( .DIN1(n6610), .DIN2(n803), .Q(n7574) );
  nnd2s1 U8289 ( .DIN1(n544), .DIN2(n6608), .Q(n7573) );
  nnd2s1 U8290 ( .DIN1(n555), .DIN2(n6176), .Q(n7572) );
  nnd4s1 U8291 ( .DIN1(n7575), .DIN2(n7576), .DIN3(n7577), .DIN4(n7578), 
        .Q(n6176) );
  nnd2s1 U8292 ( .DIN1(n758), .DIN2(n424), .Q(n7577) );
  nnd2s1 U8293 ( .DIN1(n7206), .DIN2(n106), .Q(n7545) );
  or2s1 U8294 ( .DIN1(n7579), .DIN2(n7006), .Q(n7543) );
  nnd4s1 U8295 ( .DIN1(n7580), .DIN2(n7581), .DIN3(n7433), .DIN4(n7582), 
        .Q(n7542) );
  and3s1 U8296 ( .DIN1(n7583), .DIN2(n7584), .DIN3(n7585), .Q(n7582) );
  nnd2s1 U8297 ( .DIN1(n7586), .DIN2(n700), .Q(n7585) );
  nnd2s1 U8298 ( .DIN1(n7587), .DIN2(n5824), .Q(n7584) );
  nnd2s1 U8299 ( .DIN1(n7588), .DIN2(n726), .Q(n7583) );
  and2s1 U8300 ( .DIN1(n730), .DIN2(n7589), .Q(n7433) );
  nnd2s1 U8301 ( .DIN1(n6253), .DIN2(n805), .Q(n7589) );
  nnd2s1 U8302 ( .DIN1(n7590), .DIN2(n544), .Q(n7581) );
  nnd2s1 U8303 ( .DIN1(n7591), .DIN2(n806), .Q(n7580) );
  nnd3s1 U8304 ( .DIN1(n7592), .DIN2(n7593), .DIN3(n7594), .Q(n7541) );
  nnd4s1 U8305 ( .DIN1(n7595), .DIN2(n7596), .DIN3(n7447), .DIN4(n7597), 
        .Q(n7593) );
  and3s1 U8306 ( .DIN1(n7598), .DIN2(n7599), .DIN3(n7600), .Q(n7597) );
  nnd2s1 U8307 ( .DIN1(n719), .DIN2(n7601), .Q(n7600) );
  nnd2s1 U8308 ( .DIN1(n7453), .DIN2(n5742), .Q(n7599) );
  nnd2s1 U8309 ( .DIN1(n5315), .DIN2(n7602), .Q(n7598) );
  nnd2s1 U8310 ( .DIN1(n398), .DIN2(n7603), .Q(n7596) );
  nnd2s1 U8311 ( .DIN1(n5306), .DIN2(n7604), .Q(n7595) );
  nnd2s1 U8312 ( .DIN1(n7605), .DIN2(n7606), .Q(n7592) );
  nnd3s1 U8313 ( .DIN1(n6379), .DIN2(n736), .DIN3(n6465), .Q(n7606) );
  nnd3s1 U8314 ( .DIN1(n7607), .DIN2(n7608), .DIN3(n7609), .Q(\EXinst/n1443 )
         );
  nnd2s1 U8315 ( .DIN1(n727), .DIN2(\DM_addr[11] ), .Q(n7609) );
  nnd2s1 U8316 ( .DIN1(n5324), .DIN2(n7610), .Q(n7608) );
  nnd4s1 U8317 ( .DIN1(n7611), .DIN2(n7612), .DIN3(n7613), .DIN4(n7614), 
        .Q(n7610) );
  and4s1 U8318 ( .DIN1(n7615), .DIN2(n7616), .DIN3(n7617), .DIN4(n7618), 
        .Q(n7614) );
  nnd2s1 U8319 ( .DIN1(n7619), .DIN2(n7620), .Q(n7618) );
  nnd3s1 U8320 ( .DIN1(n7621), .DIN2(n749), .DIN3(n7622), .Q(n7619) );
  nnd2s1 U8321 ( .DIN1(n705), .DIN2(n7509), .Q(n7622) );
  nnd2s1 U8322 ( .DIN1(n654), .DIN2(n7505), .Q(n7621) );
  hi1s1 U8323 ( .DIN(n7506), .Q(n7505) );
  nnd2s1 U8324 ( .DIN1(n7623), .DIN2(n7624), .Q(n7617) );
  nnd2s1 U8325 ( .DIN1(n7625), .DIN2(n7626), .Q(n7624) );
  nnd2s1 U8326 ( .DIN1(n653), .DIN2(n7506), .Q(n7626) );
  nnd2s1 U8327 ( .DIN1(n7627), .DIN2(n7628), .Q(n7506) );
  nnd2s1 U8328 ( .DIN1(reg_out_B[10]), .DIN2(n7629), .Q(n7628) );
  nnd2s1 U8329 ( .DIN1(n7630), .DIN2(n65), .Q(n7629) );
  nnd2s1 U8330 ( .DIN1(n423), .DIN2(n7631), .Q(n7627) );
  or2s1 U8331 ( .DIN1(n7509), .DIN2(n5375), .Q(n7625) );
  nnd2s1 U8332 ( .DIN1(n7632), .DIN2(n7633), .Q(n7509) );
  nnd2s1 U8333 ( .DIN1(n7634), .DIN2(n7635), .Q(n7633) );
  nnd2s1 U8334 ( .DIN1(n7138), .DIN2(n5882), .Q(n7616) );
  nnd3s1 U8335 ( .DIN1(n7636), .DIN2(n7637), .DIN3(n7638), .Q(n5882) );
  nnd2s1 U8336 ( .DIN1(n630), .DIN2(n6309), .Q(n7638) );
  nnd4s1 U8337 ( .DIN1(n7639), .DIN2(n7640), .DIN3(n7641), .DIN4(n7642), 
        .Q(n6309) );
  nnd2s1 U8338 ( .DIN1(n772), .DIN2(n424), .Q(n7642) );
  nnd2s1 U8339 ( .DIN1(n532), .DIN2(n36), .Q(n7641) );
  nnd2s1 U8340 ( .DIN1(n546), .DIN2(n6745), .Q(n7637) );
  nnd2s1 U8341 ( .DIN1(n623), .DIN2(n7143), .Q(n7636) );
  nnd2s1 U8342 ( .DIN1(n422), .DIN2(n767), .Q(n7615) );
  nnd2s1 U8343 ( .DIN1(reg_out_B[11]), .DIN2(n7643), .Q(n7613) );
  nnd2s1 U8344 ( .DIN1(n5471), .DIN2(n7644), .Q(n7643) );
  nnd2s1 U8345 ( .DIN1(n776), .DIN2(n422), .Q(n7644) );
  nnd3s1 U8346 ( .DIN1(n7645), .DIN2(n7646), .DIN3(n769), .Q(n7612) );
  nnd4s1 U8347 ( .DIN1(n7399), .DIN2(n7647), .DIN3(n7648), .DIN4(n7649), 
        .Q(n7646) );
  nnd2s1 U8348 ( .DIN1(n7650), .DIN2(n204), .Q(n7649) );
  nnd3s1 U8349 ( .DIN1(n628), .DIN2(n5863), .DIN3(n55), .Q(n7648) );
  nnd2s1 U8350 ( .DIN1(n5345), .DIN2(n7651), .Q(n7647) );
  and2s1 U8351 ( .DIN1(n5337), .DIN2(n7652), .Q(n7399) );
  nnd2s1 U8352 ( .DIN1(n752), .DIN2(n5864), .Q(n7652) );
  nnd2s1 U8353 ( .DIN1(n6294), .DIN2(n7653), .Q(n5864) );
  nnd2s1 U8354 ( .DIN1(n7156), .DIN2(n742), .Q(n7653) );
  hi1s1 U8355 ( .DIN(n6216), .Q(n6294) );
  nnd2s1 U8356 ( .DIN1(n7154), .DIN2(n7654), .Q(n7645) );
  nnd2s1 U8357 ( .DIN1(n7156), .DIN2(n5867), .Q(n7654) );
  nnd2s1 U8358 ( .DIN1(n7655), .DIN2(n7656), .Q(n7611) );
  nnd3s1 U8359 ( .DIN1(n7657), .DIN2(n807), .DIN3(n7658), .Q(n7656) );
  hi1s1 U8360 ( .DIN(n7650), .Q(n7658) );
  nnd3s1 U8361 ( .DIN1(n7659), .DIN2(n7660), .DIN3(n7661), .Q(n7650) );
  nnd2s1 U8362 ( .DIN1(n622), .DIN2(n7163), .Q(n7661) );
  nnd2s1 U8363 ( .DIN1(n5876), .DIN2(n6729), .Q(n7660) );
  nnd2s1 U8364 ( .DIN1(n547), .DIN2(n6728), .Q(n7659) );
  nnd2s1 U8365 ( .DIN1(n629), .DIN2(n7651), .Q(n7657) );
  nnd2s1 U8366 ( .DIN1(n5994), .DIN2(n7662), .Q(n7655) );
  nnd2s1 U8367 ( .DIN1(n7165), .DIN2(n5857), .Q(n7662) );
  nnd2s1 U8368 ( .DIN1(n551), .DIN2(n7663), .Q(n7607) );
  nnd4s1 U8369 ( .DIN1(n7664), .DIN2(n7665), .DIN3(n7666), .DIN4(n7667), 
        .Q(n7663) );
  and3s1 U8370 ( .DIN1(n7668), .DIN2(n7669), .DIN3(n7670), .Q(n7667) );
  nnd2s1 U8371 ( .DIN1(n400), .DIN2(n5829), .Q(n7670) );
  nnd3s1 U8372 ( .DIN1(n7671), .DIN2(n7672), .DIN3(n7673), .Q(n5829) );
  nnd2s1 U8373 ( .DIN1(n554), .DIN2(n6258), .Q(n7673) );
  nnd4s1 U8374 ( .DIN1(n7674), .DIN2(n7675), .DIN3(n7676), .DIN4(n7677), 
        .Q(n6258) );
  nnd2s1 U8375 ( .DIN1(n784), .DIN2(n424), .Q(n7677) );
  nnd2s1 U8376 ( .DIN1(n758), .DIN2(n425), .Q(n7676) );
  nnd2s1 U8377 ( .DIN1(n5826), .DIN2(n6689), .Q(n7672) );
  nnd2s1 U8378 ( .DIN1(n545), .DIN2(n6686), .Q(n7671) );
  nnd4s1 U8379 ( .DIN1(n7678), .DIN2(n7679), .DIN3(n7680), .DIN4(n7681), 
        .Q(n7669) );
  and3s1 U8380 ( .DIN1(n7682), .DIN2(n7683), .DIN3(n7188), .Q(n7681) );
  nnd2s1 U8381 ( .DIN1(n7684), .DIN2(n700), .Q(n7683) );
  or2s1 U8382 ( .DIN1(n5830), .DIN2(n739), .Q(n7682) );
  nnd2s1 U8383 ( .DIN1(n7204), .DIN2(n397), .Q(n7680) );
  nnd2s1 U8384 ( .DIN1(n7192), .DIN2(n5824), .Q(n7679) );
  nnd2s1 U8385 ( .DIN1(n7189), .DIN2(n726), .Q(n7678) );
  nnd3s1 U8386 ( .DIN1(n7685), .DIN2(n7686), .DIN3(n7594), .Q(n7668) );
  nnd4s1 U8387 ( .DIN1(n7687), .DIN2(n7688), .DIN3(n7447), .DIN4(n7689), 
        .Q(n7686) );
  and3s1 U8388 ( .DIN1(n7690), .DIN2(n7691), .DIN3(n7692), .Q(n7689) );
  nnd2s1 U8389 ( .DIN1(n5304), .DIN2(n7203), .Q(n7692) );
  nnd2s1 U8390 ( .DIN1(n7453), .DIN2(n5807), .Q(n7691) );
  nor2s1 U8391 ( .DIN1(n6253), .DIN2(n739), .Q(n7453) );
  nnd2s1 U8392 ( .DIN1(n5315), .DIN2(n7693), .Q(n7690) );
  and2s1 U8393 ( .DIN1(n9486), .DIN2(n7694), .Q(n7447) );
  nnd2s1 U8394 ( .DIN1(n5809), .DIN2(n805), .Q(n7694) );
  nnd2s1 U8395 ( .DIN1(n5556), .DIN2(n7695), .Q(n5809) );
  nnd2s1 U8396 ( .DIN1(n5321), .DIN2(n792), .Q(n7695) );
  nnd2s1 U8397 ( .DIN1(n397), .DIN2(n7696), .Q(n7688) );
  nnd2s1 U8398 ( .DIN1(n5306), .DIN2(n7697), .Q(n7687) );
  nnd2s1 U8399 ( .DIN1(n7605), .DIN2(n7698), .Q(n7685) );
  nnd3s1 U8400 ( .DIN1(n6379), .DIN2(n5811), .DIN3(n5321), .Q(n7698) );
  nnd2s1 U8401 ( .DIN1(n7206), .DIN2(n8), .Q(n7666) );
  nnd2s1 U8402 ( .DIN1(n422), .DIN2(n7699), .Q(n7665) );
  nnd4s1 U8403 ( .DIN1(n7700), .DIN2(n7701), .DIN3(n7702), .DIN4(n7059), 
        .Q(n7699) );
  nnd2s1 U8404 ( .DIN1(n7703), .DIN2(n7212), .Q(n7702) );
  xnr2s1 U8405 ( .DIN1(n7564), .DIN2(n7565), .Q(n7703) );
  hi1s1 U8406 ( .DIN(n7704), .Q(n7565) );
  nnd2s1 U8407 ( .DIN1(n7705), .DIN2(n743), .Q(n7701) );
  xnr2s1 U8408 ( .DIN1(n7570), .DIN2(n7571), .Q(n7705) );
  hi1s1 U8409 ( .DIN(n7706), .Q(n7571) );
  nor2s1 U8410 ( .DIN1(n7707), .DIN2(n7708), .Q(n7700) );
  nor2s1 U8411 ( .DIN1(n8), .DIN2(n7006), .Q(n7708) );
  nor2s1 U8412 ( .DIN1(n9480), .DIN2(n7037), .Q(n7707) );
  nnd2s1 U8413 ( .DIN1(n7709), .DIN2(n84), .Q(n7664) );
  nnd3s1 U8414 ( .DIN1(n7710), .DIN2(n7711), .DIN3(n7712), .Q(n7709) );
  nnd2s1 U8415 ( .DIN1(n7222), .DIN2(n8), .Q(n7712) );
  nnd2s1 U8416 ( .DIN1(n7713), .DIN2(n722), .Q(n7711) );
  xnr2s1 U8417 ( .DIN1(n7564), .DIN2(n7704), .Q(n7713) );
  xnr2s1 U8418 ( .DIN1(n9480), .DIN2(n786), .Q(n7704) );
  nnd2s1 U8419 ( .DIN1(n7714), .DIN2(n7715), .Q(n7564) );
  nnd2s1 U8420 ( .DIN1(n423), .DIN2(n7716), .Q(n7715) );
  nnd2s1 U8421 ( .DIN1(n7717), .DIN2(n7718), .Q(n7716) );
  or2s1 U8422 ( .DIN1(n7718), .DIN2(n7717), .Q(n7714) );
  nnd2s1 U8423 ( .DIN1(n7719), .DIN2(n7058), .Q(n7710) );
  xnr2s1 U8424 ( .DIN1(n7570), .DIN2(n7706), .Q(n7719) );
  xnr2s1 U8425 ( .DIN1(n633), .DIN2(n8), .Q(n7706) );
  nnd2s1 U8426 ( .DIN1(n7720), .DIN2(n7721), .Q(n7570) );
  nnd2s1 U8427 ( .DIN1(n423), .DIN2(n7722), .Q(n7721) );
  nnd2s1 U8428 ( .DIN1(n7723), .DIN2(n390), .Q(n7722) );
  or2s1 U8429 ( .DIN1(n390), .DIN2(n7723), .Q(n7720) );
  nnd3s1 U8430 ( .DIN1(n7724), .DIN2(n7725), .DIN3(n7726), .Q(\EXinst/n1442 )
         );
  nnd2s1 U8431 ( .DIN1(n5394), .DIN2(\DM_addr[10] ), .Q(n7726) );
  nnd2s1 U8432 ( .DIN1(n5324), .DIN2(n7727), .Q(n7725) );
  nnd4s1 U8433 ( .DIN1(n7728), .DIN2(n7729), .DIN3(n7730), .DIN4(n7731), 
        .Q(n7727) );
  and4s1 U8434 ( .DIN1(n7732), .DIN2(n7733), .DIN3(n7734), .DIN4(n7735), 
        .Q(n7731) );
  nnd2s1 U8435 ( .DIN1(n7736), .DIN2(n7737), .Q(n7735) );
  nnd3s1 U8436 ( .DIN1(n7738), .DIN2(n5372), .DIN3(n7739), .Q(n7736) );
  nnd2s1 U8437 ( .DIN1(n620), .DIN2(n7635), .Q(n7739) );
  nnd2s1 U8438 ( .DIN1(n656), .DIN2(n7630), .Q(n7738) );
  hi1s1 U8439 ( .DIN(n7631), .Q(n7630) );
  nnd2s1 U8440 ( .DIN1(n7740), .DIN2(n7741), .Q(n7734) );
  nnd2s1 U8441 ( .DIN1(n7742), .DIN2(n7743), .Q(n7741) );
  nnd2s1 U8442 ( .DIN1(n655), .DIN2(n7631), .Q(n7743) );
  nnd2s1 U8443 ( .DIN1(n7744), .DIN2(n7745), .Q(n7631) );
  nnd2s1 U8444 ( .DIN1(reg_out_B[9]), .DIN2(n7746), .Q(n7745) );
  nnd2s1 U8445 ( .DIN1(n7747), .DIN2(n66), .Q(n7746) );
  nnd2s1 U8446 ( .DIN1(n424), .DIN2(n7748), .Q(n7744) );
  or2s1 U8447 ( .DIN1(n7635), .DIN2(n5375), .Q(n7742) );
  nnd2s1 U8448 ( .DIN1(n7749), .DIN2(n7750), .Q(n7635) );
  nnd2s1 U8449 ( .DIN1(n7751), .DIN2(n7752), .Q(n7750) );
  nnd2s1 U8450 ( .DIN1(n7138), .DIN2(n6018), .Q(n7733) );
  nnd3s1 U8451 ( .DIN1(n7753), .DIN2(n7754), .DIN3(n7755), .Q(n6018) );
  nnd2s1 U8452 ( .DIN1(n630), .DIN2(n6445), .Q(n7755) );
  nnd4s1 U8453 ( .DIN1(n7756), .DIN2(n7757), .DIN3(n7758), .DIN4(n7759), 
        .Q(n6445) );
  nnd2s1 U8454 ( .DIN1(n771), .DIN2(n36), .Q(n7759) );
  nnd2s1 U8455 ( .DIN1(n546), .DIN2(n6879), .Q(n7754) );
  nnd2s1 U8456 ( .DIN1(n621), .DIN2(n7267), .Q(n7753) );
  nnd2s1 U8457 ( .DIN1(n423), .DIN2(n768), .Q(n7732) );
  nnd2s1 U8458 ( .DIN1(reg_out_B[10]), .DIN2(n7760), .Q(n7730) );
  nnd2s1 U8459 ( .DIN1(n5471), .DIN2(n7761), .Q(n7760) );
  nnd2s1 U8460 ( .DIN1(n775), .DIN2(n423), .Q(n7761) );
  nnd3s1 U8461 ( .DIN1(n7762), .DIN2(n7763), .DIN3(n5336), .Q(n7729) );
  nnd2s1 U8462 ( .DIN1(n7154), .DIN2(n7764), .Q(n7763) );
  nnd2s1 U8463 ( .DIN1(n7156), .DIN2(n7765), .Q(n7764) );
  nnd4s1 U8464 ( .DIN1(n7276), .DIN2(n7766), .DIN3(n7767), .DIN4(n7768), 
        .Q(n7762) );
  nnd2s1 U8465 ( .DIN1(n7769), .DIN2(n808), .Q(n7768) );
  nnd3s1 U8466 ( .DIN1(n6000), .DIN2(n337), .DIN3(n752), .Q(n7767) );
  nnd2s1 U8467 ( .DIN1(n5345), .DIN2(n7770), .Q(n7766) );
  nnd2s1 U8468 ( .DIN1(n7771), .DIN2(n7772), .Q(n7728) );
  nnd3s1 U8469 ( .DIN1(n7773), .DIN2(n807), .DIN3(n7774), .Q(n7772) );
  hi1s1 U8470 ( .DIN(n7769), .Q(n7774) );
  nnd3s1 U8471 ( .DIN1(n7775), .DIN2(n7776), .DIN3(n7777), .Q(n7769) );
  nnd2s1 U8472 ( .DIN1(n623), .DIN2(n7281), .Q(n7777) );
  nnd2s1 U8473 ( .DIN1(n5876), .DIN2(n7293), .Q(n7776) );
  nnd2s1 U8474 ( .DIN1(n547), .DIN2(n7291), .Q(n7775) );
  nnd2s1 U8475 ( .DIN1(n629), .DIN2(n7770), .Q(n7773) );
  nnd2s1 U8476 ( .DIN1(n5994), .DIN2(n7778), .Q(n7771) );
  nnd2s1 U8477 ( .DIN1(n7165), .DIN2(n5993), .Q(n7778) );
  and2s1 U8478 ( .DIN1(n386), .DIN2(n801), .Q(n7165) );
  nnd2s1 U8479 ( .DIN1(n551), .DIN2(n7779), .Q(n7724) );
  nnd4s1 U8480 ( .DIN1(n7780), .DIN2(n7781), .DIN3(n7782), .DIN4(n7783), 
        .Q(n7779) );
  and4s1 U8481 ( .DIN1(n7784), .DIN2(n7785), .DIN3(n7786), .DIN4(n7787), 
        .Q(n7783) );
  nnd2s1 U8482 ( .DIN1(n423), .DIN2(n7788), .Q(n7787) );
  nnd4s1 U8483 ( .DIN1(n7789), .DIN2(n7790), .DIN3(n7791), .DIN4(n7059), 
        .Q(n7788) );
  nnd2s1 U8484 ( .DIN1(n7792), .DIN2(n7212), .Q(n7791) );
  xnr2s1 U8485 ( .DIN1(n7718), .DIN2(n7717), .Q(n7792) );
  hi1s1 U8486 ( .DIN(n7793), .Q(n7717) );
  nnd2s1 U8487 ( .DIN1(n7794), .DIN2(n743), .Q(n7790) );
  xnr2s1 U8488 ( .DIN1(n390), .DIN2(n7723), .Q(n7794) );
  hi1s1 U8489 ( .DIN(n7795), .Q(n7723) );
  nnd2s1 U8490 ( .DIN1(n7314), .DIN2(n104), .Q(n7789) );
  nnd2s1 U8491 ( .DIN1(n7796), .DIN2(n65), .Q(n7786) );
  nnd2s1 U8492 ( .DIN1(n7797), .DIN2(n7798), .Q(n7796) );
  nnd2s1 U8493 ( .DIN1(n7799), .DIN2(n722), .Q(n7798) );
  xnr2s1 U8494 ( .DIN1(n7793), .DIN2(n7718), .Q(n7799) );
  xor2s1 U8495 ( .DIN1(n9481), .DIN2(n5413), .Q(n7718) );
  nnd2s1 U8496 ( .DIN1(n7800), .DIN2(n7801), .Q(n7793) );
  nnd2s1 U8497 ( .DIN1(n424), .DIN2(n7802), .Q(n7801) );
  or2s1 U8498 ( .DIN1(n7803), .DIN2(n7804), .Q(n7802) );
  nnd2s1 U8499 ( .DIN1(n7804), .DIN2(n7803), .Q(n7800) );
  nnd2s1 U8500 ( .DIN1(n7805), .DIN2(n7058), .Q(n7797) );
  xnr2s1 U8501 ( .DIN1(n7795), .DIN2(n390), .Q(n7805) );
  nnd2s1 U8502 ( .DIN1(n7806), .DIN2(n7807), .Q(n7795) );
  nnd2s1 U8503 ( .DIN1(n424), .DIN2(n7808), .Q(n7807) );
  or2s1 U8504 ( .DIN1(n7809), .DIN2(n7810), .Q(n7808) );
  nnd2s1 U8505 ( .DIN1(n7810), .DIN2(n7809), .Q(n7806) );
  nnd2s1 U8506 ( .DIN1(n400), .DIN2(n5966), .Q(n7785) );
  nnd3s1 U8507 ( .DIN1(n7811), .DIN2(n7812), .DIN3(n7813), .Q(n5966) );
  nnd2s1 U8508 ( .DIN1(n555), .DIN2(n6399), .Q(n7813) );
  nnd4s1 U8509 ( .DIN1(n7814), .DIN2(n7815), .DIN3(n7816), .DIN4(n7817), 
        .Q(n6399) );
  nnd2s1 U8510 ( .DIN1(n783), .DIN2(n425), .Q(n7817) );
  nnd2s1 U8511 ( .DIN1(n5826), .DIN2(n6830), .Q(n7812) );
  nnd2s1 U8512 ( .DIN1(n544), .DIN2(n6828), .Q(n7811) );
  nnd2s1 U8513 ( .DIN1(n7206), .DIN2(n104), .Q(n7784) );
  or2s1 U8514 ( .DIN1(n7818), .DIN2(n7006), .Q(n7782) );
  nnd4s1 U8515 ( .DIN1(n7819), .DIN2(n7188), .DIN3(n7820), .DIN4(n7821), 
        .Q(n7781) );
  or2s1 U8516 ( .DIN1(n5943), .DIN2(n740), .Q(n7821) );
  nor2s1 U8517 ( .DIN1(n7822), .DIN2(n7823), .Q(n7820) );
  and2s1 U8518 ( .DIN1(n726), .DIN2(n7356), .Q(n7823) );
  and2s1 U8519 ( .DIN1(n5824), .DIN2(n6386), .Q(n7822) );
  and2s1 U8520 ( .DIN1(n730), .DIN2(n7824), .Q(n7188) );
  nnd2s1 U8521 ( .DIN1(n4840), .DIN2(n806), .Q(n7824) );
  nnd4s1 U8522 ( .DIN1(n7346), .DIN2(n7825), .DIN3(n7826), .DIN4(n7827), 
        .Q(n7780) );
  nnd2s1 U8523 ( .DIN1(n7350), .DIN2(n5951), .Q(n7827) );
  and2s1 U8524 ( .DIN1(n7828), .DIN2(n7196), .Q(n7826) );
  nnd3s1 U8525 ( .DIN1(n5741), .DIN2(n707), .DIN3(n7205), .Q(n7828) );
  nnd2s1 U8526 ( .DIN1(n733), .DIN2(n7829), .Q(n7825) );
  nnd3s1 U8527 ( .DIN1(n7830), .DIN2(n7831), .DIN3(n7819), .Q(n7829) );
  and2s1 U8528 ( .DIN1(n7832), .DIN2(n7833), .Q(n7819) );
  nnd2s1 U8529 ( .DIN1(n7357), .DIN2(n398), .Q(n7833) );
  nnd2s1 U8530 ( .DIN1(n7834), .DIN2(n700), .Q(n7832) );
  nnd2s1 U8531 ( .DIN1(n7356), .DIN2(n763), .Q(n7831) );
  nnd2s1 U8532 ( .DIN1(n6386), .DIN2(n719), .Q(n7830) );
  and2s1 U8533 ( .DIN1(n7193), .DIN2(n7835), .Q(n7346) );
  nnd2s1 U8534 ( .DIN1(n7350), .DIN2(n735), .Q(n7835) );
  and2s1 U8535 ( .DIN1(n7836), .DIN2(n5556), .Q(n7350) );
  nnd3s1 U8536 ( .DIN1(n7837), .DIN2(n7838), .DIN3(n7839), .Q(\EXinst/n1441 )
         );
  nnd2s1 U8537 ( .DIN1(n727), .DIN2(\DM_addr[9] ), .Q(n7839) );
  nnd2s1 U8538 ( .DIN1(n5324), .DIN2(n7840), .Q(n7838) );
  nnd4s1 U8539 ( .DIN1(n7841), .DIN2(n7842), .DIN3(n7843), .DIN4(n7844), 
        .Q(n7840) );
  and4s1 U8540 ( .DIN1(n7845), .DIN2(n7846), .DIN3(n7847), .DIN4(n7848), 
        .Q(n7844) );
  nnd2s1 U8541 ( .DIN1(n7849), .DIN2(n7850), .Q(n7848) );
  nnd3s1 U8542 ( .DIN1(n7851), .DIN2(n749), .DIN3(n7852), .Q(n7849) );
  nnd2s1 U8543 ( .DIN1(n705), .DIN2(n7751), .Q(n7852) );
  nnd2s1 U8544 ( .DIN1(n654), .DIN2(n7747), .Q(n7851) );
  hi1s1 U8545 ( .DIN(n7748), .Q(n7747) );
  nnd2s1 U8546 ( .DIN1(n7853), .DIN2(n7854), .Q(n7847) );
  nnd2s1 U8547 ( .DIN1(n7855), .DIN2(n7856), .Q(n7854) );
  nnd2s1 U8548 ( .DIN1(n653), .DIN2(n7748), .Q(n7856) );
  nnd2s1 U8549 ( .DIN1(n7857), .DIN2(n7858), .Q(n7748) );
  nnd2s1 U8550 ( .DIN1(reg_out_B[8]), .DIN2(n7859), .Q(n7858) );
  nnd2s1 U8551 ( .DIN1(n7860), .DIN2(n332), .Q(n7859) );
  nnd2s1 U8552 ( .DIN1(n425), .DIN2(n7861), .Q(n7857) );
  or2s1 U8553 ( .DIN1(n7751), .DIN2(n5375), .Q(n7855) );
  nnd2s1 U8554 ( .DIN1(n7862), .DIN2(n7863), .Q(n7751) );
  nnd2s1 U8555 ( .DIN1(n7864), .DIN2(n7865), .Q(n7863) );
  nnd2s1 U8556 ( .DIN1(n7138), .DIN2(n6102), .Q(n7846) );
  nnd3s1 U8557 ( .DIN1(n7866), .DIN2(n7867), .DIN3(n7868), .Q(n6102) );
  nnd2s1 U8558 ( .DIN1(n630), .DIN2(n6524), .Q(n7868) );
  nnd4s1 U8559 ( .DIN1(n7869), .DIN2(n7870), .DIN3(n7871), .DIN4(n7872), 
        .Q(n6524) );
  nnd2s1 U8560 ( .DIN1(n772), .DIN2(n429), .Q(n7872) );
  nnd2s1 U8561 ( .DIN1(n546), .DIN2(n7873), .Q(n7867) );
  nnd2s1 U8562 ( .DIN1(n622), .DIN2(n6957), .Q(n7866) );
  nnd2s1 U8563 ( .DIN1(n424), .DIN2(n767), .Q(n7845) );
  nnd2s1 U8564 ( .DIN1(reg_out_B[9]), .DIN2(n7874), .Q(n7843) );
  nnd2s1 U8565 ( .DIN1(n5471), .DIN2(n7875), .Q(n7874) );
  nnd2s1 U8566 ( .DIN1(n776), .DIN2(n424), .Q(n7875) );
  nnd3s1 U8567 ( .DIN1(n7876), .DIN2(n7877), .DIN3(n769), .Q(n7842) );
  nnd4s1 U8568 ( .DIN1(n7276), .DIN2(n7878), .DIN3(n7879), .DIN4(n7880), 
        .Q(n7877) );
  nnd2s1 U8569 ( .DIN1(n753), .DIN2(n6085), .Q(n7880) );
  nnd2s1 U8570 ( .DIN1(n7881), .DIN2(n7882), .Q(n6085) );
  nnd2s1 U8571 ( .DIN1(n621), .DIN2(n5651), .Q(n7882) );
  nnd2s1 U8572 ( .DIN1(n629), .DIN2(n7413), .Q(n7881) );
  nnd2s1 U8573 ( .DIN1(n7883), .DIN2(n204), .Q(n7879) );
  nnd2s1 U8574 ( .DIN1(n5345), .DIN2(n7884), .Q(n7878) );
  nnd2s1 U8575 ( .DIN1(n7154), .DIN2(n7885), .Q(n7876) );
  nnd2s1 U8576 ( .DIN1(n7156), .DIN2(n6087), .Q(n7885) );
  hi1s1 U8577 ( .DIN(n7089), .Q(n7154) );
  nnd2s1 U8578 ( .DIN1(n7886), .DIN2(n7887), .Q(n7841) );
  nnd3s1 U8579 ( .DIN1(n7888), .DIN2(n807), .DIN3(n7889), .Q(n7887) );
  hi1s1 U8580 ( .DIN(n7883), .Q(n7889) );
  nnd3s1 U8581 ( .DIN1(n7890), .DIN2(n7891), .DIN3(n7892), .Q(n7883) );
  nnd2s1 U8582 ( .DIN1(n623), .DIN2(n7404), .Q(n7892) );
  nnd2s1 U8583 ( .DIN1(n5876), .DIN2(n7414), .Q(n7891) );
  nnd2s1 U8584 ( .DIN1(n547), .DIN2(n7412), .Q(n7890) );
  nnd2s1 U8585 ( .DIN1(n630), .DIN2(n7884), .Q(n7888) );
  nnd2s1 U8586 ( .DIN1(n5994), .DIN2(n7893), .Q(n7886) );
  nnd2s1 U8587 ( .DIN1(n386), .DIN2(n6079), .Q(n7893) );
  and3s1 U8588 ( .DIN1(n7894), .DIN2(n7895), .DIN3(n801), .Q(n6079) );
  or2s1 U8589 ( .DIN1(n5654), .DIN2(n5490), .Q(n7894) );
  nnd2s1 U8590 ( .DIN1(n550), .DIN2(n7896), .Q(n7837) );
  nnd4s1 U8591 ( .DIN1(n7897), .DIN2(n7898), .DIN3(n7899), .DIN4(n7900), 
        .Q(n7896) );
  and3s1 U8592 ( .DIN1(n7901), .DIN2(n7902), .DIN3(n7903), .Q(n7900) );
  nnd2s1 U8593 ( .DIN1(n400), .DIN2(n6051), .Q(n7903) );
  nnd3s1 U8594 ( .DIN1(n7904), .DIN2(n7905), .DIN3(n7906), .Q(n6051) );
  nnd2s1 U8595 ( .DIN1(n554), .DIN2(n6479), .Q(n7906) );
  nnd4s1 U8596 ( .DIN1(n7907), .DIN2(n7908), .DIN3(n7909), .DIN4(n7910), 
        .Q(n6479) );
  nnd2s1 U8597 ( .DIN1(n784), .DIN2(n429), .Q(n7910) );
  nnd2s1 U8598 ( .DIN1(n759), .DIN2(n427), .Q(n7909) );
  nnd2s1 U8599 ( .DIN1(n5826), .DIN2(n7911), .Q(n7905) );
  nnd2s1 U8600 ( .DIN1(n545), .DIN2(n6911), .Q(n7904) );
  nnd4s1 U8601 ( .DIN1(n7912), .DIN2(n7913), .DIN3(n7914), .DIN4(n7915), 
        .Q(n7902) );
  and3s1 U8602 ( .DIN1(n7916), .DIN2(n7917), .DIN3(n730), .Q(n7915) );
  nnd2s1 U8603 ( .DIN1(n7918), .DIN2(n700), .Q(n7917) );
  nnd2s1 U8604 ( .DIN1(n6052), .DIN2(n805), .Q(n7916) );
  nnd3s1 U8605 ( .DIN1(n7919), .DIN2(n7920), .DIN3(n736), .Q(n6052) );
  nnd2s1 U8606 ( .DIN1(n7442), .DIN2(n792), .Q(n7920) );
  hi1s1 U8607 ( .DIN(n5569), .Q(n7442) );
  nnd2s1 U8608 ( .DIN1(n7438), .DIN2(n397), .Q(n7914) );
  nnd2s1 U8609 ( .DIN1(n7441), .DIN2(n5315), .Q(n7913) );
  nnd2s1 U8610 ( .DIN1(n7440), .DIN2(n5304), .Q(n7912) );
  nnd3s1 U8611 ( .DIN1(n7921), .DIN2(n7922), .DIN3(n7594), .Q(n7901) );
  nnd4s1 U8612 ( .DIN1(n7923), .DIN2(n7924), .DIN3(n733), .DIN4(n7925), 
        .Q(n7922) );
  and3s1 U8613 ( .DIN1(n7926), .DIN2(n7927), .DIN3(n7928), .Q(n7925) );
  nnd2s1 U8614 ( .DIN1(n719), .DIN2(n7454), .Q(n7928) );
  nnd2s1 U8615 ( .DIN1(n6032), .DIN2(n806), .Q(n7927) );
  nnd3s1 U8616 ( .DIN1(n7929), .DIN2(n5556), .DIN3(n7930), .Q(n6032) );
  nnd2s1 U8617 ( .DIN1(n555), .DIN2(n7452), .Q(n7930) );
  nnd2s1 U8618 ( .DIN1(n544), .DIN2(n5575), .Q(n7929) );
  nnd2s1 U8619 ( .DIN1(n5315), .DIN2(n7455), .Q(n7926) );
  nnd2s1 U8620 ( .DIN1(n398), .DIN2(n7456), .Q(n7924) );
  nnd2s1 U8621 ( .DIN1(n5306), .DIN2(n7931), .Q(n7923) );
  nnd2s1 U8622 ( .DIN1(n7605), .DIN2(n7932), .Q(n7921) );
  nnd3s1 U8623 ( .DIN1(n6379), .DIN2(n6034), .DIN3(n5321), .Q(n7932) );
  hi1s1 U8624 ( .DIN(n7007), .Q(n7605) );
  nnd2s1 U8625 ( .DIN1(n6898), .DIN2(n7933), .Q(n7007) );
  nnd2s1 U8626 ( .DIN1(n6896), .DIN2(reg_out_A[31]), .Q(n7933) );
  and2s1 U8627 ( .DIN1(n6379), .DIN2(n740), .Q(n6896) );
  nnd2s1 U8628 ( .DIN1(n7206), .DIN2(n75), .Q(n7899) );
  nnd2s1 U8629 ( .DIN1(n424), .DIN2(n7934), .Q(n7898) );
  nnd4s1 U8630 ( .DIN1(n7935), .DIN2(n7936), .DIN3(n7937), .DIN4(n7059), 
        .Q(n7934) );
  nnd2s1 U8631 ( .DIN1(n7938), .DIN2(n7212), .Q(n7937) );
  xnr2s1 U8632 ( .DIN1(n7803), .DIN2(n7804), .Q(n7938) );
  hi1s1 U8633 ( .DIN(n7939), .Q(n7804) );
  nnd2s1 U8634 ( .DIN1(n7940), .DIN2(n743), .Q(n7936) );
  xnr2s1 U8635 ( .DIN1(n7809), .DIN2(n7810), .Q(n7940) );
  hi1s1 U8636 ( .DIN(n7941), .Q(n7810) );
  nor2s1 U8637 ( .DIN1(n7942), .DIN2(n7943), .Q(n7935) );
  nor2s1 U8638 ( .DIN1(n75), .DIN2(n7006), .Q(n7943) );
  nor2s1 U8639 ( .DIN1(n9482), .DIN2(n7037), .Q(n7942) );
  nnd2s1 U8640 ( .DIN1(n7944), .DIN2(n66), .Q(n7897) );
  nnd3s1 U8641 ( .DIN1(n7945), .DIN2(n7946), .DIN3(n7947), .Q(n7944) );
  nnd2s1 U8642 ( .DIN1(n7222), .DIN2(n75), .Q(n7947) );
  nnd2s1 U8643 ( .DIN1(n7948), .DIN2(n722), .Q(n7946) );
  xnr2s1 U8644 ( .DIN1(n7803), .DIN2(n7939), .Q(n7948) );
  xnr2s1 U8645 ( .DIN1(n9482), .DIN2(n785), .Q(n7939) );
  nnd2s1 U8646 ( .DIN1(n7949), .DIN2(n7950), .Q(n7803) );
  nnd2s1 U8647 ( .DIN1(n36), .DIN2(n7951), .Q(n7950) );
  nnd2s1 U8648 ( .DIN1(n7952), .DIN2(n7953), .Q(n7951) );
  or2s1 U8649 ( .DIN1(n7953), .DIN2(n7952), .Q(n7949) );
  nnd2s1 U8650 ( .DIN1(n7954), .DIN2(n7058), .Q(n7945) );
  xnr2s1 U8651 ( .DIN1(n7809), .DIN2(n7941), .Q(n7954) );
  xnr2s1 U8652 ( .DIN1(n5423), .DIN2(n75), .Q(n7941) );
  nnd2s1 U8653 ( .DIN1(n7955), .DIN2(n7956), .Q(n7809) );
  nnd2s1 U8654 ( .DIN1(n425), .DIN2(n7957), .Q(n7956) );
  nnd2s1 U8655 ( .DIN1(n7958), .DIN2(n391), .Q(n7957) );
  or2s1 U8656 ( .DIN1(n391), .DIN2(n7958), .Q(n7955) );
  nnd3s1 U8657 ( .DIN1(n7959), .DIN2(n7960), .DIN3(n7961), .Q(\EXinst/n1440 )
         );
  nnd2s1 U8658 ( .DIN1(n5394), .DIN2(\DM_addr[8] ), .Q(n7961) );
  nnd2s1 U8659 ( .DIN1(n5324), .DIN2(n7962), .Q(n7960) );
  nnd4s1 U8660 ( .DIN1(n7963), .DIN2(n7964), .DIN3(n7965), .DIN4(n7966), 
        .Q(n7962) );
  and4s1 U8661 ( .DIN1(n7967), .DIN2(n7968), .DIN3(n7969), .DIN4(n7970), 
        .Q(n7966) );
  nnd2s1 U8662 ( .DIN1(n7971), .DIN2(n7972), .Q(n7970) );
  nnd3s1 U8663 ( .DIN1(n7973), .DIN2(n5372), .DIN3(n7974), .Q(n7971) );
  nnd2s1 U8664 ( .DIN1(n620), .DIN2(n7865), .Q(n7974) );
  nnd2s1 U8665 ( .DIN1(n656), .DIN2(n7860), .Q(n7973) );
  hi1s1 U8666 ( .DIN(n7861), .Q(n7860) );
  nnd2s1 U8667 ( .DIN1(n7975), .DIN2(n7976), .Q(n7969) );
  nnd2s1 U8668 ( .DIN1(n7977), .DIN2(n7978), .Q(n7976) );
  nnd2s1 U8669 ( .DIN1(n655), .DIN2(n7861), .Q(n7978) );
  nnd2s1 U8670 ( .DIN1(n7979), .DIN2(n7980), .Q(n7861) );
  nnd2s1 U8671 ( .DIN1(reg_out_B[7]), .DIN2(n7981), .Q(n7980) );
  nnd2s1 U8672 ( .DIN1(n7982), .DIN2(n63), .Q(n7981) );
  nnd2s1 U8673 ( .DIN1(n429), .DIN2(n7983), .Q(n7979) );
  or2s1 U8674 ( .DIN1(n7865), .DIN2(n5375), .Q(n7977) );
  nnd2s1 U8675 ( .DIN1(n7984), .DIN2(n7985), .Q(n7865) );
  nnd2s1 U8676 ( .DIN1(n7986), .DIN2(n7987), .Q(n7985) );
  nnd2s1 U8677 ( .DIN1(n7138), .DIN2(n6231), .Q(n7968) );
  nnd3s1 U8678 ( .DIN1(n7988), .DIN2(n7989), .DIN3(n7990), .Q(n6231) );
  nnd2s1 U8679 ( .DIN1(n629), .DIN2(n6652), .Q(n7990) );
  nnd4s1 U8680 ( .DIN1(n7991), .DIN2(n7992), .DIN3(n7993), .DIN4(n7994), 
        .Q(n6652) );
  nnd2s1 U8681 ( .DIN1(n7106), .DIN2(n547), .Q(n7989) );
  nnd2s1 U8682 ( .DIN1(n622), .DIN2(n7100), .Q(n7988) );
  nnd2s1 U8683 ( .DIN1(n36), .DIN2(n768), .Q(n7967) );
  nnd2s1 U8684 ( .DIN1(reg_out_B[8]), .DIN2(n7995), .Q(n7965) );
  nnd2s1 U8685 ( .DIN1(n5471), .DIN2(n7996), .Q(n7995) );
  nnd2s1 U8686 ( .DIN1(n775), .DIN2(n36), .Q(n7996) );
  nnd3s1 U8687 ( .DIN1(n7997), .DIN2(n7998), .DIN3(n7398), .Q(n7964) );
  nnd4s1 U8688 ( .DIN1(n7276), .DIN2(n7999), .DIN3(n8000), .DIN4(n8001), 
        .Q(n7998) );
  nnd2s1 U8689 ( .DIN1(n6210), .DIN2(n753), .Q(n8001) );
  nnd2s1 U8690 ( .DIN1(n8002), .DIN2(n808), .Q(n8000) );
  nnd2s1 U8691 ( .DIN1(n5345), .DIN2(n8003), .Q(n7999) );
  nnd2s1 U8692 ( .DIN1(n6723), .DIN2(n6301), .Q(n7997) );
  hi1s1 U8693 ( .DIN(n7156), .Q(n6301) );
  nor2s1 U8694 ( .DIN1(n5337), .DIN2(n807), .Q(n6723) );
  nnd2s1 U8695 ( .DIN1(n8004), .DIN2(n8005), .Q(n7963) );
  nnd3s1 U8696 ( .DIN1(n8006), .DIN2(n807), .DIN3(n8007), .Q(n8005) );
  hi1s1 U8697 ( .DIN(n8002), .Q(n8007) );
  nnd3s1 U8698 ( .DIN1(n8008), .DIN2(n8009), .DIN3(n8010), .Q(n8002) );
  nnd2s1 U8699 ( .DIN1(n621), .DIN2(n7526), .Q(n8010) );
  nnd2s1 U8700 ( .DIN1(n5876), .DIN2(n7537), .Q(n8009) );
  nnd2s1 U8701 ( .DIN1(n546), .DIN2(n7535), .Q(n8008) );
  nnd2s1 U8702 ( .DIN1(n630), .DIN2(n8003), .Q(n8006) );
  nnd2s1 U8703 ( .DIN1(n5994), .DIN2(n8011), .Q(n8004) );
  nnd2s1 U8704 ( .DIN1(n386), .DIN2(n6210), .Q(n8011) );
  and3s1 U8705 ( .DIN1(n8012), .DIN2(n8013), .DIN3(n801), .Q(n6210) );
  or2s1 U8706 ( .DIN1(n7536), .DIN2(n32), .Q(n8013) );
  nnd2s1 U8707 ( .DIN1(n8014), .DIN2(n32), .Q(n8012) );
  nnd2s1 U8708 ( .DIN1(n9453), .DIN2(n8015), .Q(n7959) );
  nnd4s1 U8709 ( .DIN1(n8016), .DIN2(n8017), .DIN3(n8018), .DIN4(n8019), 
        .Q(n8015) );
  and4s1 U8710 ( .DIN1(n8020), .DIN2(n8021), .DIN3(n8022), .DIN4(n8023), 
        .Q(n8019) );
  nnd2s1 U8711 ( .DIN1(n425), .DIN2(n8024), .Q(n8023) );
  nnd4s1 U8712 ( .DIN1(n8025), .DIN2(n8026), .DIN3(n8027), .DIN4(n7059), 
        .Q(n8024) );
  nnd2s1 U8713 ( .DIN1(n8028), .DIN2(n7212), .Q(n8027) );
  xnr2s1 U8714 ( .DIN1(n7953), .DIN2(n7952), .Q(n8028) );
  hi1s1 U8715 ( .DIN(n8029), .Q(n7952) );
  nnd2s1 U8716 ( .DIN1(n8030), .DIN2(n743), .Q(n8026) );
  xnr2s1 U8717 ( .DIN1(n391), .DIN2(n7958), .Q(n8030) );
  hi1s1 U8718 ( .DIN(n8031), .Q(n7958) );
  nnd2s1 U8719 ( .DIN1(n7314), .DIN2(n107), .Q(n8025) );
  nnd2s1 U8720 ( .DIN1(n8032), .DIN2(n332), .Q(n8022) );
  nnd2s1 U8721 ( .DIN1(n8033), .DIN2(n8034), .Q(n8032) );
  nnd2s1 U8722 ( .DIN1(n8035), .DIN2(n722), .Q(n8034) );
  xnr2s1 U8723 ( .DIN1(n8029), .DIN2(n7953), .Q(n8035) );
  xor2s1 U8724 ( .DIN1(n9483), .DIN2(n745), .Q(n7953) );
  nnd2s1 U8725 ( .DIN1(n8036), .DIN2(n8037), .Q(n8029) );
  nnd2s1 U8726 ( .DIN1(n429), .DIN2(n8038), .Q(n8037) );
  or2s1 U8727 ( .DIN1(n8039), .DIN2(n8040), .Q(n8038) );
  nnd2s1 U8728 ( .DIN1(n8040), .DIN2(n8039), .Q(n8036) );
  nnd2s1 U8729 ( .DIN1(n8041), .DIN2(n7058), .Q(n8033) );
  xnr2s1 U8730 ( .DIN1(n8031), .DIN2(n391), .Q(n8041) );
  nnd2s1 U8731 ( .DIN1(n8042), .DIN2(n8043), .Q(n8031) );
  nnd2s1 U8732 ( .DIN1(n429), .DIN2(n8044), .Q(n8043) );
  or2s1 U8733 ( .DIN1(n8045), .DIN2(n8046), .Q(n8044) );
  nnd2s1 U8734 ( .DIN1(n8046), .DIN2(n8045), .Q(n8042) );
  nnd2s1 U8735 ( .DIN1(n400), .DIN2(n6183), .Q(n8021) );
  nnd3s1 U8736 ( .DIN1(n8047), .DIN2(n8048), .DIN3(n8049), .Q(n6183) );
  nnd2s1 U8737 ( .DIN1(n554), .DIN2(n6608), .Q(n8049) );
  nnd4s1 U8738 ( .DIN1(n8050), .DIN2(n8051), .DIN3(n8052), .DIN4(n8053), 
        .Q(n6608) );
  nnd2s1 U8739 ( .DIN1(n759), .DIN2(n428), .Q(n8052) );
  nnd2s1 U8740 ( .DIN1(n7026), .DIN2(n726), .Q(n8048) );
  nnd2s1 U8741 ( .DIN1(n545), .DIN2(n7024), .Q(n8047) );
  nnd2s1 U8742 ( .DIN1(n7206), .DIN2(n107), .Q(n8020) );
  or2s1 U8743 ( .DIN1(n8054), .DIN2(n7006), .Q(n8018) );
  nnd4s1 U8744 ( .DIN1(n8055), .DIN2(n8056), .DIN3(n8057), .DIN4(n8058), 
        .Q(n8017) );
  and3s1 U8745 ( .DIN1(n8059), .DIN2(n8060), .DIN3(n730), .Q(n8058) );
  nnd2s1 U8746 ( .DIN1(n8061), .DIN2(n5306), .Q(n8060) );
  nnd2s1 U8747 ( .DIN1(n6232), .DIN2(n805), .Q(n8059) );
  nnd2s1 U8748 ( .DIN1(n7586), .DIN2(n398), .Q(n8057) );
  nnd2s1 U8749 ( .DIN1(n7590), .DIN2(n5315), .Q(n8056) );
  nnd2s1 U8750 ( .DIN1(n7588), .DIN2(n719), .Q(n8055) );
  hi1s1 U8751 ( .DIN(n7602), .Q(n7588) );
  nnd3s1 U8752 ( .DIN1(n8062), .DIN2(n8063), .DIN3(n7193), .Q(n8016) );
  nnd4s1 U8753 ( .DIN1(n8064), .DIN2(n8065), .DIN3(n9486), .DIN4(n8066), 
        .Q(n8062) );
  and3s1 U8754 ( .DIN1(n8067), .DIN2(n8068), .DIN3(n8069), .Q(n8066) );
  nnd2s1 U8755 ( .DIN1(n5304), .DIN2(n7602), .Q(n8069) );
  nnd2s1 U8756 ( .DIN1(n6167), .DIN2(n806), .Q(n8068) );
  nnd2s1 U8757 ( .DIN1(n5556), .DIN2(n6232), .Q(n6167) );
  nnd3s1 U8758 ( .DIN1(n8070), .DIN2(n8071), .DIN3(n736), .Q(n6232) );
  nnd2s1 U8759 ( .DIN1(n7591), .DIN2(n792), .Q(n8071) );
  nnd2s1 U8760 ( .DIN1(n7587), .DIN2(n29), .Q(n8070) );
  hi1s1 U8761 ( .DIN(n7601), .Q(n7587) );
  nnd2s1 U8762 ( .DIN1(n5315), .DIN2(n7603), .Q(n8067) );
  nnd2s1 U8763 ( .DIN1(n397), .DIN2(n7604), .Q(n8065) );
  nnd2s1 U8764 ( .DIN1(n5306), .DIN2(n8072), .Q(n8064) );
  nnd3s1 U8765 ( .DIN1(n8073), .DIN2(n8074), .DIN3(n8075), .Q(\EXinst/n1439 )
         );
  nnd2s1 U8766 ( .DIN1(n727), .DIN2(\DM_addr[7] ), .Q(n8075) );
  nnd2s1 U8767 ( .DIN1(n5324), .DIN2(n8076), .Q(n8074) );
  nnd4s1 U8768 ( .DIN1(n8077), .DIN2(n8078), .DIN3(n8079), .DIN4(n8080), 
        .Q(n8076) );
  and4s1 U8769 ( .DIN1(n8081), .DIN2(n8082), .DIN3(n8083), .DIN4(n8084), 
        .Q(n8080) );
  nnd2s1 U8770 ( .DIN1(n8085), .DIN2(n8086), .Q(n8084) );
  nnd3s1 U8771 ( .DIN1(n8087), .DIN2(n749), .DIN3(n8088), .Q(n8085) );
  nnd2s1 U8772 ( .DIN1(n705), .DIN2(n7986), .Q(n8088) );
  nnd2s1 U8773 ( .DIN1(n654), .DIN2(n7982), .Q(n8087) );
  hi1s1 U8774 ( .DIN(n7983), .Q(n7982) );
  nnd2s1 U8775 ( .DIN1(n8089), .DIN2(n8090), .Q(n8083) );
  nnd2s1 U8776 ( .DIN1(n8091), .DIN2(n8092), .Q(n8090) );
  nnd2s1 U8777 ( .DIN1(n653), .DIN2(n7983), .Q(n8092) );
  nnd2s1 U8778 ( .DIN1(n8093), .DIN2(n8094), .Q(n7983) );
  nnd2s1 U8779 ( .DIN1(reg_out_B[6]), .DIN2(n8095), .Q(n8094) );
  nnd2s1 U8780 ( .DIN1(n8096), .DIN2(n333), .Q(n8095) );
  nnd2s1 U8781 ( .DIN1(n427), .DIN2(n8097), .Q(n8093) );
  or2s1 U8782 ( .DIN1(n7986), .DIN2(n706), .Q(n8091) );
  nnd2s1 U8783 ( .DIN1(n8098), .DIN2(n8099), .Q(n7986) );
  nnd2s1 U8784 ( .DIN1(n8100), .DIN2(n8101), .Q(n8099) );
  nnd2s1 U8785 ( .DIN1(n7138), .DIN2(n6315), .Q(n8082) );
  and3s1 U8786 ( .DIN1(n8102), .DIN2(n8103), .DIN3(n801), .Q(n6315) );
  nnd2s1 U8787 ( .DIN1(n6738), .DIN2(n205), .Q(n8103) );
  hi1s1 U8788 ( .DIN(n7143), .Q(n6738) );
  nnd4s1 U8789 ( .DIN1(n8104), .DIN2(n8105), .DIN3(n8106), .DIN4(n8107), 
        .Q(n7143) );
  or2s1 U8790 ( .DIN1(n6745), .DIN2(n5490), .Q(n8102) );
  nnd2s1 U8791 ( .DIN1(n429), .DIN2(n767), .Q(n8081) );
  nnd2s1 U8792 ( .DIN1(reg_out_B[7]), .DIN2(n8108), .Q(n8079) );
  nnd2s1 U8793 ( .DIN1(n5471), .DIN2(n8109), .Q(n8108) );
  nnd2s1 U8794 ( .DIN1(n776), .DIN2(n429), .Q(n8109) );
  nnd3s1 U8795 ( .DIN1(n8110), .DIN2(n8111), .DIN3(n5336), .Q(n8078) );
  nnd2s1 U8796 ( .DIN1(n8112), .DIN2(n6300), .Q(n8111) );
  hi1s1 U8797 ( .DIN(n5362), .Q(n6300) );
  nnd4s1 U8798 ( .DIN1(n7276), .DIN2(n8113), .DIN3(n8114), .DIN4(n8115), 
        .Q(n8110) );
  nnd2s1 U8799 ( .DIN1(n752), .DIN2(n8116), .Q(n8115) );
  nnd2s1 U8800 ( .DIN1(n8117), .DIN2(n204), .Q(n8114) );
  nnd2s1 U8801 ( .DIN1(n5345), .DIN2(n8118), .Q(n8113) );
  and2s1 U8802 ( .DIN1(n5337), .DIN2(n8119), .Q(n7276) );
  nnd2s1 U8803 ( .DIN1(n6216), .DIN2(n55), .Q(n8119) );
  nnd2s1 U8804 ( .DIN1(n8120), .DIN2(n8121), .Q(n8077) );
  nnd3s1 U8805 ( .DIN1(n8122), .DIN2(n807), .DIN3(n8123), .Q(n8121) );
  hi1s1 U8806 ( .DIN(n8117), .Q(n8123) );
  nnd3s1 U8807 ( .DIN1(n8124), .DIN2(n8125), .DIN3(n8126), .Q(n8117) );
  nnd2s1 U8808 ( .DIN1(n623), .DIN2(n7651), .Q(n8126) );
  nnd2s1 U8809 ( .DIN1(n5876), .DIN2(n6728), .Q(n8125) );
  nnd2s1 U8810 ( .DIN1(n547), .DIN2(n7163), .Q(n8124) );
  nnd2s1 U8811 ( .DIN1(n629), .DIN2(n8118), .Q(n8122) );
  nnd2s1 U8812 ( .DIN1(n5994), .DIN2(n8127), .Q(n8120) );
  nnd2s1 U8813 ( .DIN1(n386), .DIN2(n6288), .Q(n8127) );
  nnd2s1 U8814 ( .DIN1(n8128), .DIN2(n8129), .Q(n6288) );
  nnd2s1 U8815 ( .DIN1(n5362), .DIN2(n438), .Q(n8129) );
  nor2s1 U8816 ( .DIN1(n6863), .DIN2(n5353), .Q(n5362) );
  hi1s1 U8817 ( .DIN(n8116), .Q(n8128) );
  nnd2s1 U8818 ( .DIN1(n8130), .DIN2(n8131), .Q(n8116) );
  nnd2s1 U8819 ( .DIN1(n622), .DIN2(n5863), .Q(n8131) );
  nnd2s1 U8820 ( .DIN1(n630), .DIN2(n6729), .Q(n8130) );
  nnd2s1 U8821 ( .DIN1(n551), .DIN2(n8132), .Q(n8073) );
  nnd4s1 U8822 ( .DIN1(n8133), .DIN2(n8134), .DIN3(n8135), .DIN4(n8136), 
        .Q(n8132) );
  and3s1 U8823 ( .DIN1(n8137), .DIN2(n8138), .DIN3(n8139), .Q(n8136) );
  nnd2s1 U8824 ( .DIN1(n400), .DIN2(n6260), .Q(n8139) );
  and3s1 U8825 ( .DIN1(n8140), .DIN2(n8141), .DIN3(n736), .Q(n6260) );
  or2s1 U8826 ( .DIN1(n6689), .DIN2(n29), .Q(n8141) );
  or2s1 U8827 ( .DIN1(n6686), .DIN2(n792), .Q(n8140) );
  nnd4s1 U8828 ( .DIN1(n8142), .DIN2(n8143), .DIN3(n8144), .DIN4(n8145), 
        .Q(n6686) );
  nnd2s1 U8829 ( .DIN1(n783), .DIN2(n428), .Q(n8145) );
  nnd2s1 U8830 ( .DIN1(n758), .DIN2(n433), .Q(n8144) );
  nnd4s1 U8831 ( .DIN1(n8146), .DIN2(n8147), .DIN3(n7339), .DIN4(n8148), 
        .Q(n8138) );
  and3s1 U8832 ( .DIN1(n8149), .DIN2(n8150), .DIN3(n8151), .Q(n8148) );
  nnd2s1 U8833 ( .DIN1(n7189), .DIN2(n5304), .Q(n8151) );
  nnd3s1 U8834 ( .DIN1(n8152), .DIN2(n8153), .DIN3(n5306), .Q(n8150) );
  nnd2s1 U8835 ( .DIN1(n8154), .DIN2(n712), .Q(n8152) );
  nnd2s1 U8836 ( .DIN1(n7204), .DIN2(n5315), .Q(n8149) );
  nnd2s1 U8837 ( .DIN1(n7684), .DIN2(n397), .Q(n8147) );
  or2s1 U8838 ( .DIN1(n6261), .DIN2(n740), .Q(n8146) );
  nnd2s1 U8839 ( .DIN1(n8155), .DIN2(n8156), .Q(n6261) );
  nnd2s1 U8840 ( .DIN1(n5317), .DIN2(n735), .Q(n8156) );
  nnd3s1 U8841 ( .DIN1(n8157), .DIN2(n8158), .DIN3(n7193), .Q(n8137) );
  nnd4s1 U8842 ( .DIN1(n8159), .DIN2(n8160), .DIN3(n733), .DIN4(n8161), 
        .Q(n8158) );
  and3s1 U8843 ( .DIN1(n8162), .DIN2(n8163), .DIN3(n8164), .Q(n8161) );
  nnd2s1 U8844 ( .DIN1(n5315), .DIN2(n7696), .Q(n8164) );
  nnd2s1 U8845 ( .DIN1(n5306), .DIN2(n8165), .Q(n8163) );
  nnd2s1 U8846 ( .DIN1(n8166), .DIN2(n8142), .Q(n8165) );
  nnd2s1 U8847 ( .DIN1(n552), .DIN2(n429), .Q(n8142) );
  nnd2s1 U8848 ( .DIN1(n6244), .DIN2(n805), .Q(n8162) );
  nnd2s1 U8849 ( .DIN1(n8155), .DIN2(n5556), .Q(n6244) );
  hi1s1 U8850 ( .DIN(n8167), .Q(n5556) );
  and2s1 U8851 ( .DIN1(n8168), .DIN2(n8169), .Q(n8155) );
  nnd2s1 U8852 ( .DIN1(n544), .DIN2(n5807), .Q(n8169) );
  nnd2s1 U8853 ( .DIN1(n555), .DIN2(n7203), .Q(n8168) );
  nnd2s1 U8854 ( .DIN1(n719), .DIN2(n7693), .Q(n8160) );
  nnd2s1 U8855 ( .DIN1(n398), .DIN2(n7697), .Q(n8159) );
  nnd2s1 U8856 ( .DIN1(n8170), .DIN2(n7190), .Q(n8157) );
  hi1s1 U8857 ( .DIN(n5317), .Q(n7190) );
  nor2s1 U8858 ( .DIN1(n5741), .DIN2(n213), .Q(n5317) );
  nnd2s1 U8859 ( .DIN1(n7206), .DIN2(n76), .Q(n8135) );
  nnd2s1 U8860 ( .DIN1(n429), .DIN2(n8171), .Q(n8134) );
  nnd4s1 U8861 ( .DIN1(n7059), .DIN2(n8173), .DIN3(n8174), .DIN4(n8172), 
        .Q(n8171) );
  nnd2s1 U8862 ( .DIN1(n8175), .DIN2(n7212), .Q(n8174) );
  xnr2s1 U8863 ( .DIN1(n8039), .DIN2(n8040), .Q(n8175) );
  hi1s1 U8864 ( .DIN(n8176), .Q(n8040) );
  nnd2s1 U8865 ( .DIN1(n8177), .DIN2(n743), .Q(n8173) );
  xnr2s1 U8866 ( .DIN1(n8045), .DIN2(n8046), .Q(n8177) );
  hi1s1 U8867 ( .DIN(n8178), .Q(n8046) );
  nor2s1 U8868 ( .DIN1(n8179), .DIN2(n8180), .Q(n8172) );
  nor2s1 U8869 ( .DIN1(n76), .DIN2(n7006), .Q(n8180) );
  nor2s1 U8870 ( .DIN1(n9484), .DIN2(n7037), .Q(n8179) );
  nnd2s1 U8871 ( .DIN1(n8181), .DIN2(n63), .Q(n8133) );
  nnd3s1 U8872 ( .DIN1(n8182), .DIN2(n8183), .DIN3(n8184), .Q(n8181) );
  nnd2s1 U8873 ( .DIN1(n7222), .DIN2(n76), .Q(n8184) );
  nnd2s1 U8874 ( .DIN1(n8185), .DIN2(n722), .Q(n8183) );
  xnr2s1 U8875 ( .DIN1(n8039), .DIN2(n8176), .Q(n8185) );
  xnr2s1 U8876 ( .DIN1(n9484), .DIN2(n787), .Q(n8176) );
  nnd2s1 U8877 ( .DIN1(n8186), .DIN2(n8187), .Q(n8039) );
  nnd2s1 U8878 ( .DIN1(n34), .DIN2(n8188), .Q(n8187) );
  nnd2s1 U8879 ( .DIN1(n8189), .DIN2(n8190), .Q(n8188) );
  or2s1 U8880 ( .DIN1(n8190), .DIN2(n8189), .Q(n8186) );
  nnd2s1 U8881 ( .DIN1(n8191), .DIN2(n7058), .Q(n8182) );
  xnr2s1 U8882 ( .DIN1(n8045), .DIN2(n8178), .Q(n8191) );
  xnr2s1 U8883 ( .DIN1(n633), .DIN2(n76), .Q(n8178) );
  nnd2s1 U8884 ( .DIN1(n8192), .DIN2(n8193), .Q(n8045) );
  nnd2s1 U8885 ( .DIN1(n427), .DIN2(n8194), .Q(n8193) );
  nnd2s1 U8886 ( .DIN1(n8195), .DIN2(n392), .Q(n8194) );
  or2s1 U8887 ( .DIN1(n392), .DIN2(n8195), .Q(n8192) );
  nnd3s1 U8888 ( .DIN1(n8196), .DIN2(n8197), .DIN3(n8198), .Q(\EXinst/n1438 )
         );
  nnd2s1 U8889 ( .DIN1(n5394), .DIN2(\DM_addr[6] ), .Q(n8198) );
  nnd2s1 U8890 ( .DIN1(n5324), .DIN2(n8199), .Q(n8197) );
  nnd4s1 U8891 ( .DIN1(n8200), .DIN2(n8201), .DIN3(n8202), .DIN4(n8203), 
        .Q(n8199) );
  and4s1 U8892 ( .DIN1(n8204), .DIN2(n8205), .DIN3(n8206), .DIN4(n8207), 
        .Q(n8203) );
  nnd2s1 U8893 ( .DIN1(n8208), .DIN2(n8209), .Q(n8207) );
  nnd3s1 U8894 ( .DIN1(n8210), .DIN2(n5372), .DIN3(n8211), .Q(n8208) );
  nnd2s1 U8895 ( .DIN1(n620), .DIN2(n8101), .Q(n8211) );
  nnd2s1 U8896 ( .DIN1(n656), .DIN2(n8096), .Q(n8210) );
  hi1s1 U8897 ( .DIN(n8097), .Q(n8096) );
  nnd2s1 U8898 ( .DIN1(n8212), .DIN2(n8213), .Q(n8206) );
  nnd2s1 U8899 ( .DIN1(n8214), .DIN2(n8215), .Q(n8213) );
  nnd2s1 U8900 ( .DIN1(n655), .DIN2(n8097), .Q(n8215) );
  nnd2s1 U8901 ( .DIN1(n8216), .DIN2(n8217), .Q(n8097) );
  nnd2s1 U8902 ( .DIN1(n716), .DIN2(n8218), .Q(n8217) );
  nnd2s1 U8903 ( .DIN1(n8219), .DIN2(n81), .Q(n8218) );
  nnd2s1 U8904 ( .DIN1(n428), .DIN2(n8220), .Q(n8216) );
  or2s1 U8905 ( .DIN1(n8101), .DIN2(n5375), .Q(n8214) );
  nnd2s1 U8906 ( .DIN1(n8221), .DIN2(n8222), .Q(n8101) );
  nnd2s1 U8907 ( .DIN1(n8223), .DIN2(n8224), .Q(n8222) );
  nnd2s1 U8908 ( .DIN1(n7138), .DIN2(n6451), .Q(n8205) );
  and3s1 U8909 ( .DIN1(n8225), .DIN2(n8226), .DIN3(n801), .Q(n6451) );
  nnd2s1 U8910 ( .DIN1(n6873), .DIN2(n205), .Q(n8226) );
  hi1s1 U8911 ( .DIN(n7267), .Q(n6873) );
  nnd4s1 U8912 ( .DIN1(n8227), .DIN2(n8228), .DIN3(n8229), .DIN4(n8230), 
        .Q(n7267) );
  nnd2s1 U8913 ( .DIN1(n531), .DIN2(n431), .Q(n8229) );
  or2s1 U8914 ( .DIN1(n6879), .DIN2(n205), .Q(n8225) );
  nnd2s1 U8915 ( .DIN1(n34), .DIN2(n768), .Q(n8204) );
  nnd2s1 U8916 ( .DIN1(reg_out_B[6]), .DIN2(n8231), .Q(n8202) );
  nnd2s1 U8917 ( .DIN1(n5471), .DIN2(n8232), .Q(n8231) );
  nnd2s1 U8918 ( .DIN1(n775), .DIN2(n34), .Q(n8232) );
  nnd3s1 U8919 ( .DIN1(n8233), .DIN2(n8234), .DIN3(n769), .Q(n8201) );
  nnd4s1 U8920 ( .DIN1(n8235), .DIN2(n5337), .DIN3(n8236), .DIN4(n8237), 
        .Q(n8233) );
  nnd2s1 U8921 ( .DIN1(n752), .DIN2(n6435), .Q(n8237) );
  nnd2s1 U8922 ( .DIN1(n8238), .DIN2(n8239), .Q(n6435) );
  nnd2s1 U8923 ( .DIN1(n438), .DIN2(n5477), .Q(n8239) );
  nnd3s1 U8924 ( .DIN1(n8240), .DIN2(n8241), .DIN3(n8242), .Q(n5477) );
  nnd2s1 U8925 ( .DIN1(n734), .DIN2(n5353), .Q(n8242) );
  hi1s1 U8926 ( .DIN(n8243), .Q(n8241) );
  nnd2s1 U8927 ( .DIN1(n5495), .DIN2(n205), .Q(n8240) );
  nnd2s1 U8928 ( .DIN1(n8244), .DIN2(n808), .Q(n8236) );
  nnd2s1 U8929 ( .DIN1(n5345), .DIN2(n8245), .Q(n8235) );
  nnd2s1 U8930 ( .DIN1(n8246), .DIN2(n8247), .Q(n8200) );
  nnd3s1 U8931 ( .DIN1(n8248), .DIN2(n807), .DIN3(n8249), .Q(n8247) );
  hi1s1 U8932 ( .DIN(n8244), .Q(n8249) );
  nnd3s1 U8933 ( .DIN1(n8250), .DIN2(n8251), .DIN3(n8252), .Q(n8244) );
  nnd2s1 U8934 ( .DIN1(n621), .DIN2(n7770), .Q(n8252) );
  nnd2s1 U8935 ( .DIN1(n5876), .DIN2(n7291), .Q(n8251) );
  nnd2s1 U8936 ( .DIN1(n546), .DIN2(n7281), .Q(n8250) );
  nnd2s1 U8937 ( .DIN1(n628), .DIN2(n8245), .Q(n8248) );
  nnd2s1 U8938 ( .DIN1(n5994), .DIN2(n8253), .Q(n8246) );
  nnd2s1 U8939 ( .DIN1(n386), .DIN2(n6428), .Q(n8253) );
  nnd3s1 U8940 ( .DIN1(n8254), .DIN2(n8255), .DIN3(n8238), .Q(n6428) );
  and2s1 U8941 ( .DIN1(n8256), .DIN2(n8257), .Q(n8238) );
  nnd2s1 U8942 ( .DIN1(n623), .DIN2(n7292), .Q(n8257) );
  nnd2s1 U8943 ( .DIN1(n628), .DIN2(n7293), .Q(n8256) );
  nnd3s1 U8944 ( .DIN1(n773), .DIN2(n5490), .DIN3(n6216), .Q(n8255) );
  nor2s1 U8945 ( .DIN1(n801), .DIN2(n401), .Q(n6216) );
  nnd2s1 U8946 ( .DIN1(n5495), .DIN2(n546), .Q(n8254) );
  nnd2s1 U8947 ( .DIN1(n550), .DIN2(n8258), .Q(n8196) );
  nnd4s1 U8948 ( .DIN1(n8259), .DIN2(n8260), .DIN3(n8261), .DIN4(n8262), 
        .Q(n8258) );
  and4s1 U8949 ( .DIN1(n8263), .DIN2(n8264), .DIN3(n8265), .DIN4(n8266), 
        .Q(n8262) );
  nnd2s1 U8950 ( .DIN1(n427), .DIN2(n8267), .Q(n8266) );
  nnd4s1 U8951 ( .DIN1(n8268), .DIN2(n8269), .DIN3(n8270), .DIN4(n7059), 
        .Q(n8267) );
  nnd2s1 U8952 ( .DIN1(n8271), .DIN2(n7212), .Q(n8270) );
  xnr2s1 U8953 ( .DIN1(n8190), .DIN2(n8189), .Q(n8271) );
  hi1s1 U8954 ( .DIN(n8272), .Q(n8189) );
  nnd2s1 U8955 ( .DIN1(n8273), .DIN2(n743), .Q(n8269) );
  xnr2s1 U8956 ( .DIN1(n392), .DIN2(n8195), .Q(n8273) );
  hi1s1 U8957 ( .DIN(n8274), .Q(n8195) );
  nnd2s1 U8958 ( .DIN1(n7314), .DIN2(n105), .Q(n8268) );
  nnd2s1 U8959 ( .DIN1(n8275), .DIN2(n333), .Q(n8265) );
  nnd2s1 U8960 ( .DIN1(n8276), .DIN2(n8277), .Q(n8275) );
  nnd2s1 U8961 ( .DIN1(n8278), .DIN2(n722), .Q(n8277) );
  xnr2s1 U8962 ( .DIN1(n8272), .DIN2(n8190), .Q(n8278) );
  xor2s1 U8963 ( .DIN1(n9485), .DIN2(n744), .Q(n8190) );
  nnd2s1 U8964 ( .DIN1(n8279), .DIN2(n8280), .Q(n8272) );
  nnd2s1 U8965 ( .DIN1(n428), .DIN2(n8281), .Q(n8280) );
  or2s1 U8966 ( .DIN1(n8282), .DIN2(n8283), .Q(n8281) );
  nnd2s1 U8967 ( .DIN1(n8283), .DIN2(n8282), .Q(n8279) );
  nnd2s1 U8968 ( .DIN1(n8284), .DIN2(n7058), .Q(n8276) );
  xnr2s1 U8969 ( .DIN1(n8274), .DIN2(n392), .Q(n8284) );
  nnd2s1 U8970 ( .DIN1(n8285), .DIN2(n8286), .Q(n8274) );
  nnd2s1 U8971 ( .DIN1(n428), .DIN2(n8287), .Q(n8286) );
  or2s1 U8972 ( .DIN1(n8288), .DIN2(n8289), .Q(n8287) );
  nnd2s1 U8973 ( .DIN1(n8289), .DIN2(n8288), .Q(n8285) );
  nnd2s1 U8974 ( .DIN1(n400), .DIN2(n6401), .Q(n8264) );
  and3s1 U8975 ( .DIN1(n8290), .DIN2(n8291), .DIN3(n736), .Q(n6401) );
  or2s1 U8976 ( .DIN1(n6830), .DIN2(n747), .Q(n8291) );
  or2s1 U8977 ( .DIN1(n6828), .DIN2(n792), .Q(n8290) );
  nnd4s1 U8978 ( .DIN1(n8292), .DIN2(n8293), .DIN3(n8294), .DIN4(n8295), 
        .Q(n6828) );
  nnd2s1 U8979 ( .DIN1(n784), .DIN2(n10), .Q(n8295) );
  nnd2s1 U8980 ( .DIN1(n759), .DIN2(n431), .Q(n8294) );
  nnd2s1 U8981 ( .DIN1(n7206), .DIN2(n105), .Q(n8263) );
  or2s1 U8982 ( .DIN1(n8296), .DIN2(n7006), .Q(n8261) );
  nnd4s1 U8983 ( .DIN1(n8297), .DIN2(n8298), .DIN3(n7339), .DIN4(n8299), 
        .Q(n8260) );
  and3s1 U8984 ( .DIN1(n8300), .DIN2(n8301), .DIN3(n8302), .Q(n8299) );
  nnd2s1 U8985 ( .DIN1(n7356), .DIN2(n719), .Q(n8302) );
  nnd3s1 U8986 ( .DIN1(n8303), .DIN2(n8304), .DIN3(n5306), .Q(n8301) );
  nnd3s1 U8987 ( .DIN1(n8305), .DIN2(n8306), .DIN3(n712), .Q(n8303) );
  nnd2s1 U8988 ( .DIN1(n9489), .DIN2(n333), .Q(n8306) );
  nnd2s1 U8989 ( .DIN1(n439), .DIN2(n63), .Q(n8305) );
  nnd2s1 U8990 ( .DIN1(n7357), .DIN2(n5315), .Q(n8300) );
  nnd2s1 U8991 ( .DIN1(n7834), .DIN2(n398), .Q(n8298) );
  nnd2s1 U8992 ( .DIN1(n6452), .DIN2(n806), .Q(n8297) );
  and3s1 U8993 ( .DIN1(n8307), .DIN2(n8308), .DIN3(n8309), .Q(n6452) );
  nnd3s1 U8994 ( .DIN1(n789), .DIN2(n29), .DIN3(n8167), .Q(n8308) );
  nor2s1 U8995 ( .DIN1(n401), .DIN2(n9487), .Q(n8167) );
  nnd2s1 U8996 ( .DIN1(n5546), .DIN2(n726), .Q(n8307) );
  nnd3s1 U8997 ( .DIN1(n8310), .DIN2(n8311), .DIN3(n8312), .Q(n8259) );
  nnd4s1 U8998 ( .DIN1(n8313), .DIN2(n8314), .DIN3(n733), .DIN4(n8315), 
        .Q(n8310) );
  and3s1 U8999 ( .DIN1(n8316), .DIN2(n8317), .DIN3(n8318), .Q(n8315) );
  nnd2s1 U9000 ( .DIN1(n5315), .DIN2(n8319), .Q(n8318) );
  nnd2s1 U9001 ( .DIN1(n8320), .DIN2(n805), .Q(n8317) );
  nnd2s1 U9002 ( .DIN1(n8309), .DIN2(n8321), .Q(n8320) );
  nnd2s1 U9003 ( .DIN1(n5557), .DIN2(n803), .Q(n8321) );
  nnd3s1 U9004 ( .DIN1(n8322), .DIN2(n8323), .DIN3(n8324), .Q(n5557) );
  nnd2s1 U9005 ( .DIN1(n734), .DIN2(n213), .Q(n8324) );
  hi1s1 U9006 ( .DIN(n8325), .Q(n8323) );
  nnd2s1 U9007 ( .DIN1(n5546), .DIN2(n747), .Q(n8322) );
  and2s1 U9008 ( .DIN1(n8326), .DIN2(n8327), .Q(n8309) );
  nnd2s1 U9009 ( .DIN1(n545), .DIN2(n7355), .Q(n8327) );
  nnd2s1 U9010 ( .DIN1(n554), .DIN2(n8328), .Q(n8326) );
  nnd2s1 U9011 ( .DIN1(n5306), .DIN2(n8329), .Q(n8316) );
  nnd3s1 U9012 ( .DIN1(n8051), .DIN2(n8304), .DIN3(n8292), .Q(n8329) );
  nnd2s1 U9013 ( .DIN1(n553), .DIN2(n427), .Q(n8292) );
  nnd2s1 U9014 ( .DIN1(n790), .DIN2(n429), .Q(n8051) );
  nnd2s1 U9015 ( .DIN1(n5304), .DIN2(n8330), .Q(n8314) );
  nnd2s1 U9016 ( .DIN1(n397), .DIN2(n8331), .Q(n8313) );
  nnd3s1 U9017 ( .DIN1(n8332), .DIN2(n8333), .DIN3(n8334), .Q(\EXinst/n1437 )
         );
  nnd2s1 U9018 ( .DIN1(n727), .DIN2(\DM_addr[5] ), .Q(n8334) );
  nnd2s1 U9019 ( .DIN1(n5324), .DIN2(n8335), .Q(n8333) );
  nnd4s1 U9020 ( .DIN1(n8336), .DIN2(n8337), .DIN3(n8338), .DIN4(n8339), 
        .Q(n8335) );
  and4s1 U9021 ( .DIN1(n8340), .DIN2(n8341), .DIN3(n8342), .DIN4(n8343), 
        .Q(n8339) );
  nnd2s1 U9022 ( .DIN1(n8344), .DIN2(n8345), .Q(n8343) );
  nnd3s1 U9023 ( .DIN1(n8346), .DIN2(n749), .DIN3(n8347), .Q(n8344) );
  nnd2s1 U9024 ( .DIN1(n705), .DIN2(n8223), .Q(n8347) );
  nnd2s1 U9025 ( .DIN1(n654), .DIN2(n8219), .Q(n8346) );
  hi1s1 U9026 ( .DIN(n8220), .Q(n8219) );
  nnd2s1 U9027 ( .DIN1(n8348), .DIN2(n8349), .Q(n8342) );
  nnd2s1 U9028 ( .DIN1(n8350), .DIN2(n8351), .Q(n8349) );
  nnd2s1 U9029 ( .DIN1(n653), .DIN2(n8220), .Q(n8351) );
  nnd2s1 U9030 ( .DIN1(n8352), .DIN2(n8353), .Q(n8220) );
  nnd2s1 U9031 ( .DIN1(n753), .DIN2(n8354), .Q(n8353) );
  nnd2s1 U9032 ( .DIN1(n8355), .DIN2(n334), .Q(n8354) );
  nnd2s1 U9033 ( .DIN1(n10), .DIN2(n8356), .Q(n8352) );
  or2s1 U9034 ( .DIN1(n8223), .DIN2(n5375), .Q(n8350) );
  nnd2s1 U9035 ( .DIN1(n8357), .DIN2(n8358), .Q(n8223) );
  nnd2s1 U9036 ( .DIN1(n8359), .DIN2(n8360), .Q(n8358) );
  nnd2s1 U9037 ( .DIN1(n716), .DIN2(n8361), .Q(n8341) );
  nnd2s1 U9038 ( .DIN1(n5471), .DIN2(n8362), .Q(n8361) );
  nnd2s1 U9039 ( .DIN1(n776), .DIN2(n428), .Q(n8362) );
  nnd2s1 U9040 ( .DIN1(n428), .DIN2(n767), .Q(n8340) );
  nnd2s1 U9041 ( .DIN1(n8363), .DIN2(n8364), .Q(n8338) );
  nnd3s1 U9042 ( .DIN1(n8365), .DIN2(n807), .DIN3(n8366), .Q(n8364) );
  hi1s1 U9043 ( .DIN(n8367), .Q(n8366) );
  nnd2s1 U9044 ( .DIN1(n628), .DIN2(n8368), .Q(n8365) );
  nnd2s1 U9045 ( .DIN1(n5994), .DIN2(n8369), .Q(n8363) );
  nnd2s1 U9046 ( .DIN1(n386), .DIN2(n6509), .Q(n8369) );
  nnd2s1 U9047 ( .DIN1(n8370), .DIN2(n8371), .Q(n6509) );
  nnd2s1 U9048 ( .DIN1(n547), .DIN2(n5654), .Q(n8371) );
  nnd3s1 U9049 ( .DIN1(n6530), .DIN2(n801), .DIN3(n7138), .Q(n8337) );
  nnd2s1 U9050 ( .DIN1(n8372), .DIN2(n8373), .Q(n6530) );
  nnd2s1 U9051 ( .DIN1(n6957), .DIN2(n205), .Q(n8373) );
  nnd4s1 U9052 ( .DIN1(n8374), .DIN2(n8375), .DIN3(n8376), .DIN4(n8377), 
        .Q(n6957) );
  nnd2s1 U9053 ( .DIN1(n532), .DIN2(n426), .Q(n8376) );
  nnd2s1 U9054 ( .DIN1(n741), .DIN2(n7873), .Q(n8372) );
  nnd2s1 U9055 ( .DIN1(n8378), .DIN2(n8379), .Q(n7873) );
  nnd2s1 U9056 ( .DIN1(n774), .DIN2(n33), .Q(n8379) );
  nnd3s1 U9057 ( .DIN1(n8380), .DIN2(n8381), .DIN3(n5336), .Q(n8336) );
  nnd2s1 U9058 ( .DIN1(n8382), .DIN2(n8383), .Q(n8381) );
  nnd2s1 U9059 ( .DIN1(n7283), .DIN2(n1), .Q(n8383) );
  hi1s1 U9060 ( .DIN(n8234), .Q(n8382) );
  nnd2s1 U9061 ( .DIN1(n8112), .DIN2(n8384), .Q(n8234) );
  nnd2s1 U9062 ( .DIN1(n7283), .DIN2(n714), .Q(n8384) );
  nnd4s1 U9063 ( .DIN1(n8385), .DIN2(n5337), .DIN3(n8386), .DIN4(n8387), 
        .Q(n8380) );
  nnd2s1 U9064 ( .DIN1(n753), .DIN2(n6516), .Q(n8387) );
  nnd2s1 U9065 ( .DIN1(n8370), .DIN2(n8388), .Q(n6516) );
  nnd2s1 U9066 ( .DIN1(n8389), .DIN2(n8390), .Q(n8388) );
  nnd2s1 U9067 ( .DIN1(n8391), .DIN2(n205), .Q(n8390) );
  and2s1 U9068 ( .DIN1(n8392), .DIN2(n8393), .Q(n8370) );
  nnd2s1 U9069 ( .DIN1(n622), .DIN2(n7413), .Q(n8393) );
  nnd2s1 U9070 ( .DIN1(n628), .DIN2(n7414), .Q(n8392) );
  nnd2s1 U9071 ( .DIN1(n8367), .DIN2(n204), .Q(n8386) );
  nnd3s1 U9072 ( .DIN1(n8394), .DIN2(n8395), .DIN3(n8396), .Q(n8367) );
  nnd2s1 U9073 ( .DIN1(n621), .DIN2(n7884), .Q(n8396) );
  nnd2s1 U9074 ( .DIN1(n5876), .DIN2(n7412), .Q(n8395) );
  nnd2s1 U9075 ( .DIN1(n546), .DIN2(n7404), .Q(n8394) );
  nnd2s1 U9076 ( .DIN1(n5345), .DIN2(n8368), .Q(n8385) );
  nnd2s1 U9077 ( .DIN1(n551), .DIN2(n8397), .Q(n8332) );
  nnd4s1 U9078 ( .DIN1(n8398), .DIN2(n8399), .DIN3(n8400), .DIN4(n8401), 
        .Q(n8397) );
  and3s1 U9079 ( .DIN1(n8402), .DIN2(n8403), .DIN3(n8404), .Q(n8401) );
  nnd3s1 U9080 ( .DIN1(n9487), .DIN2(n6481), .DIN3(n400), .Q(n8404) );
  nnd2s1 U9081 ( .DIN1(n8405), .DIN2(n8406), .Q(n6481) );
  nnd2s1 U9082 ( .DIN1(n29), .DIN2(n6911), .Q(n8406) );
  nnd4s1 U9083 ( .DIN1(n8407), .DIN2(n8408), .DIN3(n8409), .DIN4(n8410), 
        .Q(n6911) );
  nnd2s1 U9084 ( .DIN1(n783), .DIN2(n431), .Q(n8410) );
  nnd2s1 U9085 ( .DIN1(n759), .DIN2(n426), .Q(n8409) );
  nnd2s1 U9086 ( .DIN1(n789), .DIN2(n433), .Q(n8408) );
  nnd2s1 U9087 ( .DIN1(n7911), .DIN2(n792), .Q(n8405) );
  nnd2s1 U9088 ( .DIN1(n8411), .DIN2(n8412), .Q(n7911) );
  nnd2s1 U9089 ( .DIN1(n790), .DIN2(n430), .Q(n8412) );
  nnd2s1 U9090 ( .DIN1(n552), .DIN2(n35), .Q(n8411) );
  nnd4s1 U9091 ( .DIN1(n8413), .DIN2(n8414), .DIN3(n7339), .DIN4(n8415), 
        .Q(n8403) );
  and3s1 U9092 ( .DIN1(n8416), .DIN2(n8417), .DIN3(n8418), .Q(n8415) );
  nnd2s1 U9093 ( .DIN1(n7441), .DIN2(n5304), .Q(n8418) );
  nnd3s1 U9094 ( .DIN1(n8419), .DIN2(n8420), .DIN3(n5306), .Q(n8417) );
  nnd3s1 U9095 ( .DIN1(n8421), .DIN2(n8422), .DIN3(n712), .Q(n8419) );
  nnd2s1 U9096 ( .DIN1(n9489), .DIN2(n81), .Q(n8422) );
  nnd2s1 U9097 ( .DIN1(n440), .DIN2(n333), .Q(n8421) );
  nnd2s1 U9098 ( .DIN1(n7438), .DIN2(n5315), .Q(n8416) );
  nnd2s1 U9099 ( .DIN1(n7918), .DIN2(n397), .Q(n8414) );
  or2s1 U9100 ( .DIN1(n6482), .DIN2(n739), .Q(n8413) );
  nnd2s1 U9101 ( .DIN1(n8423), .DIN2(n8424), .Q(n6482) );
  nnd2s1 U9102 ( .DIN1(n5826), .DIN2(n5569), .Q(n8424) );
  nnd3s1 U9103 ( .DIN1(n8425), .DIN2(n8426), .DIN3(n8312), .Q(n8402) );
  nnd4s1 U9104 ( .DIN1(n8427), .DIN2(n8428), .DIN3(n9486), .DIN4(n8429), 
        .Q(n8426) );
  and3s1 U9105 ( .DIN1(n8430), .DIN2(n8431), .DIN3(n8432), .Q(n8429) );
  nnd2s1 U9106 ( .DIN1(n5315), .DIN2(n7456), .Q(n8432) );
  nnd2s1 U9107 ( .DIN1(n5306), .DIN2(n8433), .Q(n8431) );
  nnd2s1 U9108 ( .DIN1(n8434), .DIN2(n8143), .Q(n8433) );
  nnd2s1 U9109 ( .DIN1(n789), .DIN2(n34), .Q(n8143) );
  nnd2s1 U9110 ( .DIN1(n6467), .DIN2(n806), .Q(n8430) );
  nnd2s1 U9111 ( .DIN1(n8423), .DIN2(n8435), .Q(n6467) );
  nnd2s1 U9112 ( .DIN1(n8436), .DIN2(n8437), .Q(n8435) );
  nnd2s1 U9113 ( .DIN1(n8438), .DIN2(n29), .Q(n8437) );
  and2s1 U9114 ( .DIN1(n8439), .DIN2(n8440), .Q(n8423) );
  nnd2s1 U9115 ( .DIN1(n544), .DIN2(n7452), .Q(n8440) );
  nnd2s1 U9116 ( .DIN1(n555), .DIN2(n7454), .Q(n8439) );
  nnd2s1 U9117 ( .DIN1(n719), .DIN2(n7455), .Q(n8428) );
  nnd2s1 U9118 ( .DIN1(n398), .DIN2(n7931), .Q(n8427) );
  nnd2s1 U9119 ( .DIN1(n8170), .DIN2(n759), .Q(n8425) );
  nnd2s1 U9120 ( .DIN1(n7206), .DIN2(n4831), .Q(n8400) );
  nnd2s1 U9121 ( .DIN1(n428), .DIN2(n8441), .Q(n8399) );
  nnd4s1 U9122 ( .DIN1(n8442), .DIN2(n8443), .DIN3(n8444), .DIN4(n7059), 
        .Q(n8441) );
  nnd2s1 U9123 ( .DIN1(n8445), .DIN2(n7212), .Q(n8444) );
  xnr2s1 U9124 ( .DIN1(n8282), .DIN2(n8283), .Q(n8445) );
  hi1s1 U9125 ( .DIN(n8446), .Q(n8283) );
  nnd2s1 U9126 ( .DIN1(n8447), .DIN2(n743), .Q(n8443) );
  xnr2s1 U9127 ( .DIN1(n8288), .DIN2(n8289), .Q(n8447) );
  hi1s1 U9128 ( .DIN(n8448), .Q(n8289) );
  nor2s1 U9129 ( .DIN1(n8449), .DIN2(n8450), .Q(n8442) );
  nor2s1 U9130 ( .DIN1(n4831), .DIN2(n7006), .Q(n8450) );
  nor2s1 U9131 ( .DIN1(n9486), .DIN2(n7037), .Q(n8449) );
  nnd2s1 U9132 ( .DIN1(n8451), .DIN2(n81), .Q(n8398) );
  nnd3s1 U9133 ( .DIN1(n8452), .DIN2(n8453), .DIN3(n8454), .Q(n8451) );
  nnd2s1 U9134 ( .DIN1(n7222), .DIN2(n4831), .Q(n8454) );
  nnd2s1 U9135 ( .DIN1(n8455), .DIN2(n722), .Q(n8453) );
  xnr2s1 U9136 ( .DIN1(n8282), .DIN2(n8446), .Q(n8455) );
  xnr2s1 U9137 ( .DIN1(n9486), .DIN2(n786), .Q(n8446) );
  nnd2s1 U9138 ( .DIN1(n8456), .DIN2(n8457), .Q(n8282) );
  nnd2s1 U9139 ( .DIN1(n433), .DIN2(n8458), .Q(n8457) );
  nnd2s1 U9140 ( .DIN1(n8459), .DIN2(n8460), .Q(n8458) );
  or2s1 U9141 ( .DIN1(n8460), .DIN2(n8459), .Q(n8456) );
  nnd2s1 U9142 ( .DIN1(n8461), .DIN2(n7058), .Q(n8452) );
  xnr2s1 U9143 ( .DIN1(n8448), .DIN2(n8288), .Q(n8461) );
  xnr2s1 U9144 ( .DIN1(n5423), .DIN2(n4831), .Q(n8448) );
  nnd2s1 U9145 ( .DIN1(n8462), .DIN2(n8463), .Q(n8288) );
  nnd2s1 U9146 ( .DIN1(n10), .DIN2(n8464), .Q(n8463) );
  nnd2s1 U9147 ( .DIN1(n8465), .DIN2(n393), .Q(n8464) );
  or2s1 U9148 ( .DIN1(n393), .DIN2(n8465), .Q(n8462) );
  nnd3s1 U9149 ( .DIN1(n8467), .DIN2(n8468), .DIN3(n8469), .Q(\EXinst/n1436 )
         );
  nnd2s1 U9150 ( .DIN1(n5394), .DIN2(\DM_addr[4] ), .Q(n8469) );
  nnd2s1 U9151 ( .DIN1(n5324), .DIN2(n8470), .Q(n8468) );
  nnd4s1 U9152 ( .DIN1(n8471), .DIN2(n8472), .DIN3(n8473), .DIN4(n8474), 
        .Q(n8470) );
  and4s1 U9153 ( .DIN1(n8475), .DIN2(n8476), .DIN3(n8477), .DIN4(n8478), 
        .Q(n8474) );
  nnd2s1 U9154 ( .DIN1(n8479), .DIN2(n8480), .Q(n8478) );
  nnd3s1 U9155 ( .DIN1(n8481), .DIN2(n5372), .DIN3(n8482), .Q(n8479) );
  nnd2s1 U9156 ( .DIN1(n620), .DIN2(n8360), .Q(n8482) );
  nnd2s1 U9157 ( .DIN1(n656), .DIN2(n8355), .Q(n8481) );
  hi1s1 U9158 ( .DIN(n8356), .Q(n8355) );
  nnd2s1 U9159 ( .DIN1(n8483), .DIN2(n8484), .Q(n8477) );
  nnd2s1 U9160 ( .DIN1(n8485), .DIN2(n8486), .Q(n8484) );
  nnd2s1 U9161 ( .DIN1(n655), .DIN2(n8356), .Q(n8486) );
  nnd2s1 U9162 ( .DIN1(n8487), .DIN2(n8488), .Q(n8356) );
  nnd2s1 U9163 ( .DIN1(n61), .DIN2(n8489), .Q(n8488) );
  nnd2s1 U9164 ( .DIN1(n8490), .DIN2(n77), .Q(n8489) );
  nnd2s1 U9165 ( .DIN1(n431), .DIN2(n8491), .Q(n8487) );
  or2s1 U9166 ( .DIN1(n8360), .DIN2(n5375), .Q(n8485) );
  nnd2s1 U9167 ( .DIN1(n8492), .DIN2(n8493), .Q(n8360) );
  nnd2s1 U9168 ( .DIN1(n8494), .DIN2(n8495), .Q(n8493) );
  nnd2s1 U9169 ( .DIN1(n752), .DIN2(n8496), .Q(n8476) );
  nnd2s1 U9170 ( .DIN1(n5471), .DIN2(n8497), .Q(n8496) );
  nnd2s1 U9171 ( .DIN1(n775), .DIN2(n10), .Q(n8497) );
  nnd2s1 U9172 ( .DIN1(n433), .DIN2(n768), .Q(n8475) );
  nnd2s1 U9173 ( .DIN1(n8498), .DIN2(n8499), .Q(n8473) );
  nnd3s1 U9174 ( .DIN1(n8500), .DIN2(n807), .DIN3(n8501), .Q(n8499) );
  hi1s1 U9175 ( .DIN(n8502), .Q(n8501) );
  nnd2s1 U9176 ( .DIN1(n628), .DIN2(n8503), .Q(n8500) );
  nnd2s1 U9177 ( .DIN1(n5994), .DIN2(n8504), .Q(n8498) );
  nnd2s1 U9178 ( .DIN1(n386), .DIN2(n6637), .Q(n8504) );
  nnd2s1 U9179 ( .DIN1(n8505), .DIN2(n8506), .Q(n6637) );
  nnd2s1 U9180 ( .DIN1(n547), .DIN2(n7539), .Q(n8506) );
  nnd3s1 U9181 ( .DIN1(n6658), .DIN2(n337), .DIN3(n7138), .Q(n8472) );
  nnd2s1 U9182 ( .DIN1(n8507), .DIN2(n8508), .Q(n6658) );
  nnd2s1 U9183 ( .DIN1(n7106), .DIN2(n741), .Q(n8508) );
  nnd2s1 U9184 ( .DIN1(n7100), .DIN2(n205), .Q(n8507) );
  nnd4s1 U9185 ( .DIN1(n8509), .DIN2(n8510), .DIN3(n8511), .DIN4(n8512), 
        .Q(n7100) );
  nnd2s1 U9186 ( .DIN1(n771), .DIN2(n426), .Q(n8512) );
  nnd2s1 U9187 ( .DIN1(n531), .DIN2(n432), .Q(n8511) );
  nnd3s1 U9188 ( .DIN1(n8513), .DIN2(n8514), .DIN3(n769), .Q(n8471) );
  nnd4s1 U9189 ( .DIN1(n8515), .DIN2(n5337), .DIN3(n8516), .DIN4(n8517), 
        .Q(n8514) );
  nnd2s1 U9190 ( .DIN1(n753), .DIN2(n6643), .Q(n8517) );
  nnd2s1 U9191 ( .DIN1(n8505), .DIN2(n8518), .Q(n6643) );
  nnd2s1 U9192 ( .DIN1(n8389), .DIN2(n8519), .Q(n8518) );
  nnd2s1 U9193 ( .DIN1(n8014), .DIN2(n205), .Q(n8519) );
  hi1s1 U9194 ( .DIN(n7539), .Q(n8014) );
  and2s1 U9195 ( .DIN1(n8520), .DIN2(n8521), .Q(n8505) );
  nnd2s1 U9196 ( .DIN1(n623), .DIN2(n7536), .Q(n8521) );
  nnd2s1 U9197 ( .DIN1(n628), .DIN2(n7537), .Q(n8520) );
  nnd2s1 U9198 ( .DIN1(n8502), .DIN2(n808), .Q(n8516) );
  nnd3s1 U9199 ( .DIN1(n8522), .DIN2(n8523), .DIN3(n8524), .Q(n8502) );
  nnd2s1 U9200 ( .DIN1(n622), .DIN2(n8003), .Q(n8524) );
  nnd2s1 U9201 ( .DIN1(n5876), .DIN2(n7535), .Q(n8523) );
  nnd2s1 U9202 ( .DIN1(n546), .DIN2(n7526), .Q(n8522) );
  nnd2s1 U9203 ( .DIN1(n5345), .DIN2(n8503), .Q(n8515) );
  and2s1 U9204 ( .DIN1(n629), .DIN2(n204), .Q(n5345) );
  nnd2s1 U9205 ( .DIN1(n8112), .DIN2(n6863), .Q(n8513) );
  nnd2s1 U9206 ( .DIN1(n551), .DIN2(n8525), .Q(n8467) );
  nnd4s1 U9207 ( .DIN1(n8526), .DIN2(n8527), .DIN3(n8528), .DIN4(n8529), 
        .Q(n8525) );
  and4s1 U9208 ( .DIN1(n8530), .DIN2(n8531), .DIN3(n8532), .DIN4(n8533), 
        .Q(n8529) );
  nnd2s1 U9209 ( .DIN1(n10), .DIN2(n8534), .Q(n8533) );
  nnd4s1 U9210 ( .DIN1(n8535), .DIN2(n8536), .DIN3(n8537), .DIN4(n7059), 
        .Q(n8534) );
  nnd2s1 U9211 ( .DIN1(n8538), .DIN2(n7212), .Q(n8537) );
  xnr2s1 U9212 ( .DIN1(n8460), .DIN2(n8459), .Q(n8538) );
  hi1s1 U9213 ( .DIN(n8539), .Q(n8459) );
  nnd2s1 U9214 ( .DIN1(n8540), .DIN2(n743), .Q(n8536) );
  xnr2s1 U9215 ( .DIN1(n393), .DIN2(n8465), .Q(n8540) );
  hi1s1 U9216 ( .DIN(n8541), .Q(n8465) );
  nnd2s1 U9217 ( .DIN1(n7314), .DIN2(n805), .Q(n8535) );
  nnd2s1 U9218 ( .DIN1(n8542), .DIN2(n334), .Q(n8532) );
  nnd2s1 U9219 ( .DIN1(n8543), .DIN2(n8544), .Q(n8542) );
  nnd2s1 U9220 ( .DIN1(n8545), .DIN2(n722), .Q(n8544) );
  xnr2s1 U9221 ( .DIN1(n8539), .DIN2(n8460), .Q(n8545) );
  xor2s1 U9222 ( .DIN1(n744), .DIN2(n56), .Q(n8460) );
  nnd2s1 U9223 ( .DIN1(n8546), .DIN2(n8547), .Q(n8539) );
  nnd2s1 U9224 ( .DIN1(n431), .DIN2(n8548), .Q(n8547) );
  or2s1 U9225 ( .DIN1(n8549), .DIN2(n8550), .Q(n8548) );
  nnd2s1 U9226 ( .DIN1(n8550), .DIN2(n8549), .Q(n8546) );
  nnd2s1 U9227 ( .DIN1(n8551), .DIN2(n7058), .Q(n8543) );
  xnr2s1 U9228 ( .DIN1(n8541), .DIN2(n393), .Q(n8551) );
  nnd2s1 U9229 ( .DIN1(n8552), .DIN2(n8553), .Q(n8541) );
  nnd2s1 U9230 ( .DIN1(n431), .DIN2(n8554), .Q(n8553) );
  or2s1 U9231 ( .DIN1(n8555), .DIN2(n8556), .Q(n8554) );
  nnd2s1 U9232 ( .DIN1(n8556), .DIN2(n8555), .Q(n8552) );
  or2s1 U9233 ( .DIN1(n8557), .DIN2(n7006), .Q(n8531) );
  nnd2s1 U9234 ( .DIN1(n7206), .DIN2(n806), .Q(n8530) );
  nnd2s1 U9235 ( .DIN1(n8312), .DIN2(n8558), .Q(n8528) );
  nnd4s1 U9236 ( .DIN1(n8559), .DIN2(n8560), .DIN3(n9486), .DIN4(n8561), 
        .Q(n8558) );
  and3s1 U9237 ( .DIN1(n8562), .DIN2(n8563), .DIN3(n8564), .Q(n8561) );
  nnd2s1 U9238 ( .DIN1(n5304), .DIN2(n7603), .Q(n8564) );
  nnd2s1 U9239 ( .DIN1(n6595), .DIN2(n805), .Q(n8563) );
  nnd2s1 U9240 ( .DIN1(n8565), .DIN2(n8566), .Q(n6595) );
  or2s1 U9241 ( .DIN1(n5740), .DIN2(n736), .Q(n8566) );
  nnd2s1 U9242 ( .DIN1(n8567), .DIN2(n8568), .Q(n5740) );
  nnd2s1 U9243 ( .DIN1(n7591), .DIN2(n747), .Q(n8567) );
  hi1s1 U9244 ( .DIN(n5742), .Q(n7591) );
  nnd2s1 U9245 ( .DIN1(n5315), .DIN2(n7604), .Q(n8562) );
  nnd2s1 U9246 ( .DIN1(n397), .DIN2(n8072), .Q(n8560) );
  nnd2s1 U9247 ( .DIN1(n5306), .DIN2(n8569), .Q(n8559) );
  and2s1 U9248 ( .DIN1(n7193), .DIN2(n8570), .Q(n8312) );
  nnd2s1 U9249 ( .DIN1(n8170), .DIN2(n792), .Q(n8570) );
  nnd4s1 U9250 ( .DIN1(n8571), .DIN2(n8572), .DIN3(n8573), .DIN4(n8574), 
        .Q(n8527) );
  and3s1 U9251 ( .DIN1(n8575), .DIN2(n8576), .DIN3(n730), .Q(n8574) );
  nnd2s1 U9252 ( .DIN1(n8577), .DIN2(n5306), .Q(n8576) );
  nor2s1 U9253 ( .DIN1(n6253), .DIN2(n206), .Q(n5306) );
  nnd2s1 U9254 ( .DIN1(n6659), .DIN2(n806), .Q(n8575) );
  and2s1 U9255 ( .DIN1(n8565), .DIN2(n8578), .Q(n6659) );
  nnd2s1 U9256 ( .DIN1(n5826), .DIN2(n5742), .Q(n8578) );
  and2s1 U9257 ( .DIN1(n8579), .DIN2(n8580), .Q(n8565) );
  nnd2s1 U9258 ( .DIN1(n545), .DIN2(n7601), .Q(n8580) );
  nnd2s1 U9259 ( .DIN1(n554), .DIN2(n7602), .Q(n8579) );
  nnd2s1 U9260 ( .DIN1(n8061), .DIN2(n398), .Q(n8573) );
  nnd2s1 U9261 ( .DIN1(n544), .DIN2(n739), .Q(n5303) );
  nnd2s1 U9262 ( .DIN1(n7586), .DIN2(n5315), .Q(n8572) );
  nnd2s1 U9263 ( .DIN1(n7590), .DIN2(n719), .Q(n8571) );
  hi1s1 U9264 ( .DIN(n7603), .Q(n7590) );
  nnd3s1 U9265 ( .DIN1(n9487), .DIN2(n6610), .DIN3(n400), .Q(n8526) );
  nnd2s1 U9266 ( .DIN1(n8581), .DIN2(n8582), .Q(n6610) );
  nnd2s1 U9267 ( .DIN1(n7026), .DIN2(n792), .Q(n8582) );
  nnd2s1 U9268 ( .DIN1(n747), .DIN2(n7024), .Q(n8581) );
  nnd4s1 U9269 ( .DIN1(n8583), .DIN2(n8584), .DIN3(n8585), .DIN4(n8586), 
        .Q(n7024) );
  nnd2s1 U9270 ( .DIN1(n784), .DIN2(n426), .Q(n8586) );
  nnd2s1 U9271 ( .DIN1(n758), .DIN2(n35), .Q(n8585) );
  nnd2s1 U9272 ( .DIN1(n790), .DIN2(n431), .Q(n8584) );
  nnd3s1 U9273 ( .DIN1(n8587), .DIN2(n8588), .DIN3(n8589), .Q(\EXinst/n1435 )
         );
  nnd2s1 U9274 ( .DIN1(n727), .DIN2(\DM_addr[3] ), .Q(n8589) );
  nnd2s1 U9275 ( .DIN1(n5324), .DIN2(n8590), .Q(n8588) );
  nnd4s1 U9276 ( .DIN1(n8591), .DIN2(n8592), .DIN3(n8593), .DIN4(n8594), 
        .Q(n8590) );
  and4s1 U9277 ( .DIN1(n8595), .DIN2(n8596), .DIN3(n8597), .DIN4(n8598), 
        .Q(n8594) );
  nnd2s1 U9278 ( .DIN1(n8599), .DIN2(n8600), .Q(n8598) );
  nnd3s1 U9279 ( .DIN1(n8601), .DIN2(n749), .DIN3(n8602), .Q(n8599) );
  nnd2s1 U9280 ( .DIN1(n705), .DIN2(n8494), .Q(n8602) );
  nnd2s1 U9281 ( .DIN1(n654), .DIN2(n8490), .Q(n8601) );
  hi1s1 U9282 ( .DIN(n8491), .Q(n8490) );
  nnd2s1 U9283 ( .DIN1(n8603), .DIN2(n8604), .Q(n8597) );
  nnd2s1 U9284 ( .DIN1(n8605), .DIN2(n8606), .Q(n8604) );
  nnd2s1 U9285 ( .DIN1(n653), .DIN2(n8491), .Q(n8606) );
  nnd2s1 U9286 ( .DIN1(n8607), .DIN2(n8608), .Q(n8491) );
  nnd2s1 U9287 ( .DIN1(n742), .DIN2(n8609), .Q(n8608) );
  nnd2s1 U9288 ( .DIN1(n8610), .DIN2(n80), .Q(n8609) );
  nnd2s1 U9289 ( .DIN1(n426), .DIN2(n8611), .Q(n8607) );
  or2s1 U9290 ( .DIN1(n8494), .DIN2(n5375), .Q(n8605) );
  nnd2s1 U9291 ( .DIN1(n8612), .DIN2(n8613), .Q(n8494) );
  nnd2s1 U9292 ( .DIN1(n8614), .DIN2(n8615), .Q(n8613) );
  hi1s1 U9293 ( .DIN(n8600), .Q(n8603) );
  nnd2s1 U9294 ( .DIN1(n8616), .DIN2(n6745), .Q(n8596) );
  nnd4s1 U9295 ( .DIN1(n8617), .DIN2(n8618), .DIN3(n8619), .DIN4(n8620), 
        .Q(n6745) );
  nnd2s1 U9296 ( .DIN1(n772), .DIN2(n432), .Q(n8620) );
  nnd2s1 U9297 ( .DIN1(n431), .DIN2(n767), .Q(n8595) );
  nnd2s1 U9298 ( .DIN1(n438), .DIN2(n8621), .Q(n8593) );
  nnd2s1 U9299 ( .DIN1(n5471), .DIN2(n8622), .Q(n8621) );
  nnd2s1 U9300 ( .DIN1(n776), .DIN2(n431), .Q(n8622) );
  nnd3s1 U9301 ( .DIN1(n8623), .DIN2(n8624), .DIN3(n5336), .Q(n8592) );
  nnd2s1 U9302 ( .DIN1(n8112), .DIN2(n6730), .Q(n8624) );
  hi1s1 U9303 ( .DIN(n5867), .Q(n6730) );
  nnd2s1 U9304 ( .DIN1(n6863), .DIN2(n8625), .Q(n5867) );
  nnd2s1 U9305 ( .DIN1(n754), .DIN2(reg_out_A[31]), .Q(n8625) );
  nnd3s1 U9306 ( .DIN1(n8626), .DIN2(n8627), .DIN3(n5337), .Q(n8623) );
  nnd2s1 U9307 ( .DIN1(n752), .DIN2(n8628), .Q(n8627) );
  nnd2s1 U9308 ( .DIN1(n8629), .DIN2(n6724), .Q(n8628) );
  nnd2s1 U9309 ( .DIN1(n8389), .DIN2(n8630), .Q(n6724) );
  nnd2s1 U9310 ( .DIN1(n6299), .DIN2(n5490), .Q(n8630) );
  hi1s1 U9311 ( .DIN(n5863), .Q(n6299) );
  and2s1 U9312 ( .DIN1(n438), .DIN2(n8631), .Q(n8389) );
  nnd2s1 U9313 ( .DIN1(n32), .DIN2(n62), .Q(n8631) );
  nnd3s1 U9314 ( .DIN1(n8632), .DIN2(n8633), .DIN3(n808), .Q(n8626) );
  nnd2s1 U9315 ( .DIN1(n8634), .DIN2(n8635), .Q(n8591) );
  nnd2s1 U9316 ( .DIN1(n808), .DIN2(n8636), .Q(n8635) );
  nnd2s1 U9317 ( .DIN1(n8632), .DIN2(n8633), .Q(n8636) );
  nnd3s1 U9318 ( .DIN1(n8637), .DIN2(n8638), .DIN3(n801), .Q(n8633) );
  nnd2s1 U9319 ( .DIN1(n741), .DIN2(n8118), .Q(n8638) );
  nnd3s1 U9320 ( .DIN1(n7870), .DIN2(n8639), .DIN3(n8104), .Q(n8118) );
  nnd2s1 U9321 ( .DIN1(n755), .DIN2(n429), .Q(n8104) );
  nnd3s1 U9322 ( .DIN1(n8640), .DIN2(n8641), .DIN3(reg_out_B[1]), .Q(n8639) );
  nnd2s1 U9323 ( .DIN1(n66), .DIN2(n1), .Q(n8641) );
  nnd2s1 U9324 ( .DIN1(n399), .DIN2(n65), .Q(n8640) );
  nnd2s1 U9325 ( .DIN1(n773), .DIN2(n425), .Q(n7870) );
  nnd2s1 U9326 ( .DIN1(n8642), .DIN2(n5490), .Q(n8637) );
  nnd4s1 U9327 ( .DIN1(n8617), .DIN2(n8375), .DIN3(n7871), .DIN4(n8107), 
        .Q(n8642) );
  nnd2s1 U9328 ( .DIN1(n771), .DIN2(n428), .Q(n8107) );
  nnd2s1 U9329 ( .DIN1(n532), .DIN2(n427), .Q(n7871) );
  nnd2s1 U9330 ( .DIN1(n774), .DIN2(n433), .Q(n8375) );
  nnd2s1 U9331 ( .DIN1(n754), .DIN2(n431), .Q(n8617) );
  nnd3s1 U9332 ( .DIN1(n8643), .DIN2(n8644), .DIN3(n438), .Q(n8632) );
  nnd2s1 U9333 ( .DIN1(n742), .DIN2(n7163), .Q(n8644) );
  nnd4s1 U9334 ( .DIN1(n7144), .DIN2(n6959), .DIN3(n6527), .DIN4(n6742), 
        .Q(n7163) );
  nnd2s1 U9335 ( .DIN1(n772), .DIN2(n416), .Q(n6742) );
  nnd2s1 U9336 ( .DIN1(n531), .DIN2(n415), .Q(n6527) );
  nnd2s1 U9337 ( .DIN1(n773), .DIN2(n417), .Q(n6959) );
  nnd2s1 U9338 ( .DIN1(n755), .DIN2(n418), .Q(n7144) );
  nnd2s1 U9339 ( .DIN1(n7651), .DIN2(n5490), .Q(n8643) );
  nnd4s1 U9340 ( .DIN1(n7639), .DIN2(n7391), .DIN3(n6960), .DIN4(n7147), 
        .Q(n7651) );
  nnd2s1 U9341 ( .DIN1(n771), .DIN2(n420), .Q(n7147) );
  nnd2s1 U9342 ( .DIN1(n532), .DIN2(n419), .Q(n6960) );
  nnd2s1 U9343 ( .DIN1(n774), .DIN2(n421), .Q(n7391) );
  nnd2s1 U9344 ( .DIN1(n754), .DIN2(n422), .Q(n7639) );
  nnd2s1 U9345 ( .DIN1(n5994), .DIN2(n8645), .Q(n8634) );
  nnd2s1 U9346 ( .DIN1(n386), .DIN2(n6717), .Q(n8645) );
  nnd2s1 U9347 ( .DIN1(n8629), .DIN2(n8646), .Q(n6717) );
  nnd2s1 U9348 ( .DIN1(n61), .DIN2(n5857), .Q(n8646) );
  nnd2s1 U9349 ( .DIN1(n8647), .DIN2(n8648), .Q(n5857) );
  nnd2s1 U9350 ( .DIN1(n8243), .DIN2(n755), .Q(n8648) );
  nnd2s1 U9351 ( .DIN1(n5863), .DIN2(n5490), .Q(n8647) );
  nnd4s1 U9352 ( .DIN1(n5877), .DIN2(n5637), .DIN3(n8649), .DIN4(n8650), 
        .Q(n5863) );
  nnd2s1 U9353 ( .DIN1(n772), .DIN2(n406), .Q(n8650) );
  nnd2s1 U9354 ( .DIN1(reg_out_A[30]), .DIN2(n532), .Q(n8649) );
  nnd2s1 U9355 ( .DIN1(n773), .DIN2(n12), .Q(n5637) );
  nnd2s1 U9356 ( .DIN1(n755), .DIN2(n407), .Q(n5877) );
  and2s1 U9357 ( .DIN1(n8651), .DIN2(n8652), .Q(n8629) );
  nnd2s1 U9358 ( .DIN1(n621), .DIN2(n6729), .Q(n8652) );
  nnd4s1 U9359 ( .DIN1(n6310), .DIN2(n6096), .DIN3(n5638), .DIN4(n5880), 
        .Q(n6729) );
  nnd2s1 U9360 ( .DIN1(n771), .DIN2(n408), .Q(n5880) );
  nnd2s1 U9361 ( .DIN1(n531), .DIN2(n435), .Q(n5638) );
  nnd2s1 U9362 ( .DIN1(n774), .DIN2(n409), .Q(n6096) );
  nnd2s1 U9363 ( .DIN1(n754), .DIN2(n410), .Q(n6310) );
  nnd2s1 U9364 ( .DIN1(n628), .DIN2(n6728), .Q(n8651) );
  nnd4s1 U9365 ( .DIN1(n6739), .DIN2(n6526), .DIN3(n8653), .DIN4(n6313), 
        .Q(n6728) );
  nnd2s1 U9366 ( .DIN1(n772), .DIN2(n412), .Q(n6313) );
  nnd2s1 U9367 ( .DIN1(n532), .DIN2(n411), .Q(n8653) );
  nnd2s1 U9368 ( .DIN1(n773), .DIN2(n413), .Q(n6526) );
  nnd2s1 U9369 ( .DIN1(n755), .DIN2(n414), .Q(n6739) );
  nnd2s1 U9370 ( .DIN1(n550), .DIN2(n8654), .Q(n8587) );
  nnd4s1 U9371 ( .DIN1(n8655), .DIN2(n8656), .DIN3(n8657), .DIN4(n8658), 
        .Q(n8654) );
  and3s1 U9372 ( .DIN1(n8659), .DIN2(n8660), .DIN3(n8661), .Q(n8658) );
  nnd2s1 U9373 ( .DIN1(n7206), .DIN2(n4840), .Q(n8661) );
  nnd2s1 U9374 ( .DIN1(n431), .DIN2(n8662), .Q(n8660) );
  nnd4s1 U9375 ( .DIN1(n8663), .DIN2(n8664), .DIN3(n8665), .DIN4(n7059), 
        .Q(n8662) );
  nnd2s1 U9376 ( .DIN1(n8666), .DIN2(n7212), .Q(n8665) );
  xnr2s1 U9377 ( .DIN1(n8549), .DIN2(n8550), .Q(n8666) );
  hi1s1 U9378 ( .DIN(n8667), .Q(n8550) );
  nnd2s1 U9379 ( .DIN1(n8668), .DIN2(n743), .Q(n8664) );
  xnr2s1 U9380 ( .DIN1(n8555), .DIN2(n8556), .Q(n8668) );
  hi1s1 U9381 ( .DIN(n8669), .Q(n8556) );
  nor2s1 U9382 ( .DIN1(n8670), .DIN2(n8671), .Q(n8663) );
  nor2s1 U9383 ( .DIN1(n4840), .DIN2(n7006), .Q(n8671) );
  nor2s1 U9384 ( .DIN1(n9487), .DIN2(n7037), .Q(n8670) );
  nnd2s1 U9385 ( .DIN1(n8672), .DIN2(n77), .Q(n8659) );
  nnd3s1 U9386 ( .DIN1(n8673), .DIN2(n8674), .DIN3(n8675), .Q(n8672) );
  nnd2s1 U9387 ( .DIN1(n7222), .DIN2(n4840), .Q(n8675) );
  nnd2s1 U9388 ( .DIN1(n8676), .DIN2(n722), .Q(n8674) );
  xnr2s1 U9389 ( .DIN1(n8549), .DIN2(n8667), .Q(n8676) );
  xnr2s1 U9390 ( .DIN1(n745), .DIN2(n802), .Q(n8667) );
  nnd2s1 U9391 ( .DIN1(n8677), .DIN2(n8678), .Q(n8549) );
  nnd2s1 U9392 ( .DIN1(n426), .DIN2(n8679), .Q(n8678) );
  nnd2s1 U9393 ( .DIN1(n8680), .DIN2(n8681), .Q(n8679) );
  or2s1 U9394 ( .DIN1(n8681), .DIN2(n8680), .Q(n8677) );
  nnd2s1 U9395 ( .DIN1(n8682), .DIN2(n7058), .Q(n8673) );
  xnr2s1 U9396 ( .DIN1(n8555), .DIN2(n8669), .Q(n8682) );
  xnr2s1 U9397 ( .DIN1(n633), .DIN2(n802), .Q(n8669) );
  nnd2s1 U9398 ( .DIN1(n8683), .DIN2(n8684), .Q(n8555) );
  nnd2s1 U9399 ( .DIN1(n426), .DIN2(n8685), .Q(n8684) );
  nnd2s1 U9400 ( .DIN1(n8686), .DIN2(n395), .Q(n8685) );
  or2s1 U9401 ( .DIN1(n395), .DIN2(n8686), .Q(n8683) );
  nnd3s1 U9402 ( .DIN1(n555), .DIN2(n6689), .DIN3(n400), .Q(n8657) );
  nnd4s1 U9403 ( .DIN1(n8688), .DIN2(n8689), .DIN3(n8690), .DIN4(n8691), 
        .Q(n6689) );
  nnd2s1 U9404 ( .DIN1(n783), .DIN2(n35), .Q(n8691) );
  nnd2s1 U9405 ( .DIN1(n759), .DIN2(n33), .Q(n8690) );
  nnd2s1 U9406 ( .DIN1(n789), .DIN2(n426), .Q(n8689) );
  nnd2s1 U9407 ( .DIN1(n553), .DIN2(n431), .Q(n8688) );
  nnd3s1 U9408 ( .DIN1(n7339), .DIN2(n8692), .DIN3(n8693), .Q(n8656) );
  hi1s1 U9409 ( .DIN(n8694), .Q(n8693) );
  or2s1 U9410 ( .DIN1(n6690), .DIN2(n740), .Q(n8692) );
  nnd2s1 U9411 ( .DIN1(n6672), .DIN2(n8695), .Q(n6690) );
  nnd2s1 U9412 ( .DIN1(n5830), .DIN2(n803), .Q(n8695) );
  nnd2s1 U9413 ( .DIN1(n8696), .DIN2(n8697), .Q(n5830) );
  nnd2s1 U9414 ( .DIN1(n8325), .DIN2(n552), .Q(n8697) );
  nnd2s1 U9415 ( .DIN1(n29), .DIN2(n5807), .Q(n8696) );
  and2s1 U9416 ( .DIN1(n8698), .DIN2(n8699), .Q(n6672) );
  nnd2s1 U9417 ( .DIN1(n545), .DIN2(n7203), .Q(n8699) );
  nnd2s1 U9418 ( .DIN1(n555), .DIN2(n7693), .Q(n8698) );
  nnd4s1 U9419 ( .DIN1(n7193), .DIN2(n8700), .DIN3(n8701), .DIN4(n8702), 
        .Q(n8655) );
  nnd3s1 U9420 ( .DIN1(n8703), .DIN2(n6673), .DIN3(n7836), .Q(n8702) );
  nnd2s1 U9421 ( .DIN1(n8436), .DIN2(n8704), .Q(n6673) );
  nnd2s1 U9422 ( .DIN1(n7191), .DIN2(n29), .Q(n8704) );
  hi1s1 U9423 ( .DIN(n5807), .Q(n7191) );
  nnd4s1 U9424 ( .DIN1(n5819), .DIN2(n5594), .DIN3(n8705), .DIN4(n8706), 
        .Q(n5807) );
  nnd2s1 U9425 ( .DIN1(n784), .DIN2(n406), .Q(n8706) );
  nnd2s1 U9426 ( .DIN1(n718), .DIN2(n758), .Q(n8705) );
  nnd2s1 U9427 ( .DIN1(n790), .DIN2(n434), .Q(n5594) );
  nnd2s1 U9428 ( .DIN1(n552), .DIN2(n407), .Q(n5819) );
  and2s1 U9429 ( .DIN1(n735), .DIN2(n8568), .Q(n8436) );
  nnd2s1 U9430 ( .DIN1(n4845), .DIN2(n401), .Q(n8568) );
  nnd3s1 U9431 ( .DIN1(n8707), .DIN2(n8708), .DIN3(n736), .Q(n8703) );
  nnd2s1 U9432 ( .DIN1(n7192), .DIN2(n4845), .Q(n8708) );
  hi1s1 U9433 ( .DIN(n7203), .Q(n7192) );
  nnd4s1 U9434 ( .DIN1(n6254), .DIN2(n6045), .DIN3(n5595), .DIN4(n5822), 
        .Q(n7203) );
  nnd2s1 U9435 ( .DIN1(n783), .DIN2(n408), .Q(n5822) );
  nnd2s1 U9436 ( .DIN1(n758), .DIN2(n6), .Q(n5595) );
  nnd2s1 U9437 ( .DIN1(n789), .DIN2(n409), .Q(n6045) );
  nnd2s1 U9438 ( .DIN1(n553), .DIN2(n410), .Q(n6254) );
  nnd2s1 U9439 ( .DIN1(n7189), .DIN2(n747), .Q(n8707) );
  hi1s1 U9440 ( .DIN(n7693), .Q(n7189) );
  nnd4s1 U9441 ( .DIN1(n6682), .DIN2(n6476), .DIN3(n8709), .DIN4(n6257), 
        .Q(n7693) );
  nnd2s1 U9442 ( .DIN1(n784), .DIN2(n412), .Q(n6257) );
  nnd2s1 U9443 ( .DIN1(n758), .DIN2(n411), .Q(n8709) );
  nnd2s1 U9444 ( .DIN1(n790), .DIN2(n413), .Q(n6476) );
  nnd2s1 U9445 ( .DIN1(n552), .DIN2(n414), .Q(n6682) );
  or2s1 U9446 ( .DIN1(n5811), .DIN2(n8063), .Q(n8701) );
  hi1s1 U9447 ( .DIN(n8170), .Q(n8063) );
  nnd2s1 U9448 ( .DIN1(n5741), .DIN2(n8710), .Q(n5811) );
  nnd2s1 U9449 ( .DIN1(n553), .DIN2(n734), .Q(n8710) );
  nnd2s1 U9450 ( .DIN1(n9486), .DIN2(n8694), .Q(n8700) );
  nnd3s1 U9451 ( .DIN1(n8711), .DIN2(n8712), .DIN3(n8713), .Q(n8694) );
  nnd4s1 U9452 ( .DIN1(n8714), .DIN2(n56), .DIN3(n9487), .DIN4(n8715), 
        .Q(n8713) );
  nnd2s1 U9453 ( .DIN1(n9489), .DIN2(n8716), .Q(n8715) );
  nor2s1 U9454 ( .DIN1(n8717), .DIN2(n8718), .Q(n8714) );
  nor2s1 U9455 ( .DIN1(n8719), .DIN2(n4845), .Q(n8718) );
  nor2s1 U9456 ( .DIN1(n8720), .DIN2(n8721), .Q(n8719) );
  and2s1 U9457 ( .DIN1(n433), .DIN2(n790), .Q(n8721) );
  nor2s1 U9458 ( .DIN1(n333), .DIN2(n5313), .Q(n8720) );
  nor2s1 U9459 ( .DIN1(n747), .DIN2(n8166), .Q(n8717) );
  and2s1 U9460 ( .DIN1(n8153), .DIN2(n7908), .Q(n8166) );
  nnd2s1 U9461 ( .DIN1(n789), .DIN2(n36), .Q(n7908) );
  nnd3s1 U9462 ( .DIN1(n8722), .DIN2(n8723), .DIN3(n707), .Q(n8153) );
  nnd2s1 U9463 ( .DIN1(n9489), .DIN2(n66), .Q(n8723) );
  nnd2s1 U9464 ( .DIN1(n439), .DIN2(n65), .Q(n8722) );
  nnd2s1 U9465 ( .DIN1(n7684), .DIN2(n5315), .Q(n8712) );
  hi1s1 U9466 ( .DIN(n7697), .Q(n7684) );
  nnd4s1 U9467 ( .DIN1(n7674), .DIN2(n7428), .DIN3(n6909), .DIN4(n7181), 
        .Q(n7697) );
  nnd2s1 U9468 ( .DIN1(n783), .DIN2(n420), .Q(n7181) );
  nnd2s1 U9469 ( .DIN1(n759), .DIN2(n419), .Q(n6909) );
  nnd2s1 U9470 ( .DIN1(n790), .DIN2(n421), .Q(n7428) );
  nnd2s1 U9471 ( .DIN1(n552), .DIN2(n422), .Q(n7674) );
  nnd2s1 U9472 ( .DIN1(n7204), .DIN2(n5304), .Q(n8711) );
  hi1s1 U9473 ( .DIN(n7696), .Q(n7204) );
  nnd4s1 U9474 ( .DIN1(n7178), .DIN2(n6908), .DIN3(n6477), .DIN4(n6685), 
        .Q(n7696) );
  nnd2s1 U9475 ( .DIN1(n784), .DIN2(n416), .Q(n6685) );
  nnd2s1 U9476 ( .DIN1(n758), .DIN2(n415), .Q(n6477) );
  nnd2s1 U9477 ( .DIN1(n789), .DIN2(n417), .Q(n6908) );
  nnd2s1 U9478 ( .DIN1(n553), .DIN2(n418), .Q(n7178) );
  nnd3s1 U9479 ( .DIN1(n8724), .DIN2(n8725), .DIN3(n8726), .Q(\EXinst/n1434 )
         );
  nnd2s1 U9480 ( .DIN1(n5394), .DIN2(\DM_addr[2] ), .Q(n8726) );
  or2s1 U9481 ( .DIN1(n8727), .DIN2(n8728), .Q(n8725) );
  nor2s1 U9482 ( .DIN1(n8729), .DIN2(n8730), .Q(n8727) );
  nnd4s1 U9483 ( .DIN1(n8731), .DIN2(n8732), .DIN3(n8733), .DIN4(n8734), 
        .Q(n8730) );
  nnd2s1 U9484 ( .DIN1(n8735), .DIN2(n8736), .Q(n8734) );
  nnd3s1 U9485 ( .DIN1(n8737), .DIN2(n5372), .DIN3(n8738), .Q(n8735) );
  nnd2s1 U9486 ( .DIN1(n620), .DIN2(n8615), .Q(n8738) );
  nnd2s1 U9487 ( .DIN1(n656), .DIN2(n8610), .Q(n8737) );
  hi1s1 U9488 ( .DIN(n8611), .Q(n8610) );
  nnd3s1 U9489 ( .DIN1(n653), .DIN2(n8611), .DIN3(n8739), .Q(n8733) );
  nnd2s1 U9490 ( .DIN1(n8619), .DIN2(n8740), .Q(n8611) );
  nnd2s1 U9491 ( .DIN1(n432), .DIN2(n8741), .Q(n8740) );
  nnd2s1 U9492 ( .DIN1(n714), .DIN2(n8742), .Q(n8741) );
  nnd2s1 U9493 ( .DIN1(n531), .DIN2(n430), .Q(n8619) );
  nnd2s1 U9494 ( .DIN1(n8743), .DIN2(n705), .Q(n8732) );
  nnd2s1 U9495 ( .DIN1(n426), .DIN2(n768), .Q(n8731) );
  nnd4s1 U9496 ( .DIN1(n8744), .DIN2(n8745), .DIN3(n8746), .DIN4(n8747), 
        .Q(n8729) );
  nnd3s1 U9497 ( .DIN1(n8748), .DIN2(n8749), .DIN3(n769), .Q(n8747) );
  nnd3s1 U9498 ( .DIN1(n8750), .DIN2(n8751), .DIN3(n5337), .Q(n8749) );
  nnd2s1 U9499 ( .DIN1(n752), .DIN2(n6865), .Q(n8751) );
  nnd2s1 U9500 ( .DIN1(n8752), .DIN2(n8753), .Q(n6865) );
  nnd2s1 U9501 ( .DIN1(n438), .DIN2(n6000), .Q(n8753) );
  nnd2s1 U9502 ( .DIN1(n8754), .DIN2(n8755), .Q(n6000) );
  nnd2s1 U9503 ( .DIN1(n8243), .DIN2(n5353), .Q(n8755) );
  nnd3s1 U9504 ( .DIN1(n8756), .DIN2(n8757), .DIN3(n204), .Q(n8750) );
  nnd2s1 U9505 ( .DIN1(n8112), .DIN2(n8758), .Q(n8748) );
  nnd2s1 U9506 ( .DIN1(n734), .DIN2(n7765), .Q(n8758) );
  nnd2s1 U9507 ( .DIN1(reg_out_B[1]), .DIN2(n6863), .Q(n7765) );
  nor2s1 U9508 ( .DIN1(n7089), .DIN2(n7156), .Q(n8112) );
  nnd2s1 U9509 ( .DIN1(n8759), .DIN2(n8760), .Q(n8746) );
  nnd2s1 U9510 ( .DIN1(n204), .DIN2(n8761), .Q(n8760) );
  nnd2s1 U9511 ( .DIN1(n8756), .DIN2(n8757), .Q(n8761) );
  nnd3s1 U9512 ( .DIN1(n8762), .DIN2(n8763), .DIN3(n337), .Q(n8757) );
  nnd2s1 U9513 ( .DIN1(n32), .DIN2(n8245), .Q(n8763) );
  nnd3s1 U9514 ( .DIN1(n7992), .DIN2(n8764), .DIN3(n8227), .Q(n8245) );
  nnd2s1 U9515 ( .DIN1(n754), .DIN2(n34), .Q(n8227) );
  nnd3s1 U9516 ( .DIN1(n8765), .DIN2(n8766), .DIN3(reg_out_B[1]), .Q(n8764) );
  nnd2s1 U9517 ( .DIN1(n399), .DIN2(n66), .Q(n8766) );
  nnd2s1 U9518 ( .DIN1(n332), .DIN2(n1), .Q(n8765) );
  nnd2s1 U9519 ( .DIN1(n774), .DIN2(n429), .Q(n7992) );
  nnd2s1 U9520 ( .DIN1(n8767), .DIN2(n5490), .Q(n8762) );
  nnd4s1 U9521 ( .DIN1(n8768), .DIN2(n8510), .DIN3(n7993), .DIN4(n8230), 
        .Q(n8767) );
  nnd2s1 U9522 ( .DIN1(n771), .DIN2(n10), .Q(n8230) );
  nnd2s1 U9523 ( .DIN1(n532), .DIN2(n428), .Q(n7993) );
  nnd2s1 U9524 ( .DIN1(n773), .DIN2(n431), .Q(n8510) );
  nnd3s1 U9525 ( .DIN1(n8769), .DIN2(n8770), .DIN3(n61), .Q(n8756) );
  nnd2s1 U9526 ( .DIN1(n741), .DIN2(n7281), .Q(n8770) );
  nnd4s1 U9527 ( .DIN1(n7268), .DIN2(n7102), .DIN3(n6655), .DIN4(n6877), 
        .Q(n7281) );
  nnd2s1 U9528 ( .DIN1(n772), .DIN2(n417), .Q(n6877) );
  nnd2s1 U9529 ( .DIN1(n531), .DIN2(n416), .Q(n6655) );
  nnd2s1 U9530 ( .DIN1(n774), .DIN2(n418), .Q(n7102) );
  nnd2s1 U9531 ( .DIN1(n755), .DIN2(n419), .Q(n7268) );
  nnd2s1 U9532 ( .DIN1(n7770), .DIN2(n5490), .Q(n8769) );
  nnd4s1 U9533 ( .DIN1(n7756), .DIN2(n7515), .DIN3(n7103), .DIN4(n7271), 
        .Q(n7770) );
  nnd2s1 U9534 ( .DIN1(n771), .DIN2(n421), .Q(n7271) );
  nnd2s1 U9535 ( .DIN1(n532), .DIN2(n420), .Q(n7103) );
  nnd2s1 U9536 ( .DIN1(n773), .DIN2(n422), .Q(n7515) );
  nnd2s1 U9537 ( .DIN1(n754), .DIN2(n423), .Q(n7756) );
  nnd2s1 U9538 ( .DIN1(n5994), .DIN2(n8771), .Q(n8759) );
  nnd2s1 U9539 ( .DIN1(n386), .DIN2(n6857), .Q(n8771) );
  nnd2s1 U9540 ( .DIN1(n8752), .DIN2(n8772), .Q(n6857) );
  nnd2s1 U9541 ( .DIN1(n61), .DIN2(n5993), .Q(n8772) );
  nnd2s1 U9542 ( .DIN1(n8754), .DIN2(n8773), .Q(n5993) );
  nnd2s1 U9543 ( .DIN1(n8243), .DIN2(n773), .Q(n8773) );
  nor2s1 U9544 ( .DIN1(n5490), .DIN2(n62), .Q(n8243) );
  and2s1 U9545 ( .DIN1(n8774), .DIN2(n8775), .Q(n8754) );
  nnd2s1 U9546 ( .DIN1(n5495), .DIN2(n742), .Q(n8775) );
  nor2s1 U9547 ( .DIN1(n717), .DIN2(n5353), .Q(n5495) );
  nnd2s1 U9548 ( .DIN1(n7292), .DIN2(n5490), .Q(n8774) );
  nnd4s1 U9549 ( .DIN1(n6014), .DIN2(n5785), .DIN3(n8776), .DIN4(n5493), 
        .Q(n7292) );
  nnd2s1 U9550 ( .DIN1(n772), .DIN2(n12), .Q(n5493) );
  nnd2s1 U9551 ( .DIN1(n531), .DIN2(n406), .Q(n8776) );
  nnd2s1 U9552 ( .DIN1(n774), .DIN2(n407), .Q(n5785) );
  nnd2s1 U9553 ( .DIN1(n755), .DIN2(n435), .Q(n6014) );
  and2s1 U9554 ( .DIN1(n8777), .DIN2(n8778), .Q(n8752) );
  nnd2s1 U9555 ( .DIN1(n623), .DIN2(n7293), .Q(n8778) );
  nnd4s1 U9556 ( .DIN1(n6446), .DIN2(n6225), .DIN3(n5786), .DIN4(n8779), 
        .Q(n7293) );
  nnd2s1 U9557 ( .DIN1(n771), .DIN2(n409), .Q(n8779) );
  nnd2s1 U9558 ( .DIN1(n532), .DIN2(n408), .Q(n5786) );
  nnd2s1 U9559 ( .DIN1(n773), .DIN2(n410), .Q(n6225) );
  nnd2s1 U9560 ( .DIN1(n754), .DIN2(n411), .Q(n6446) );
  nnd2s1 U9561 ( .DIN1(n628), .DIN2(n7291), .Q(n8777) );
  nnd4s1 U9562 ( .DIN1(n6874), .DIN2(n6654), .DIN3(n8780), .DIN4(n6449), 
        .Q(n7291) );
  nnd2s1 U9563 ( .DIN1(n772), .DIN2(n413), .Q(n6449) );
  nnd2s1 U9564 ( .DIN1(n531), .DIN2(n412), .Q(n8780) );
  nnd2s1 U9565 ( .DIN1(n774), .DIN2(n414), .Q(n6654) );
  nnd2s1 U9566 ( .DIN1(n755), .DIN2(n415), .Q(n6874) );
  nnd2s1 U9567 ( .DIN1(n742), .DIN2(n8781), .Q(n8745) );
  nnd2s1 U9568 ( .DIN1(n5471), .DIN2(n8782), .Q(n8781) );
  nnd2s1 U9569 ( .DIN1(n775), .DIN2(n426), .Q(n8782) );
  nnd2s1 U9570 ( .DIN1(n8616), .DIN2(n6879), .Q(n8744) );
  nnd3s1 U9571 ( .DIN1(n8783), .DIN2(n8784), .DIN3(n8768), .Q(n6879) );
  nnd2s1 U9572 ( .DIN1(n754), .DIN2(n426), .Q(n8768) );
  nnd2s1 U9573 ( .DIN1(n771), .DIN2(n33), .Q(n8784) );
  nnd2s1 U9574 ( .DIN1(n773), .DIN2(n432), .Q(n8783) );
  nnd2s1 U9575 ( .DIN1(n9453), .DIN2(n8785), .Q(n8724) );
  nnd4s1 U9576 ( .DIN1(n8786), .DIN2(n8787), .DIN3(n8788), .DIN4(n8789), 
        .Q(n8785) );
  and4s1 U9577 ( .DIN1(n8790), .DIN2(n8791), .DIN3(n8792), .DIN4(n8793), 
        .Q(n8789) );
  nnd2s1 U9578 ( .DIN1(n426), .DIN2(n8794), .Q(n8793) );
  nnd4s1 U9579 ( .DIN1(n8795), .DIN2(n8796), .DIN3(n8797), .DIN4(n7059), 
        .Q(n8794) );
  nnd2s1 U9580 ( .DIN1(n8798), .DIN2(n7212), .Q(n8797) );
  xnr2s1 U9581 ( .DIN1(n8681), .DIN2(n8680), .Q(n8798) );
  hi1s1 U9582 ( .DIN(n8799), .Q(n8680) );
  nnd2s1 U9583 ( .DIN1(n8800), .DIN2(n743), .Q(n8796) );
  xnr2s1 U9584 ( .DIN1(n395), .DIN2(n8686), .Q(n8800) );
  hi1s1 U9585 ( .DIN(n8801), .Q(n8686) );
  nnd2s1 U9586 ( .DIN1(n7314), .DIN2(n4845), .Q(n8795) );
  nnd2s1 U9587 ( .DIN1(n8802), .DIN2(n80), .Q(n8792) );
  nnd2s1 U9588 ( .DIN1(n8803), .DIN2(n8804), .Q(n8802) );
  nnd2s1 U9589 ( .DIN1(n8805), .DIN2(n722), .Q(n8804) );
  xnr2s1 U9590 ( .DIN1(n8799), .DIN2(n8681), .Q(n8805) );
  xor2s1 U9591 ( .DIN1(n744), .DIN2(n746), .Q(n8681) );
  nnd2s1 U9592 ( .DIN1(n8806), .DIN2(n8807), .Q(n8799) );
  nnd2s1 U9593 ( .DIN1(n35), .DIN2(n8808), .Q(n8807) );
  or2s1 U9594 ( .DIN1(n8809), .DIN2(n8810), .Q(n8808) );
  nnd2s1 U9595 ( .DIN1(n8810), .DIN2(n8809), .Q(n8806) );
  nnd2s1 U9596 ( .DIN1(n8811), .DIN2(n7058), .Q(n8803) );
  xnr2s1 U9597 ( .DIN1(n8801), .DIN2(n395), .Q(n8811) );
  xor2s1 U9598 ( .DIN1(n632), .DIN2(n746), .Q(n8687) );
  nnd2s1 U9599 ( .DIN1(n8812), .DIN2(n8813), .Q(n8801) );
  nnd2s1 U9600 ( .DIN1(n432), .DIN2(n8814), .Q(n8813) );
  or2s1 U9601 ( .DIN1(n8815), .DIN2(n8816), .Q(n8814) );
  nnd2s1 U9602 ( .DIN1(n8816), .DIN2(n8815), .Q(n8812) );
  nnd2s1 U9603 ( .DIN1(n7222), .DIN2(n8817), .Q(n8791) );
  nnd2s1 U9604 ( .DIN1(n7206), .DIN2(n4845), .Q(n8790) );
  nnd3s1 U9605 ( .DIN1(n554), .DIN2(n6830), .DIN3(n400), .Q(n8788) );
  nnd3s1 U9606 ( .DIN1(n8818), .DIN2(n8819), .DIN3(n8820), .Q(n6830) );
  nnd2s1 U9607 ( .DIN1(n552), .DIN2(n426), .Q(n8820) );
  nnd2s1 U9608 ( .DIN1(n783), .DIN2(n430), .Q(n8819) );
  nnd2s1 U9609 ( .DIN1(n790), .DIN2(n35), .Q(n8818) );
  nnd3s1 U9610 ( .DIN1(n7339), .DIN2(n8821), .DIN3(n8822), .Q(n8787) );
  hi1s1 U9611 ( .DIN(n8823), .Q(n8822) );
  nnd2s1 U9612 ( .DIN1(n6880), .DIN2(n805), .Q(n8821) );
  and2s1 U9613 ( .DIN1(n6814), .DIN2(n8824), .Q(n6880) );
  nnd2s1 U9614 ( .DIN1(n5943), .DIN2(n735), .Q(n8824) );
  nnd2s1 U9615 ( .DIN1(n8825), .DIN2(n8826), .Q(n5943) );
  nnd2s1 U9616 ( .DIN1(n8325), .DIN2(n789), .Q(n8826) );
  and2s1 U9617 ( .DIN1(n8827), .DIN2(n8828), .Q(n6814) );
  nnd2s1 U9618 ( .DIN1(n544), .DIN2(n8328), .Q(n8828) );
  nnd2s1 U9619 ( .DIN1(n554), .DIN2(n8330), .Q(n8827) );
  nnd4s1 U9620 ( .DIN1(n7193), .DIN2(n8829), .DIN3(n8830), .DIN4(n8831), 
        .Q(n8786) );
  or2s1 U9621 ( .DIN1(n8311), .DIN2(n6465), .Q(n8831) );
  nnd2s1 U9622 ( .DIN1(n8170), .DIN2(n707), .Q(n8311) );
  nor2s1 U9623 ( .DIN1(n6380), .DIN2(n5321), .Q(n8170) );
  nor2s1 U9624 ( .DIN1(n803), .DIN2(n401), .Q(n5321) );
  hi1s1 U9625 ( .DIN(n7205), .Q(n6380) );
  nnd2s1 U9626 ( .DIN1(n7836), .DIN2(n8832), .Q(n8830) );
  nnd3s1 U9627 ( .DIN1(n8833), .DIN2(n8834), .DIN3(n8835), .Q(n8832) );
  nnd2s1 U9628 ( .DIN1(n5951), .DIN2(n735), .Q(n8835) );
  hi1s1 U9629 ( .DIN(n6816), .Q(n5951) );
  nnd2s1 U9630 ( .DIN1(n8825), .DIN2(n8836), .Q(n6816) );
  nnd2s1 U9631 ( .DIN1(n8325), .DIN2(n213), .Q(n8836) );
  nor2s1 U9632 ( .DIN1(n62), .DIN2(n746), .Q(n8325) );
  and2s1 U9633 ( .DIN1(n8837), .DIN2(n8838), .Q(n8825) );
  nnd2s1 U9634 ( .DIN1(n5546), .DIN2(n4845), .Q(n8838) );
  nor2s1 U9635 ( .DIN1(n717), .DIN2(n213), .Q(n5546) );
  nnd2s1 U9636 ( .DIN1(n747), .DIN2(n7355), .Q(n8837) );
  nnd4s1 U9637 ( .DIN1(n5962), .DIN2(n5731), .DIN3(n8839), .DIN4(n5544), 
        .Q(n7355) );
  nnd2s1 U9638 ( .DIN1(n784), .DIN2(n434), .Q(n5544) );
  nnd2s1 U9639 ( .DIN1(n758), .DIN2(n406), .Q(n8839) );
  nnd2s1 U9640 ( .DIN1(n789), .DIN2(n407), .Q(n5731) );
  nnd2s1 U9641 ( .DIN1(n553), .DIN2(n435), .Q(n5962) );
  nnd2s1 U9642 ( .DIN1(n6386), .DIN2(n545), .Q(n8834) );
  hi1s1 U9643 ( .DIN(n8328), .Q(n6386) );
  nnd4s1 U9644 ( .DIN1(n6395), .DIN2(n6177), .DIN3(n5732), .DIN4(n8840), 
        .Q(n8328) );
  nnd2s1 U9645 ( .DIN1(n783), .DIN2(n409), .Q(n8840) );
  nnd2s1 U9646 ( .DIN1(n759), .DIN2(n408), .Q(n5732) );
  nnd2s1 U9647 ( .DIN1(n790), .DIN2(n410), .Q(n6177) );
  nnd2s1 U9648 ( .DIN1(n552), .DIN2(n411), .Q(n6395) );
  nnd2s1 U9649 ( .DIN1(n7356), .DIN2(n555), .Q(n8833) );
  hi1s1 U9650 ( .DIN(n8330), .Q(n7356) );
  nnd4s1 U9651 ( .DIN1(n6824), .DIN2(n6605), .DIN3(n8841), .DIN4(n6398), 
        .Q(n8330) );
  nnd2s1 U9652 ( .DIN1(n784), .DIN2(n413), .Q(n6398) );
  nnd2s1 U9653 ( .DIN1(n759), .DIN2(n412), .Q(n8841) );
  nnd2s1 U9654 ( .DIN1(n789), .DIN2(n414), .Q(n6605) );
  nnd2s1 U9655 ( .DIN1(n553), .DIN2(n415), .Q(n6824) );
  nnd2s1 U9656 ( .DIN1(n9486), .DIN2(n8823), .Q(n8829) );
  nnd3s1 U9657 ( .DIN1(n8842), .DIN2(n8843), .DIN3(n8844), .Q(n8823) );
  nnd4s1 U9658 ( .DIN1(n8845), .DIN2(n8846), .DIN3(n740), .DIN4(n8847), 
        .Q(n8844) );
  nor2s1 U9659 ( .DIN1(n8848), .DIN2(n802), .Q(n8847) );
  nor2s1 U9660 ( .DIN1(n29), .DIN2(n8304), .Q(n8848) );
  nnd3s1 U9661 ( .DIN1(n8849), .DIN2(n8850), .DIN3(n707), .Q(n8304) );
  nnd2s1 U9662 ( .DIN1(n9489), .DIN2(n332), .Q(n8850) );
  nnd2s1 U9663 ( .DIN1(n440), .DIN2(n66), .Q(n8849) );
  nnd2s1 U9664 ( .DIN1(n8716), .DIN2(n439), .Q(n8846) );
  nnd2s1 U9665 ( .DIN1(n8851), .DIN2(n8852), .Q(n8716) );
  nnd3s1 U9666 ( .DIN1(n429), .DIN2(n712), .DIN3(n4845), .Q(n8852) );
  nnd2s1 U9667 ( .DIN1(n8853), .DIN2(n29), .Q(n8851) );
  nnd2s1 U9668 ( .DIN1(n8854), .DIN2(n8855), .Q(n8853) );
  nnd2s1 U9669 ( .DIN1(n428), .DIN2(n707), .Q(n8855) );
  nnd2s1 U9670 ( .DIN1(n431), .DIN2(n712), .Q(n8854) );
  nnd2s1 U9671 ( .DIN1(n8856), .DIN2(n9489), .Q(n8845) );
  nnd2s1 U9672 ( .DIN1(n7834), .DIN2(n5315), .Q(n8843) );
  hi1s1 U9673 ( .DIN(n8331), .Q(n7834) );
  nnd4s1 U9674 ( .DIN1(n7814), .DIN2(n7576), .DIN3(n7022), .DIN4(n7337), 
        .Q(n8331) );
  nnd2s1 U9675 ( .DIN1(n783), .DIN2(n421), .Q(n7337) );
  nnd2s1 U9676 ( .DIN1(n758), .DIN2(n420), .Q(n7022) );
  nnd2s1 U9677 ( .DIN1(n790), .DIN2(n422), .Q(n7576) );
  nnd2s1 U9678 ( .DIN1(n552), .DIN2(n423), .Q(n7814) );
  nnd2s1 U9679 ( .DIN1(n7357), .DIN2(n719), .Q(n8842) );
  hi1s1 U9680 ( .DIN(n8319), .Q(n7357) );
  nnd4s1 U9681 ( .DIN1(n7334), .DIN2(n7021), .DIN3(n6606), .DIN4(n6827), 
        .Q(n8319) );
  nnd2s1 U9682 ( .DIN1(n784), .DIN2(n417), .Q(n6827) );
  nnd2s1 U9683 ( .DIN1(n759), .DIN2(n416), .Q(n6606) );
  nnd2s1 U9684 ( .DIN1(n789), .DIN2(n418), .Q(n7021) );
  nnd2s1 U9685 ( .DIN1(n553), .DIN2(n419), .Q(n7334) );
  nnd3s1 U9686 ( .DIN1(n8857), .DIN2(n8858), .DIN3(n8859), .Q(\EXinst/n1433 )
         );
  nnd2s1 U9687 ( .DIN1(n727), .DIN2(\DM_addr[1] ), .Q(n8859) );
  nnd2s1 U9688 ( .DIN1(n5324), .DIN2(n8860), .Q(n8858) );
  nnd4s1 U9689 ( .DIN1(n8861), .DIN2(n8862), .DIN3(n8863), .DIN4(n8864), 
        .Q(n8860) );
  and4s1 U9690 ( .DIN1(n8865), .DIN2(n8866), .DIN3(n8867), .DIN4(n8868), 
        .Q(n8864) );
  nnd2s1 U9691 ( .DIN1(n8869), .DIN2(n8870), .Q(n8868) );
  nnd3s1 U9692 ( .DIN1(n8871), .DIN2(n749), .DIN3(n8872), .Q(n8870) );
  nnd2s1 U9693 ( .DIN1(n705), .DIN2(n8873), .Q(n8872) );
  nnd2s1 U9694 ( .DIN1(n655), .DIN2(n8742), .Q(n8871) );
  nnd2s1 U9695 ( .DIN1(n399), .DIN2(n33), .Q(n8742) );
  nnd2s1 U9696 ( .DIN1(n8874), .DIN2(n8875), .Q(n8867) );
  nnd2s1 U9697 ( .DIN1(n8876), .DIN2(n8877), .Q(n8875) );
  nnd3s1 U9698 ( .DIN1(n399), .DIN2(n430), .DIN3(n654), .Q(n8877) );
  nnd2s1 U9699 ( .DIN1(n620), .DIN2(n8878), .Q(n8876) );
  hi1s1 U9700 ( .DIN(n8869), .Q(n8874) );
  nnd2s1 U9701 ( .DIN1(n7138), .DIN2(n6963), .Q(n8866) );
  and4s1 U9702 ( .DIN1(n629), .DIN2(n8879), .DIN3(n8873), .DIN4(n714), 
        .Q(n6963) );
  nnd2s1 U9703 ( .DIN1(n330), .DIN2(n1), .Q(n8879) );
  nnd2s1 U9704 ( .DIN1(n35), .DIN2(n767), .Q(n8865) );
  nnd2s1 U9705 ( .DIN1(reg_out_B[1]), .DIN2(n8880), .Q(n8863) );
  nnd2s1 U9706 ( .DIN1(n5471), .DIN2(n8881), .Q(n8880) );
  nnd2s1 U9707 ( .DIN1(n776), .DIN2(n432), .Q(n8881) );
  nnd3s1 U9708 ( .DIN1(n8882), .DIN2(n8883), .DIN3(n5336), .Q(n8862) );
  nnd3s1 U9709 ( .DIN1(n8884), .DIN2(n8885), .DIN3(n5337), .Q(n8883) );
  nnd2s1 U9710 ( .DIN1(n753), .DIN2(n6948), .Q(n8885) );
  nnd2s1 U9711 ( .DIN1(n8886), .DIN2(n8887), .Q(n6948) );
  nnd3s1 U9712 ( .DIN1(n8888), .DIN2(n7895), .DIN3(n438), .Q(n8887) );
  nnd2s1 U9713 ( .DIN1(n8889), .DIN2(n5490), .Q(n7895) );
  hi1s1 U9714 ( .DIN(n7413), .Q(n8889) );
  nnd2s1 U9715 ( .DIN1(n8391), .DIN2(n32), .Q(n8888) );
  hi1s1 U9716 ( .DIN(n5651), .Q(n8391) );
  nnd2s1 U9717 ( .DIN1(n8890), .DIN2(n8891), .Q(n5651) );
  nnd2s1 U9718 ( .DIN1(n715), .DIN2(n734), .Q(n8891) );
  nnd3s1 U9719 ( .DIN1(n8892), .DIN2(n8893), .DIN3(n808), .Q(n8884) );
  or3s1 U9720 ( .DIN1(n7089), .DIN2(n7156), .DIN3(n6087), .Q(n8882) );
  nnd2s1 U9721 ( .DIN1(n8894), .DIN2(n6863), .Q(n6087) );
  hi1s1 U9722 ( .DIN(n7283), .Q(n6863) );
  nor2s1 U9723 ( .DIN1(n401), .DIN2(n741), .Q(n7283) );
  nnd2s1 U9724 ( .DIN1(n734), .DIN2(n211), .Q(n8894) );
  nor2s1 U9725 ( .DIN1(n62), .DIN2(n61), .Q(n7156) );
  nnd2s1 U9726 ( .DIN1(n716), .DIN2(n8895), .Q(n7089) );
  nnd2s1 U9727 ( .DIN1(n734), .DIN2(n204), .Q(n8895) );
  nnd2s1 U9728 ( .DIN1(n8896), .DIN2(n8897), .Q(n8861) );
  nnd2s1 U9729 ( .DIN1(n808), .DIN2(n8898), .Q(n8897) );
  nnd2s1 U9730 ( .DIN1(n8892), .DIN2(n8893), .Q(n8898) );
  nnd3s1 U9731 ( .DIN1(n8899), .DIN2(n8900), .DIN3(n801), .Q(n8893) );
  nnd2s1 U9732 ( .DIN1(n32), .DIN2(n8368), .Q(n8900) );
  nnd3s1 U9733 ( .DIN1(n8105), .DIN2(n8901), .DIN3(n8374), .Q(n8368) );
  nnd2s1 U9734 ( .DIN1(n755), .DIN2(n428), .Q(n8374) );
  nnd3s1 U9735 ( .DIN1(n8902), .DIN2(n8903), .DIN3(reg_out_B[1]), .Q(n8901) );
  nnd2s1 U9736 ( .DIN1(n399), .DIN2(n332), .Q(n8903) );
  nnd2s1 U9737 ( .DIN1(n63), .DIN2(n1), .Q(n8902) );
  nnd2s1 U9738 ( .DIN1(n774), .DIN2(n427), .Q(n8105) );
  nnd2s1 U9739 ( .DIN1(n8904), .DIN2(n5490), .Q(n8899) );
  nnd4s1 U9740 ( .DIN1(n8378), .DIN2(n8618), .DIN3(n8106), .DIN4(n8377), 
        .Q(n8904) );
  nnd2s1 U9741 ( .DIN1(n772), .DIN2(n431), .Q(n8377) );
  nnd2s1 U9742 ( .DIN1(n532), .DIN2(n433), .Q(n8106) );
  nnd2s1 U9743 ( .DIN1(n773), .DIN2(n426), .Q(n8618) );
  nnd2s1 U9744 ( .DIN1(n754), .DIN2(n35), .Q(n8378) );
  nnd3s1 U9745 ( .DIN1(n8905), .DIN2(n8906), .DIN3(n61), .Q(n8892) );
  nnd2s1 U9746 ( .DIN1(n741), .DIN2(n7404), .Q(n8906) );
  nnd4s1 U9747 ( .DIN1(n7390), .DIN2(n7145), .DIN3(n6741), .DIN4(n6961), 
        .Q(n7404) );
  nnd2s1 U9748 ( .DIN1(n771), .DIN2(n418), .Q(n6961) );
  nnd2s1 U9749 ( .DIN1(n531), .DIN2(n417), .Q(n6741) );
  nnd2s1 U9750 ( .DIN1(n774), .DIN2(n419), .Q(n7145) );
  nnd2s1 U9751 ( .DIN1(n755), .DIN2(n420), .Q(n7390) );
  nnd2s1 U9752 ( .DIN1(n7884), .DIN2(n5490), .Q(n8905) );
  nnd4s1 U9753 ( .DIN1(n7869), .DIN2(n7640), .DIN3(n7146), .DIN4(n7393), 
        .Q(n7884) );
  nnd2s1 U9754 ( .DIN1(n772), .DIN2(n422), .Q(n7393) );
  nnd2s1 U9755 ( .DIN1(n532), .DIN2(n421), .Q(n7146) );
  nnd2s1 U9756 ( .DIN1(n773), .DIN2(n423), .Q(n7640) );
  nnd2s1 U9757 ( .DIN1(n754), .DIN2(n424), .Q(n7869) );
  nnd2s1 U9758 ( .DIN1(n5994), .DIN2(n8907), .Q(n8896) );
  nnd2s1 U9759 ( .DIN1(n386), .DIN2(n6942), .Q(n8907) );
  nnd3s1 U9760 ( .DIN1(n8908), .DIN2(n8909), .DIN3(n8886), .Q(n6942) );
  and2s1 U9761 ( .DIN1(n8910), .DIN2(n8911), .Q(n8886) );
  nnd2s1 U9762 ( .DIN1(n622), .DIN2(n7414), .Q(n8911) );
  nnd4s1 U9763 ( .DIN1(n6525), .DIN2(n6311), .DIN3(n5879), .DIN4(n8912), 
        .Q(n7414) );
  nnd2s1 U9764 ( .DIN1(n771), .DIN2(n410), .Q(n8912) );
  nnd2s1 U9765 ( .DIN1(n531), .DIN2(n409), .Q(n5879) );
  nnd2s1 U9766 ( .DIN1(n774), .DIN2(n411), .Q(n6311) );
  nnd2s1 U9767 ( .DIN1(n755), .DIN2(n412), .Q(n6525) );
  nnd2s1 U9768 ( .DIN1(n628), .DIN2(n7412), .Q(n8910) );
  nnd4s1 U9769 ( .DIN1(n6958), .DIN2(n6740), .DIN3(n6312), .DIN4(n6528), 
        .Q(n7412) );
  nnd2s1 U9770 ( .DIN1(n772), .DIN2(n414), .Q(n6528) );
  nnd2s1 U9771 ( .DIN1(n532), .DIN2(n413), .Q(n6312) );
  nnd2s1 U9772 ( .DIN1(n773), .DIN2(n415), .Q(n6740) );
  nnd2s1 U9773 ( .DIN1(n754), .DIN2(n416), .Q(n6958) );
  nnd2s1 U9774 ( .DIN1(n5876), .DIN2(n5654), .Q(n8909) );
  nnd2s1 U9775 ( .DIN1(n8890), .DIN2(n8913), .Q(n5654) );
  nnd2s1 U9776 ( .DIN1(n771), .DIN2(n734), .Q(n8913) );
  and2s1 U9777 ( .DIN1(n5636), .DIN2(n8914), .Q(n8890) );
  nnd2s1 U9778 ( .DIN1(n718), .DIN2(n774), .Q(n8914) );
  nnd2s1 U9779 ( .DIN1(n755), .DIN2(n406), .Q(n5636) );
  nnd2s1 U9780 ( .DIN1(n547), .DIN2(n7413), .Q(n8908) );
  nnd4s1 U9781 ( .DIN1(n6098), .DIN2(n5878), .DIN3(n8915), .DIN4(n5639), 
        .Q(n7413) );
  nnd2s1 U9782 ( .DIN1(n772), .DIN2(n407), .Q(n5639) );
  nnd2s1 U9783 ( .DIN1(n531), .DIN2(n12), .Q(n8915) );
  nnd2s1 U9784 ( .DIN1(n774), .DIN2(n435), .Q(n5878) );
  nnd2s1 U9785 ( .DIN1(n754), .DIN2(n408), .Q(n6098) );
  nnd2s1 U9786 ( .DIN1(n551), .DIN2(n8916), .Q(n8857) );
  nnd4s1 U9787 ( .DIN1(n8917), .DIN2(n8918), .DIN3(n8919), .DIN4(n8920), 
        .Q(n8916) );
  and3s1 U9788 ( .DIN1(n8921), .DIN2(n8922), .DIN3(n8923), .Q(n8920) );
  nnd2s1 U9789 ( .DIN1(n7206), .DIN2(n707), .Q(n8923) );
  nnd2s1 U9790 ( .DIN1(n432), .DIN2(n8924), .Q(n8922) );
  nnd4s1 U9791 ( .DIN1(n8925), .DIN2(n8926), .DIN3(n8927), .DIN4(n7059), 
        .Q(n8924) );
  nnd2s1 U9792 ( .DIN1(n8928), .DIN2(n7212), .Q(n8927) );
  xnr2s1 U9793 ( .DIN1(n8809), .DIN2(n8810), .Q(n8928) );
  hi1s1 U9794 ( .DIN(n8929), .Q(n8810) );
  nnd2s1 U9795 ( .DIN1(n8930), .DIN2(n743), .Q(n8926) );
  xnr2s1 U9796 ( .DIN1(n8815), .DIN2(n8816), .Q(n8930) );
  hi1s1 U9797 ( .DIN(n8931), .Q(n8816) );
  nor2s1 U9798 ( .DIN1(n8932), .DIN2(n8933), .Q(n8925) );
  nor2s1 U9799 ( .DIN1(n711), .DIN2(n7006), .Q(n8933) );
  nor2s1 U9800 ( .DIN1(n712), .DIN2(n7037), .Q(n8932) );
  nnd2s1 U9801 ( .DIN1(n8934), .DIN2(n330), .Q(n8921) );
  nnd3s1 U9802 ( .DIN1(n8935), .DIN2(n8936), .DIN3(n8937), .Q(n8934) );
  nnd2s1 U9803 ( .DIN1(n7222), .DIN2(n707), .Q(n8937) );
  hi1s1 U9804 ( .DIN(n7006), .Q(n7222) );
  nnd2s1 U9805 ( .DIN1(n8938), .DIN2(n722), .Q(n8936) );
  xnr2s1 U9806 ( .DIN1(n8809), .DIN2(n8929), .Q(n8938) );
  xnr2s1 U9807 ( .DIN1(n712), .DIN2(n785), .Q(n8929) );
  nnd2s1 U9808 ( .DIN1(n8939), .DIN2(n8940), .Q(n8809) );
  nnd2s1 U9809 ( .DIN1(n430), .DIN2(n8941), .Q(n8940) );
  nnd2s1 U9810 ( .DIN1(n8942), .DIN2(n785), .Q(n8941) );
  or2s1 U9811 ( .DIN1(n8942), .DIN2(n5514), .Q(n8939) );
  nnd2s1 U9812 ( .DIN1(n8943), .DIN2(n7058), .Q(n8935) );
  xnr2s1 U9813 ( .DIN1(n8815), .DIN2(n8931), .Q(n8943) );
  xnr2s1 U9814 ( .DIN1(n5423), .DIN2(n711), .Q(n8931) );
  nnd2s1 U9815 ( .DIN1(n8944), .DIN2(n8945), .Q(n8815) );
  nnd2s1 U9816 ( .DIN1(n33), .DIN2(n8946), .Q(n8945) );
  nnd2s1 U9817 ( .DIN1(n8947), .DIN2(n5426), .Q(n8946) );
  or2s1 U9818 ( .DIN1(n8947), .DIN2(n5426), .Q(n8944) );
  nnd2s1 U9819 ( .DIN1(n400), .DIN2(n6913), .Q(n8919) );
  and3s1 U9820 ( .DIN1(n8948), .DIN2(n8949), .DIN3(n7345), .Q(n6913) );
  nor2s1 U9821 ( .DIN1(n6253), .DIN2(n711), .Q(n7345) );
  hi1s1 U9822 ( .DIN(n554), .Q(n6253) );
  nnd2s1 U9823 ( .DIN1(n9489), .DIN2(n330), .Q(n8949) );
  nnd2s1 U9824 ( .DIN1(n439), .DIN2(n331), .Q(n8948) );
  nnd3s1 U9825 ( .DIN1(n7339), .DIN2(n8951), .DIN3(n8952), .Q(n8918) );
  hi1s1 U9826 ( .DIN(n8953), .Q(n8952) );
  or2s1 U9827 ( .DIN1(n6915), .DIN2(n740), .Q(n8951) );
  nnd3s1 U9828 ( .DIN1(n8954), .DIN2(n8955), .DIN3(n6893), .Q(n6915) );
  and2s1 U9829 ( .DIN1(n8956), .DIN2(n8957), .Q(n6893) );
  nnd2s1 U9830 ( .DIN1(n545), .DIN2(n7454), .Q(n8957) );
  nnd2s1 U9831 ( .DIN1(n555), .DIN2(n7455), .Q(n8956) );
  nnd2s1 U9832 ( .DIN1(n5824), .DIN2(n5569), .Q(n8955) );
  nnd2s1 U9833 ( .DIN1(n8958), .DIN2(n8959), .Q(n5569) );
  nnd2s1 U9834 ( .DIN1(n783), .DIN2(n734), .Q(n8959) );
  nnd2s1 U9835 ( .DIN1(n5826), .DIN2(n7452), .Q(n8954) );
  and3s1 U9836 ( .DIN1(n8960), .DIN2(n4878), .DIN3(n6036), .Q(n7339) );
  nnd4s1 U9837 ( .DIN1(n7193), .DIN2(n8961), .DIN3(n8962), .DIN4(n8963), 
        .Q(n8917) );
  nnd3s1 U9838 ( .DIN1(n8964), .DIN2(n6894), .DIN3(n7836), .Q(n8963) );
  nnd3s1 U9839 ( .DIN1(n7919), .DIN2(n8965), .DIN3(n735), .Q(n6894) );
  nnd2s1 U9840 ( .DIN1(n8438), .DIN2(n4845), .Q(n8965) );
  hi1s1 U9841 ( .DIN(n5575), .Q(n8438) );
  nnd2s1 U9842 ( .DIN1(n8958), .DIN2(n8966), .Q(n5575) );
  nnd2s1 U9843 ( .DIN1(n734), .DIN2(n707), .Q(n8966) );
  and2s1 U9844 ( .DIN1(n5593), .DIN2(n8967), .Q(n8958) );
  nnd2s1 U9845 ( .DIN1(n718), .DIN2(n790), .Q(n8967) );
  nnd2s1 U9846 ( .DIN1(n552), .DIN2(n406), .Q(n5593) );
  nnd2s1 U9847 ( .DIN1(n7439), .DIN2(n747), .Q(n7919) );
  hi1s1 U9848 ( .DIN(n7452), .Q(n7439) );
  nnd4s1 U9849 ( .DIN1(n6047), .DIN2(n5820), .DIN3(n8968), .DIN4(n5596), 
        .Q(n7452) );
  nnd2s1 U9850 ( .DIN1(n784), .DIN2(n407), .Q(n5596) );
  nnd2s1 U9851 ( .DIN1(n759), .DIN2(n434), .Q(n8968) );
  nnd2s1 U9852 ( .DIN1(n790), .DIN2(n6), .Q(n5820) );
  nnd2s1 U9853 ( .DIN1(n553), .DIN2(n408), .Q(n6047) );
  nnd3s1 U9854 ( .DIN1(n8969), .DIN2(n8970), .DIN3(n736), .Q(n8964) );
  nnd2s1 U9855 ( .DIN1(n7440), .DIN2(n4845), .Q(n8970) );
  hi1s1 U9856 ( .DIN(n7454), .Q(n7440) );
  nnd4s1 U9857 ( .DIN1(n6475), .DIN2(n6255), .DIN3(n5821), .DIN4(n8971), 
        .Q(n7454) );
  nnd2s1 U9858 ( .DIN1(n783), .DIN2(n410), .Q(n8971) );
  nnd2s1 U9859 ( .DIN1(n758), .DIN2(n409), .Q(n5821) );
  nnd2s1 U9860 ( .DIN1(n789), .DIN2(n411), .Q(n6255) );
  nnd2s1 U9861 ( .DIN1(n552), .DIN2(n412), .Q(n6475) );
  nnd2s1 U9862 ( .DIN1(n7441), .DIN2(n29), .Q(n8969) );
  hi1s1 U9863 ( .DIN(n7455), .Q(n7441) );
  nnd4s1 U9864 ( .DIN1(n6907), .DIN2(n6683), .DIN3(n6256), .DIN4(n6478), 
        .Q(n7455) );
  nnd2s1 U9865 ( .DIN1(n784), .DIN2(n414), .Q(n6478) );
  nnd2s1 U9866 ( .DIN1(n759), .DIN2(n413), .Q(n6256) );
  nnd2s1 U9867 ( .DIN1(n790), .DIN2(n415), .Q(n6683) );
  nnd2s1 U9868 ( .DIN1(n553), .DIN2(n416), .Q(n6907) );
  or2s1 U9869 ( .DIN1(n6034), .DIN2(n7196), .Q(n8962) );
  nnd2s1 U9870 ( .DIN1(n7205), .DIN2(n803), .Q(n7196) );
  nor2s1 U9871 ( .DIN1(n56), .DIN2(n733), .Q(n7205) );
  nnd2s1 U9872 ( .DIN1(n8972), .DIN2(n5741), .Q(n6034) );
  hi1s1 U9873 ( .DIN(n6465), .Q(n5741) );
  nor2s1 U9874 ( .DIN1(n4845), .DIN2(n62), .Q(n6465) );
  nnd2s1 U9875 ( .DIN1(n734), .DIN2(n5313), .Q(n8972) );
  nnd2s1 U9876 ( .DIN1(n733), .DIN2(n8953), .Q(n8961) );
  nnd3s1 U9877 ( .DIN1(n8973), .DIN2(n8974), .DIN3(n8975), .Q(n8953) );
  nnd4s1 U9878 ( .DIN1(n8976), .DIN2(n739), .DIN3(n9487), .DIN4(n8977), 
        .Q(n8975) );
  nnd2s1 U9879 ( .DIN1(n8856), .DIN2(n440), .Q(n8977) );
  nnd2s1 U9880 ( .DIN1(n8978), .DIN2(n8979), .Q(n8856) );
  nnd2s1 U9881 ( .DIN1(n712), .DIN2(n8980), .Q(n8979) );
  nnd2s1 U9882 ( .DIN1(n8981), .DIN2(n8982), .Q(n8980) );
  nnd2s1 U9883 ( .DIN1(n34), .DIN2(n4845), .Q(n8982) );
  nnd3s1 U9884 ( .DIN1(n10), .DIN2(n747), .DIN3(n707), .Q(n8978) );
  nor2s1 U9885 ( .DIN1(n8983), .DIN2(n8984), .Q(n8976) );
  nor2s1 U9886 ( .DIN1(n8985), .DIN2(n4845), .Q(n8984) );
  nor2s1 U9887 ( .DIN1(n8986), .DIN2(n8987), .Q(n8985) );
  nor2s1 U9888 ( .DIN1(n330), .DIN2(n213), .Q(n8987) );
  and2s1 U9889 ( .DIN1(n431), .DIN2(n783), .Q(n8986) );
  nor2s1 U9890 ( .DIN1(n747), .DIN2(n8434), .Q(n8983) );
  and2s1 U9891 ( .DIN1(n8420), .DIN2(n8407), .Q(n8434) );
  nnd2s1 U9892 ( .DIN1(n552), .DIN2(n428), .Q(n8407) );
  nnd2s1 U9893 ( .DIN1(n8154), .DIN2(n707), .Q(n8420) );
  and2s1 U9894 ( .DIN1(n8988), .DIN2(n8989), .Q(n8154) );
  nnd2s1 U9895 ( .DIN1(n9489), .DIN2(n63), .Q(n8989) );
  nnd2s1 U9896 ( .DIN1(n440), .DIN2(n332), .Q(n8988) );
  nnd2s1 U9897 ( .DIN1(n7918), .DIN2(n5315), .Q(n8974) );
  hi1s1 U9898 ( .DIN(n7202), .Q(n5315) );
  nnd2s1 U9899 ( .DIN1(n5949), .DIN2(n747), .Q(n7202) );
  hi1s1 U9900 ( .DIN(n7931), .Q(n7918) );
  nnd4s1 U9901 ( .DIN1(n7907), .DIN2(n7675), .DIN3(n7180), .DIN4(n7430), 
        .Q(n7931) );
  nnd2s1 U9902 ( .DIN1(n783), .DIN2(n422), .Q(n7430) );
  nnd2s1 U9903 ( .DIN1(n758), .DIN2(n421), .Q(n7180) );
  nnd2s1 U9904 ( .DIN1(n789), .DIN2(n423), .Q(n7675) );
  nnd2s1 U9905 ( .DIN1(n553), .DIN2(n424), .Q(n7907) );
  nnd2s1 U9906 ( .DIN1(n7438), .DIN2(n5304), .Q(n8973) );
  and2s1 U9907 ( .DIN1(n5949), .DIN2(n792), .Q(n5304) );
  nor2s1 U9908 ( .DIN1(n806), .DIN2(n9487), .Q(n5949) );
  hi1s1 U9909 ( .DIN(n7456), .Q(n7438) );
  nnd4s1 U9910 ( .DIN1(n7427), .DIN2(n7179), .DIN3(n6684), .DIN4(n6910), 
        .Q(n7456) );
  nnd2s1 U9911 ( .DIN1(n784), .DIN2(n418), .Q(n6910) );
  nnd2s1 U9912 ( .DIN1(n758), .DIN2(n417), .Q(n6684) );
  nnd2s1 U9913 ( .DIN1(n790), .DIN2(n419), .Q(n7179) );
  nnd2s1 U9914 ( .DIN1(n552), .DIN2(n420), .Q(n7427) );
  and2s1 U9915 ( .DIN1(n8990), .DIN2(n7594), .Q(n7193) );
  nnd4s1 U9916 ( .DIN1(n8991), .DIN2(n8992), .DIN3(n8993), .DIN4(n8994), 
        .Q(\EXinst/n1432 ) );
  and4s1 U9917 ( .DIN1(n8995), .DIN2(n8996), .DIN3(n8997), .DIN4(n8998), 
        .Q(n8994) );
  nnd4s1 U9918 ( .DIN1(n7003), .DIN2(n6036), .DIN3(n8999), .DIN4(n9000), 
        .Q(n8998) );
  nnd2s1 U9919 ( .DIN1(n7002), .DIN2(n806), .Q(n9000) );
  nnd2s1 U9920 ( .DIN1(n740), .DIN2(n9001), .Q(n8999) );
  hi1s1 U9921 ( .DIN(n6898), .Q(n6036) );
  and3s1 U9922 ( .DIN1(n4878), .DIN2(n551), .DIN3(n8960), .Q(n7003) );
  nnd4s1 U9923 ( .DIN1(n8990), .DIN2(n6035), .DIN3(n9002), .DIN4(n9003), 
        .Q(n8997) );
  nnd3s1 U9924 ( .DIN1(n740), .DIN2(n9001), .DIN3(n733), .Q(n9003) );
  nnd4s1 U9925 ( .DIN1(n9004), .DIN2(n9005), .DIN3(n9006), .DIN4(n9007), 
        .Q(n9001) );
  nnd2s1 U9926 ( .DIN1(n554), .DIN2(n9008), .Q(n9007) );
  nnd4s1 U9927 ( .DIN1(n9009), .DIN2(n9010), .DIN3(n9011), .DIN4(n9012), 
        .Q(n9008) );
  nnd2s1 U9928 ( .DIN1(n783), .DIN2(n80), .Q(n9012) );
  nnd2s1 U9929 ( .DIN1(n759), .DIN2(n77), .Q(n9011) );
  nnd2s1 U9930 ( .DIN1(n789), .DIN2(n330), .Q(n9010) );
  nnd2s1 U9931 ( .DIN1(n553), .DIN2(n331), .Q(n9009) );
  nnd2s1 U9932 ( .DIN1(n7586), .DIN2(n5824), .Q(n9006) );
  hi1s1 U9933 ( .DIN(n7604), .Q(n7586) );
  nnd4s1 U9934 ( .DIN1(n7575), .DIN2(n7335), .DIN3(n6826), .DIN4(n7023), 
        .Q(n7604) );
  nnd2s1 U9935 ( .DIN1(n784), .DIN2(n419), .Q(n7023) );
  nnd2s1 U9936 ( .DIN1(n758), .DIN2(n418), .Q(n6826) );
  nnd2s1 U9937 ( .DIN1(n790), .DIN2(n420), .Q(n7335) );
  nnd2s1 U9938 ( .DIN1(n552), .DIN2(n421), .Q(n7575) );
  nnd2s1 U9939 ( .DIN1(n8061), .DIN2(n726), .Q(n9005) );
  hi1s1 U9940 ( .DIN(n8072), .Q(n8061) );
  nnd4s1 U9941 ( .DIN1(n8050), .DIN2(n7815), .DIN3(n7336), .DIN4(n7578), 
        .Q(n8072) );
  nnd2s1 U9942 ( .DIN1(n783), .DIN2(n423), .Q(n7578) );
  nnd2s1 U9943 ( .DIN1(n758), .DIN2(n422), .Q(n7336) );
  nnd2s1 U9944 ( .DIN1(n789), .DIN2(n424), .Q(n7815) );
  nnd2s1 U9945 ( .DIN1(n553), .DIN2(n425), .Q(n8050) );
  nnd2s1 U9946 ( .DIN1(n8577), .DIN2(n544), .Q(n9004) );
  hi1s1 U9947 ( .DIN(n8569), .Q(n8577) );
  nnd4s1 U9948 ( .DIN1(n8583), .DIN2(n8293), .DIN3(n7816), .DIN4(n8053), 
        .Q(n8569) );
  nnd2s1 U9949 ( .DIN1(n784), .DIN2(n34), .Q(n8053) );
  nnd2s1 U9950 ( .DIN1(n759), .DIN2(n429), .Q(n7816) );
  nnd2s1 U9951 ( .DIN1(n790), .DIN2(n428), .Q(n8293) );
  nnd2s1 U9952 ( .DIN1(n552), .DIN2(n10), .Q(n8583) );
  nnd2s1 U9953 ( .DIN1(n7002), .DIN2(n7836), .Q(n9002) );
  nor2s1 U9954 ( .DIN1(n4831), .DIN2(n740), .Q(n7836) );
  hi1s1 U9955 ( .DIN(n7010), .Q(n7002) );
  nnd4s1 U9956 ( .DIN1(n9013), .DIN2(n9014), .DIN3(n9015), .DIN4(n9016), 
        .Q(n7010) );
  nnd2s1 U9957 ( .DIN1(n5824), .DIN2(n5742), .Q(n9016) );
  nnd4s1 U9958 ( .DIN1(n5730), .DIN2(n5542), .DIN3(n9017), .DIN4(n9018), 
        .Q(n5742) );
  nnd2s1 U9959 ( .DIN1(n718), .DIN2(n784), .Q(n9018) );
  nnd2s1 U9960 ( .DIN1(n759), .DIN2(n734), .Q(n9017) );
  nnd2s1 U9961 ( .DIN1(n789), .DIN2(n406), .Q(n5542) );
  nnd2s1 U9962 ( .DIN1(n553), .DIN2(n12), .Q(n5730) );
  nor2s1 U9963 ( .DIN1(n746), .DIN2(n9487), .Q(n5824) );
  nnd2s1 U9964 ( .DIN1(n5826), .DIN2(n7601), .Q(n9015) );
  nnd4s1 U9965 ( .DIN1(n6179), .DIN2(n5960), .DIN3(n5543), .DIN4(n5733), 
        .Q(n7601) );
  nnd2s1 U9966 ( .DIN1(n783), .DIN2(n435), .Q(n5733) );
  nnd2s1 U9967 ( .DIN1(n758), .DIN2(n407), .Q(n5543) );
  nnd2s1 U9968 ( .DIN1(n790), .DIN2(n408), .Q(n5960) );
  nnd2s1 U9969 ( .DIN1(n552), .DIN2(n409), .Q(n6179) );
  nor2s1 U9970 ( .DIN1(n4845), .DIN2(n9487), .Q(n5826) );
  nnd2s1 U9971 ( .DIN1(n544), .DIN2(n7602), .Q(n9014) );
  nnd4s1 U9972 ( .DIN1(n6604), .DIN2(n6396), .DIN3(n9019), .DIN4(n9020), 
        .Q(n7602) );
  nnd2s1 U9973 ( .DIN1(n784), .DIN2(n411), .Q(n9020) );
  nnd2s1 U9974 ( .DIN1(n759), .DIN2(n410), .Q(n9019) );
  nnd2s1 U9975 ( .DIN1(n789), .DIN2(n412), .Q(n6396) );
  nnd2s1 U9976 ( .DIN1(n553), .DIN2(n413), .Q(n6604) );
  nnd2s1 U9977 ( .DIN1(n555), .DIN2(n7603), .Q(n9013) );
  nnd4s1 U9978 ( .DIN1(n7020), .DIN2(n6825), .DIN3(n6397), .DIN4(n6607), 
        .Q(n7603) );
  nnd2s1 U9979 ( .DIN1(n783), .DIN2(n415), .Q(n6607) );
  nnd2s1 U9980 ( .DIN1(n759), .DIN2(n414), .Q(n6397) );
  nnd2s1 U9981 ( .DIN1(n790), .DIN2(n416), .Q(n6825) );
  nnd2s1 U9982 ( .DIN1(n552), .DIN2(n417), .Q(n7020) );
  and2s1 U9983 ( .DIN1(n7594), .DIN2(n550), .Q(n6035) );
  and2s1 U9984 ( .DIN1(n8960), .DIN2(n7000), .Q(n7594) );
  and2s1 U9985 ( .DIN1(n6379), .DIN2(n9021), .Q(n8990) );
  nnd2s1 U9986 ( .DIN1(n4831), .DIN2(n62), .Q(n9021) );
  nnd3s1 U9987 ( .DIN1(n7026), .DIN2(n554), .DIN3(n5299), .Q(n8996) );
  hi1s1 U9988 ( .DIN(n5547), .Q(n5299) );
  nnd2s1 U9989 ( .DIN1(n7004), .DIN2(n7027), .Q(n5547) );
  and2s1 U9990 ( .DIN1(n8950), .DIN2(n551), .Q(n7027) );
  and2s1 U9991 ( .DIN1(n8960), .DIN2(n9022), .Q(n8950) );
  and4s1 U9992 ( .DIN1(IR_opcode_field[4]), .DIN2(IR_opcode_field[2]), 
        .DIN3(n760), .DIN4(n117), .Q(n8960) );
  nor2s1 U9993 ( .DIN1(n6898), .DIN2(n206), .Q(n7004) );
  nnd2s1 U9994 ( .DIN1(n6379), .DIN2(n733), .Q(n6898) );
  nor4s1 U9995 ( .DIN1(n9023), .DIN2(n9024), .DIN3(n9025), .DIN4(n9026), 
        .Q(n6379) );
  nnd4s1 U9996 ( .DIN1(n9475), .DIN2(n9476), .DIN3(n9474), .DIN4(n9027), 
        .Q(n9026) );
  and3s1 U9997 ( .DIN1(n9478), .DIN2(n9479), .DIN3(n9477), .Q(n9027) );
  nnd4s1 U9998 ( .DIN1(n9481), .DIN2(n9482), .DIN3(n9480), .DIN4(n9028), 
        .Q(n9025) );
  and4s1 U9999 ( .DIN1(n9483), .DIN2(n9484), .DIN3(n9485), .DIN4(n9460), 
        .Q(n9028) );
  nnd4s1 U10000 ( .DIN1(n9462), .DIN2(n9463), .DIN3(n9461), .DIN4(n9029), 
        .Q(n9024) );
  and3s1 U10001 ( .DIN1(n9465), .DIN2(n9466), .DIN3(n9464), .Q(n9029) );
  nnd4s1 U10002 ( .DIN1(n9468), .DIN2(n9469), .DIN3(n9467), .DIN4(n9030), 
        .Q(n9023) );
  and4s1 U10003 ( .DIN1(n9470), .DIN2(n9471), .DIN3(n9472), .DIN4(n9473), 
        .Q(n9030) );
  nnd2s1 U10004 ( .DIN1(n9031), .DIN2(n385), .Q(n8995) );
  hi1s1 U10005 ( .DIN(n5290), .Q(n5404) );
  nnd2s1 U10006 ( .DIN1(n550), .DIN2(n7212), .Q(n5290) );
  nnd4s1 U10007 ( .DIN1(n9032), .DIN2(n9033), .DIN3(n9034), .DIN4(n788), 
        .Q(n7212) );
  nnd2s1 U10008 ( .DIN1(n9035), .DIN2(n40), .Q(n9034) );
  nnd2s1 U10009 ( .DIN1(n9022), .DIN2(n9036), .Q(n9033) );
  nnd2s1 U10010 ( .DIN1(n9037), .DIN2(n7000), .Q(n9032) );
  xor2s1 U10011 ( .DIN1(n9038), .DIN2(n8942), .Q(n9031) );
  xnr2s1 U10012 ( .DIN1(n9489), .DIN2(n5514), .Q(n8942) );
  xnr2s1 U10013 ( .DIN1(n33), .DIN2(n744), .Q(n9038) );
  hi1s1 U10014 ( .DIN(n786), .Q(n5413) );
  nnd2s1 U10015 ( .DIN1(n9036), .DIN2(n4878), .Q(n5514) );
  nnd2s1 U10016 ( .DIN1(n551), .DIN2(n9039), .Q(n8993) );
  nnd4s1 U10017 ( .DIN1(n9040), .DIN2(n9041), .DIN3(n9042), .DIN4(n9043), 
        .Q(n9039) );
  nnd4s1 U10018 ( .DIN1(n4866), .DIN2(IR_opcode_field[4]), .DIN3(n9044), 
        .DIN4(n9045), .Q(n9043) );
  nnd4s1 U10019 ( .DIN1(n9046), .DIN2(n9047), .DIN3(n9048), .DIN4(n39), 
        .Q(n9045) );
  nor2s1 U10020 ( .DIN1(n9049), .DIN2(n9050), .Q(n9048) );
  nor2s1 U10021 ( .DIN1(n9051), .DIN2(n9052), .Q(n9050) );
  and2s1 U10022 ( .DIN1(n9052), .DIN2(n9053), .Q(n9049) );
  nnd4s1 U10023 ( .DIN1(n9054), .DIN2(n9055), .DIN3(n9056), .DIN4(n9057), 
        .Q(n9052) );
  nor4s1 U10024 ( .DIN1(n9058), .DIN2(n9059), .DIN3(n9060), .DIN4(n9061), 
        .Q(n9057) );
  nnd4s1 U10025 ( .DIN1(n9062), .DIN2(n9063), .DIN3(n9064), .DIN4(n9065), 
        .Q(n9061) );
  and2s1 U10026 ( .DIN1(n9066), .DIN2(n9067), .Q(n9064) );
  nnd4s1 U10027 ( .DIN1(n9068), .DIN2(n9069), .DIN3(n9070), .DIN4(n9071), 
        .Q(n9060) );
  and3s1 U10028 ( .DIN1(n9072), .DIN2(n9073), .DIN3(n9074), .Q(n9071) );
  nnd4s1 U10029 ( .DIN1(n9075), .DIN2(n9076), .DIN3(n9077), .DIN4(n9078), 
        .Q(n9059) );
  and3s1 U10030 ( .DIN1(n9079), .DIN2(n9080), .DIN3(n9081), .Q(n9078) );
  nnd4s1 U10031 ( .DIN1(n9082), .DIN2(n9083), .DIN3(n9084), .DIN4(n9085), 
        .Q(n9058) );
  and3s1 U10032 ( .DIN1(n9086), .DIN2(n9087), .DIN3(n9088), .Q(n9085) );
  nor4s1 U10033 ( .DIN1(n9089), .DIN2(n9090), .DIN3(n8817), .DIN4(n5287), 
        .Q(n9056) );
  nnd2s1 U10034 ( .DIN1(n9091), .DIN2(n9092), .Q(n5287) );
  nnd3s1 U10035 ( .DIN1(n216), .DIN2(n8557), .DIN3(n9093), .Q(n9090) );
  xnr2s1 U10036 ( .DIN1(n330), .DIN2(n712), .Q(n9093) );
  nnd4s1 U10037 ( .DIN1(n8054), .DIN2(n7818), .DIN3(n8296), .DIN4(n9094), 
        .Q(n9089) );
  and3s1 U10038 ( .DIN1(n7338), .DIN2(n7005), .DIN3(n7579), .Q(n9094) );
  and4s1 U10039 ( .DIN1(n9095), .DIN2(n9096), .DIN3(n9097), .DIN4(n9098), 
        .Q(n9055) );
  and3s1 U10040 ( .DIN1(n9099), .DIN2(n9100), .DIN3(n5560), .Q(n9095) );
  nor4s1 U10041 ( .DIN1(n9101), .DIN2(n6806), .DIN3(n6376), .DIN4(n6591), 
        .Q(n9054) );
  hi1s1 U10042 ( .DIN(n9102), .Q(n6591) );
  hi1s1 U10043 ( .DIN(n9103), .Q(n6376) );
  hi1s1 U10044 ( .DIN(n9104), .Q(n6806) );
  nnd3s1 U10045 ( .DIN1(n6019), .DIN2(n5795), .DIN3(n6163), .Q(n9101) );
  nnd2s1 U10046 ( .DIN1(n4878), .DIN2(n9105), .Q(n9047) );
  nnd2s1 U10047 ( .DIN1(n7000), .DIN2(n9106), .Q(n9046) );
  nnd3s1 U10048 ( .DIN1(n9107), .DIN2(n9108), .DIN3(IR_opcode_field[2]), 
        .Q(n9044) );
  or2s1 U10049 ( .DIN1(n9105), .DIN2(n4884), .Q(n9108) );
  hi1s1 U10050 ( .DIN(n9053), .Q(n4884) );
  nnd2s1 U10051 ( .DIN1(n9092), .DIN2(n9109), .Q(n9105) );
  nnd2s1 U10052 ( .DIN1(n9110), .DIN2(n9091), .Q(n9109) );
  nnd2s1 U10053 ( .DIN1(n9111), .DIN2(n9112), .Q(n9110) );
  nnd3s1 U10054 ( .DIN1(n9113), .DIN2(n9082), .DIN3(n5560), .Q(n9112) );
  nnd3s1 U10055 ( .DIN1(n9114), .DIN2(n9083), .DIN3(n9115), .Q(n9113) );
  nnd2s1 U10056 ( .DIN1(n102), .DIN2(n335), .Q(n9115) );
  nnd3s1 U10057 ( .DIN1(n9116), .DIN2(n9087), .DIN3(n5795), .Q(n9114) );
  nnd3s1 U10058 ( .DIN1(n9117), .DIN2(n9084), .DIN3(n9118), .Q(n9116) );
  nnd2s1 U10059 ( .DIN1(n103), .DIN2(n336), .Q(n9118) );
  nnd3s1 U10060 ( .DIN1(n9119), .DIN2(n9088), .DIN3(n6019), .Q(n9117) );
  nnd3s1 U10061 ( .DIN1(n9120), .DIN2(n9086), .DIN3(n9121), .Q(n9119) );
  nnd2s1 U10062 ( .DIN1(n120), .DIN2(n30), .Q(n9121) );
  nnd3s1 U10063 ( .DIN1(n9122), .DIN2(n9075), .DIN3(n6163), .Q(n9120) );
  nnd3s1 U10064 ( .DIN1(n9123), .DIN2(n9076), .DIN3(n9124), .Q(n9122) );
  nnd2s1 U10065 ( .DIN1(n121), .DIN2(n67), .Q(n9124) );
  nnd3s1 U10066 ( .DIN1(n9125), .DIN2(n9080), .DIN3(n9103), .Q(n9123) );
  nnd3s1 U10067 ( .DIN1(n9126), .DIN2(n9077), .DIN3(n9127), .Q(n9125) );
  nnd2s1 U10068 ( .DIN1(n123), .DIN2(n69), .Q(n9127) );
  nnd3s1 U10069 ( .DIN1(n9128), .DIN2(n9081), .DIN3(n9102), .Q(n9126) );
  nnd3s1 U10070 ( .DIN1(n9129), .DIN2(n9079), .DIN3(n9130), .Q(n9128) );
  nnd2s1 U10071 ( .DIN1(n122), .DIN2(n70), .Q(n9130) );
  nnd3s1 U10072 ( .DIN1(n9131), .DIN2(n9072), .DIN3(n9104), .Q(n9129) );
  nnd3s1 U10073 ( .DIN1(n9132), .DIN2(n9073), .DIN3(n9133), .Q(n9131) );
  nnd2s1 U10074 ( .DIN1(n109), .DIN2(n71), .Q(n9133) );
  nnd3s1 U10075 ( .DIN1(n9134), .DIN2(n9097), .DIN3(n7005), .Q(n9132) );
  nnd3s1 U10076 ( .DIN1(n9135), .DIN2(n9062), .DIN3(n9136), .Q(n9134) );
  nnd2s1 U10077 ( .DIN1(n108), .DIN2(n31), .Q(n9136) );
  nnd3s1 U10078 ( .DIN1(n9137), .DIN2(n9096), .DIN3(n7338), .Q(n9135) );
  nnd3s1 U10079 ( .DIN1(n9138), .DIN2(n9098), .DIN3(n9139), .Q(n9137) );
  nnd2s1 U10080 ( .DIN1(n106), .DIN2(n64), .Q(n9139) );
  nnd3s1 U10081 ( .DIN1(n9140), .DIN2(n9099), .DIN3(n7579), .Q(n9138) );
  nnd3s1 U10082 ( .DIN1(n9141), .DIN2(n9100), .DIN3(n9142), .Q(n9140) );
  nnd2s1 U10083 ( .DIN1(n104), .DIN2(n65), .Q(n9142) );
  nnd3s1 U10084 ( .DIN1(n9143), .DIN2(n9069), .DIN3(n7818), .Q(n9141) );
  nnd3s1 U10085 ( .DIN1(n9144), .DIN2(n9074), .DIN3(n9145), .Q(n9143) );
  nnd2s1 U10086 ( .DIN1(n107), .DIN2(n332), .Q(n9145) );
  nnd3s1 U10087 ( .DIN1(n9146), .DIN2(n9070), .DIN3(n8054), .Q(n9144) );
  nnd3s1 U10088 ( .DIN1(n9147), .DIN2(n9068), .DIN3(n9148), .Q(n9146) );
  nnd2s1 U10089 ( .DIN1(n105), .DIN2(n333), .Q(n9148) );
  nnd3s1 U10090 ( .DIN1(n9149), .DIN2(n9067), .DIN3(n8296), .Q(n9147) );
  nnd3s1 U10091 ( .DIN1(n9150), .DIN2(n9066), .DIN3(n9151), .Q(n9149) );
  nnd2s1 U10092 ( .DIN1(n805), .DIN2(n334), .Q(n9151) );
  nnd3s1 U10093 ( .DIN1(n9152), .DIN2(n9063), .DIN3(n8557), .Q(n9150) );
  nnd3s1 U10094 ( .DIN1(n9153), .DIN2(n9065), .DIN3(n9154), .Q(n9152) );
  nnd4s1 U10095 ( .DIN1(n9155), .DIN2(n9156), .DIN3(n9157), .DIN4(n213), 
        .Q(n9153) );
  nnd2s1 U10096 ( .DIN1(n35), .DIN2(n9158), .Q(n9157) );
  nnd2s1 U10097 ( .DIN1(n758), .DIN2(n331), .Q(n9158) );
  nnd2s1 U10098 ( .DIN1(n712), .DIN2(n430), .Q(n9156) );
  nnd2s1 U10099 ( .DIN1(n96), .DIN2(n717), .Q(n9111) );
  or2s1 U10100 ( .DIN1(n9106), .DIN2(n9051), .Q(n9107) );
  hi1s1 U10101 ( .DIN(n9022), .Q(n9051) );
  nnd2s1 U10102 ( .DIN1(n9091), .DIN2(n9159), .Q(n9106) );
  nnd2s1 U10103 ( .DIN1(n9160), .DIN2(n9092), .Q(n9159) );
  nnd2s1 U10104 ( .DIN1(n734), .DIN2(n9460), .Q(n9092) );
  nnd2s1 U10105 ( .DIN1(n9161), .DIN2(n9162), .Q(n9160) );
  nnd3s1 U10106 ( .DIN1(n9163), .DIN2(n9083), .DIN3(n5560), .Q(n9162) );
  xnr2s1 U10107 ( .DIN1(n96), .DIN2(reg_out_A[30]), .Q(n5560) );
  nnd2s1 U10108 ( .DIN1(n14), .DIN2(n79), .Q(n9083) );
  nnd3s1 U10109 ( .DIN1(n9164), .DIN2(n9082), .DIN3(n9165), .Q(n9163) );
  nnd2s1 U10110 ( .DIN1(n434), .DIN2(n9463), .Q(n9165) );
  nnd2s1 U10111 ( .DIN1(n406), .DIN2(n9462), .Q(n9082) );
  nnd3s1 U10112 ( .DIN1(n9166), .DIN2(n9084), .DIN3(n5795), .Q(n9164) );
  xnr2s1 U10113 ( .DIN1(n102), .DIN2(n434), .Q(n5795) );
  nnd2s1 U10114 ( .DIN1(n95), .DIN2(n38), .Q(n9084) );
  nnd3s1 U10115 ( .DIN1(n9167), .DIN2(n9087), .DIN3(n9168), .Q(n9166) );
  nnd2s1 U10116 ( .DIN1(n6), .DIN2(n9465), .Q(n9168) );
  nnd2s1 U10117 ( .DIN1(n407), .DIN2(n9464), .Q(n9087) );
  nnd3s1 U10118 ( .DIN1(n9169), .DIN2(n9086), .DIN3(n6019), .Q(n9167) );
  xnr2s1 U10119 ( .DIN1(n103), .DIN2(n6), .Q(n6019) );
  nnd2s1 U10120 ( .DIN1(n15), .DIN2(n83), .Q(n9086) );
  nnd3s1 U10121 ( .DIN1(n9170), .DIN2(n9088), .DIN3(n9171), .Q(n9169) );
  nnd2s1 U10122 ( .DIN1(n409), .DIN2(n9467), .Q(n9171) );
  nnd2s1 U10123 ( .DIN1(n408), .DIN2(n9466), .Q(n9088) );
  nnd3s1 U10124 ( .DIN1(n9172), .DIN2(n9076), .DIN3(n6163), .Q(n9170) );
  xnr2s1 U10125 ( .DIN1(n9467), .DIN2(n30), .Q(n6163) );
  nnd2s1 U10126 ( .DIN1(n93), .DIN2(n68), .Q(n9076) );
  nnd3s1 U10127 ( .DIN1(n9173), .DIN2(n9075), .DIN3(n9174), .Q(n9172) );
  nnd2s1 U10128 ( .DIN1(n411), .DIN2(n9469), .Q(n9174) );
  nnd2s1 U10129 ( .DIN1(n410), .DIN2(n9468), .Q(n9075) );
  nnd3s1 U10130 ( .DIN1(n9175), .DIN2(n9077), .DIN3(n9103), .Q(n9173) );
  xnr2s1 U10131 ( .DIN1(n9469), .DIN2(n67), .Q(n9103) );
  nnd2s1 U10132 ( .DIN1(n16), .DIN2(n78), .Q(n9077) );
  nnd3s1 U10133 ( .DIN1(n9176), .DIN2(n9080), .DIN3(n9177), .Q(n9175) );
  nnd2s1 U10134 ( .DIN1(n413), .DIN2(n9471), .Q(n9177) );
  nnd2s1 U10135 ( .DIN1(n412), .DIN2(n9470), .Q(n9080) );
  nnd3s1 U10136 ( .DIN1(n9178), .DIN2(n9079), .DIN3(n9102), .Q(n9176) );
  xnr2s1 U10137 ( .DIN1(n9471), .DIN2(n69), .Q(n9102) );
  nnd2s1 U10138 ( .DIN1(n94), .DIN2(n37), .Q(n9079) );
  nnd3s1 U10139 ( .DIN1(n9179), .DIN2(n9081), .DIN3(n9180), .Q(n9178) );
  nnd2s1 U10140 ( .DIN1(n415), .DIN2(n9473), .Q(n9180) );
  nnd2s1 U10141 ( .DIN1(n414), .DIN2(n9472), .Q(n9081) );
  nnd3s1 U10142 ( .DIN1(n9181), .DIN2(n9073), .DIN3(n9104), .Q(n9179) );
  xnr2s1 U10143 ( .DIN1(n9473), .DIN2(n70), .Q(n9104) );
  nnd2s1 U10144 ( .DIN1(n13), .DIN2(n82), .Q(n9073) );
  nnd3s1 U10145 ( .DIN1(n9182), .DIN2(n9072), .DIN3(n9183), .Q(n9181) );
  nnd2s1 U10146 ( .DIN1(n417), .DIN2(n9475), .Q(n9183) );
  nnd2s1 U10147 ( .DIN1(n416), .DIN2(n9474), .Q(n9072) );
  nnd3s1 U10148 ( .DIN1(n9184), .DIN2(n9062), .DIN3(n7005), .Q(n9182) );
  xnr2s1 U10149 ( .DIN1(n9475), .DIN2(n71), .Q(n7005) );
  nnd2s1 U10150 ( .DIN1(n7), .DIN2(n85), .Q(n9062) );
  nnd3s1 U10151 ( .DIN1(n9185), .DIN2(n9097), .DIN3(n9186), .Q(n9184) );
  nnd2s1 U10152 ( .DIN1(n419), .DIN2(n9477), .Q(n9186) );
  nnd2s1 U10153 ( .DIN1(n418), .DIN2(n9476), .Q(n9097) );
  nnd3s1 U10154 ( .DIN1(n9187), .DIN2(n9098), .DIN3(n7338), .Q(n9185) );
  xnr2s1 U10155 ( .DIN1(n9477), .DIN2(n31), .Q(n7338) );
  nnd2s1 U10156 ( .DIN1(n9), .DIN2(n86), .Q(n9098) );
  nnd3s1 U10157 ( .DIN1(n9188), .DIN2(n9096), .DIN3(n9189), .Q(n9187) );
  nnd2s1 U10158 ( .DIN1(n421), .DIN2(n9479), .Q(n9189) );
  nnd2s1 U10159 ( .DIN1(n420), .DIN2(n9478), .Q(n9096) );
  nnd3s1 U10160 ( .DIN1(n9190), .DIN2(n9100), .DIN3(n7579), .Q(n9188) );
  xnr2s1 U10161 ( .DIN1(n9479), .DIN2(n64), .Q(n7579) );
  nnd2s1 U10162 ( .DIN1(n8), .DIN2(n84), .Q(n9100) );
  nnd3s1 U10163 ( .DIN1(n9191), .DIN2(n9099), .DIN3(n9192), .Q(n9190) );
  nnd2s1 U10164 ( .DIN1(n423), .DIN2(n9481), .Q(n9192) );
  nnd2s1 U10165 ( .DIN1(n422), .DIN2(n9480), .Q(n9099) );
  nnd3s1 U10166 ( .DIN1(n9193), .DIN2(n9074), .DIN3(n7818), .Q(n9191) );
  xnr2s1 U10167 ( .DIN1(n9481), .DIN2(n65), .Q(n7818) );
  nnd2s1 U10168 ( .DIN1(n75), .DIN2(n66), .Q(n9074) );
  nnd3s1 U10169 ( .DIN1(n9194), .DIN2(n9069), .DIN3(n9195), .Q(n9193) );
  nnd2s1 U10170 ( .DIN1(n36), .DIN2(n9483), .Q(n9195) );
  nnd2s1 U10171 ( .DIN1(n424), .DIN2(n9482), .Q(n9069) );
  nnd3s1 U10172 ( .DIN1(n9196), .DIN2(n9068), .DIN3(n8054), .Q(n9194) );
  xnr2s1 U10173 ( .DIN1(n9483), .DIN2(n332), .Q(n8054) );
  nnd2s1 U10174 ( .DIN1(n76), .DIN2(n63), .Q(n9068) );
  nnd3s1 U10175 ( .DIN1(n9197), .DIN2(n9070), .DIN3(n9198), .Q(n9196) );
  nnd2s1 U10176 ( .DIN1(n427), .DIN2(n9485), .Q(n9198) );
  nnd2s1 U10177 ( .DIN1(n429), .DIN2(n9484), .Q(n9070) );
  nnd3s1 U10178 ( .DIN1(n9199), .DIN2(n9066), .DIN3(n8296), .Q(n9197) );
  xnr2s1 U10179 ( .DIN1(n9485), .DIN2(n333), .Q(n8296) );
  nnd2s1 U10180 ( .DIN1(n4831), .DIN2(n81), .Q(n9066) );
  hi1s1 U10181 ( .DIN(n733), .Q(n4831) );
  nnd3s1 U10182 ( .DIN1(n9200), .DIN2(n9067), .DIN3(n9201), .Q(n9199) );
  nnd2s1 U10183 ( .DIN1(n433), .DIN2(n740), .Q(n9201) );
  nnd2s1 U10184 ( .DIN1(n428), .DIN2(n9486), .Q(n9067) );
  nnd3s1 U10185 ( .DIN1(n9202), .DIN2(n9065), .DIN3(n8557), .Q(n9200) );
  xnr2s1 U10186 ( .DIN1(n433), .DIN2(n206), .Q(n8557) );
  nnd2s1 U10187 ( .DIN1(n803), .DIN2(n77), .Q(n9065) );
  hi1s1 U10188 ( .DIN(n736), .Q(n4840) );
  nnd3s1 U10189 ( .DIN1(n8981), .DIN2(n9063), .DIN3(n9203), .Q(n9202) );
  nnd4s1 U10190 ( .DIN1(n9155), .DIN2(n9204), .DIN3(n9205), .DIN4(n5313), 
        .Q(n9203) );
  or2s1 U10191 ( .DIN1(n7026), .DIN2(n35), .Q(n9205) );
  nor2s1 U10192 ( .DIN1(n213), .DIN2(n331), .Q(n7026) );
  nnd2s1 U10193 ( .DIN1(n707), .DIN2(n331), .Q(n9204) );
  hi1s1 U10194 ( .DIN(n8817), .Q(n9155) );
  nnd2s1 U10195 ( .DIN1(n8981), .DIN2(n9154), .Q(n8817) );
  nnd2s1 U10196 ( .DIN1(n4845), .DIN2(n80), .Q(n9154) );
  hi1s1 U10197 ( .DIN(n747), .Q(n4845) );
  nnd2s1 U10198 ( .DIN1(n431), .DIN2(n736), .Q(n9063) );
  nnd2s1 U10199 ( .DIN1(n426), .DIN2(n29), .Q(n8981) );
  nnd2s1 U10200 ( .DIN1(n718), .DIN2(n9461), .Q(n9161) );
  nnd2s1 U10201 ( .DIN1(n401), .DIN2(n124), .Q(n9091) );
  or2s1 U10202 ( .DIN1(n216), .DIN2(n7006), .Q(n9042) );
  nnd2s1 U10203 ( .DIN1(n7001), .DIN2(n4878), .Q(n7006) );
  nor2s1 U10204 ( .DIN1(n40), .DIN2(IR_opcode_field[0]), .Q(n4878) );
  nnd2s1 U10205 ( .DIN1(n7206), .DIN2(n439), .Q(n9041) );
  hi1s1 U10206 ( .DIN(n7059), .Q(n7206) );
  and2s1 U10207 ( .DIN1(n9206), .DIN2(n9207), .Q(n9040) );
  nnd2s1 U10208 ( .DIN1(n430), .DIN2(n9208), .Q(n9207) );
  nnd3s1 U10209 ( .DIN1(n9209), .DIN2(n7059), .DIN3(n9210), .Q(n9208) );
  nnd2s1 U10210 ( .DIN1(n7314), .DIN2(n440), .Q(n9210) );
  hi1s1 U10211 ( .DIN(n7037), .Q(n7314) );
  nnd2s1 U10212 ( .DIN1(n7001), .DIN2(n9022), .Q(n7037) );
  nnd2s1 U10213 ( .DIN1(n9053), .DIN2(n7001), .Q(n7059) );
  and3s1 U10214 ( .DIN1(IR_opcode_field[2]), .DIN2(n101), .DIN3(n4866), 
        .Q(n7001) );
  nnd2s1 U10215 ( .DIN1(n9211), .DIN2(n743), .Q(n9209) );
  nnd3s1 U10216 ( .DIN1(n381), .DIN2(n7058), .DIN3(n331), .Q(n9206) );
  nnd2s1 U10217 ( .DIN1(n5426), .DIN2(n9212), .Q(n7058) );
  nnd2s1 U10218 ( .DIN1(n9053), .DIN2(n9036), .Q(n9212) );
  xor2s1 U10219 ( .DIN1(n632), .DIN2(n8947), .Q(n9211) );
  xnr2s1 U10220 ( .DIN1(n633), .DIN2(n439), .Q(n8947) );
  hi1s1 U10221 ( .DIN(n5426), .Q(n5423) );
  nnd2s1 U10222 ( .DIN1(n7000), .DIN2(n9036), .Q(n5426) );
  and3s1 U10223 ( .DIN1(n39), .DIN2(n101), .DIN3(n4866), .Q(n9036) );
  nor2s1 U10224 ( .DIN1(n760), .DIN2(IR_opcode_field[5]), .Q(n4866) );
  nor2s1 U10225 ( .DIN1(n132), .DIN2(n40), .Q(n7000) );
  nnd2s1 U10226 ( .DIN1(n5394), .DIN2(\DM_addr[0] ), .Q(n8992) );
  nor2s1 U10227 ( .DIN1(n9213), .DIN2(n9214), .Q(n5394) );
  nnd4s1 U10228 ( .DIN1(n5324), .DIN2(n5469), .DIN3(n9215), .DIN4(n9216), 
        .Q(n9214) );
  nnd2s1 U10229 ( .DIN1(n9457), .DIN2(n9217), .Q(n9216) );
  nnd4s1 U10230 ( .DIN1(n9218), .DIN2(n5372), .DIN3(n9219), .DIN4(n9220), 
        .Q(n9213) );
  nnd2s1 U10231 ( .DIN1(n5324), .DIN2(n9221), .Q(n8991) );
  nnd4s1 U10232 ( .DIN1(n9222), .DIN2(n9223), .DIN3(n9224), .DIN4(n9225), 
        .Q(n9221) );
  and3s1 U10233 ( .DIN1(n9226), .DIN2(n9227), .DIN3(n9228), .Q(n9225) );
  nnd2s1 U10234 ( .DIN1(n5368), .DIN2(n399), .Q(n9228) );
  hi1s1 U10235 ( .DIN(n5471), .Q(n5368) );
  nnd2s1 U10236 ( .DIN1(n33), .DIN2(n9229), .Q(n9227) );
  nnd3s1 U10237 ( .DIN1(n9230), .DIN2(n9231), .DIN3(n5469), .Q(n9229) );
  nnd2s1 U10238 ( .DIN1(n9233), .DIN2(n9234), .Q(n5471) );
  nnd4s1 U10239 ( .DIN1(n9457), .DIN2(n9233), .DIN3(n9235), .DIN4(n9456), 
        .Q(n9232) );
  nor2s1 U10240 ( .DIN1(n9416), .DIN2(n9454), .Q(n9235) );
  nnd2s1 U10241 ( .DIN1(n8616), .DIN2(n754), .Q(n9231) );
  and2s1 U10242 ( .DIN1(n7138), .DIN2(n629), .Q(n8616) );
  hi1s1 U10243 ( .DIN(n5342), .Q(n7138) );
  nnd2s1 U10244 ( .DIN1(n9236), .DIN2(n7107), .Q(n5342) );
  hi1s1 U10245 ( .DIN(n9219), .Q(n7107) );
  nnd2s1 U10246 ( .DIN1(n9237), .DIN2(n9238), .Q(n9219) );
  nnd2s1 U10247 ( .DIN1(n775), .DIN2(n399), .Q(n9230) );
  nnd2s1 U10248 ( .DIN1(n7398), .DIN2(n9239), .Q(n9226) );
  nnd2s1 U10249 ( .DIN1(n9240), .DIN2(n5337), .Q(n9239) );
  nnd2s1 U10250 ( .DIN1(n9241), .DIN2(n9242), .Q(n9240) );
  or2s1 U10251 ( .DIN1(n7086), .DIN2(n204), .Q(n9242) );
  and2s1 U10252 ( .DIN1(n769), .DIN2(n9243), .Q(n7398) );
  nnd2s1 U10253 ( .DIN1(n716), .DIN2(n401), .Q(n9243) );
  nor2s1 U10254 ( .DIN1(n9218), .DIN2(n9244), .Q(n5336) );
  nnd3s1 U10255 ( .DIN1(n19), .DIN2(n2), .DIN3(n9238), .Q(n9218) );
  nnd2s1 U10256 ( .DIN1(n9245), .DIN2(n9246), .Q(n9224) );
  nnd3s1 U10257 ( .DIN1(n5375), .DIN2(n5381), .DIN3(n5372), .Q(n9245) );
  nnd3s1 U10258 ( .DIN1(n9458), .DIN2(n2), .DIN3(n9234), .Q(n5372) );
  and3s1 U10259 ( .DIN1(n9456), .DIN2(n17), .DIN3(n9217), .Q(n9234) );
  or3s1 U10260 ( .DIN1(n17), .DIN2(n137), .DIN3(n9215), .Q(n5381) );
  nnd2s1 U10261 ( .DIN1(n9217), .DIN2(n9247), .Q(n9215) );
  or2s1 U10262 ( .DIN1(n9233), .DIN2(n9237), .Q(n9247) );
  nnd4s1 U10263 ( .DIN1(n9457), .DIN2(n9217), .DIN3(n9456), .DIN4(n2), 
        .Q(n5375) );
  nnd4s1 U10264 ( .DIN1(n9217), .DIN2(n137), .DIN3(n9248), .DIN4(n9249), 
        .Q(n9223) );
  nnd3s1 U10265 ( .DIN1(n9250), .DIN2(n9251), .DIN3(n17), .Q(n9249) );
  nnd2s1 U10266 ( .DIN1(n9252), .DIN2(n9233), .Q(n9251) );
  nnd2s1 U10267 ( .DIN1(n9253), .DIN2(n9237), .Q(n9250) );
  nnd4s1 U10268 ( .DIN1(n9254), .DIN2(n9255), .DIN3(n9256), .DIN4(n9457), 
        .Q(n9248) );
  nnd3s1 U10269 ( .DIN1(n9257), .DIN2(n9258), .DIN3(n2), .Q(n9256) );
  nnd2s1 U10270 ( .DIN1(n9253), .DIN2(n19), .Q(n9258) );
  and2s1 U10271 ( .DIN1(n9259), .DIN2(n9260), .Q(n9253) );
  nnd2s1 U10272 ( .DIN1(n9261), .DIN2(n9262), .Q(n9260) );
  nnd2s1 U10273 ( .DIN1(n9263), .DIN2(n5390), .Q(n9261) );
  nnd3s1 U10274 ( .DIN1(n9264), .DIN2(n5466), .DIN3(n5454), .Q(n9263) );
  nnd3s1 U10275 ( .DIN1(n5621), .DIN2(n5463), .DIN3(n9265), .Q(n9264) );
  nnd3s1 U10276 ( .DIN1(n9266), .DIN2(n5768), .DIN3(n5756), .Q(n9265) );
  nnd3s1 U10277 ( .DIN1(n5853), .DIN2(n5765), .DIN3(n9267), .Q(n9266) );
  nnd3s1 U10278 ( .DIN1(n9268), .DIN2(n5992), .DIN3(n5980), .Q(n9267) );
  nnd3s1 U10279 ( .DIN1(n6075), .DIN2(n5989), .DIN3(n9269), .Q(n9268) );
  nnd3s1 U10280 ( .DIN1(n9270), .DIN2(n6209), .DIN3(n6197), .Q(n9269) );
  nnd3s1 U10281 ( .DIN1(n6284), .DIN2(n6206), .DIN3(n9271), .Q(n9270) );
  nnd3s1 U10282 ( .DIN1(n9272), .DIN2(n6427), .DIN3(n6415), .Q(n9271) );
  nnd3s1 U10283 ( .DIN1(n6505), .DIN2(n6424), .DIN3(n9273), .Q(n9272) );
  nnd3s1 U10284 ( .DIN1(n9274), .DIN2(n6636), .DIN3(n6624), .Q(n9273) );
  nnd3s1 U10285 ( .DIN1(n6713), .DIN2(n6633), .DIN3(n9275), .Q(n9274) );
  nnd3s1 U10286 ( .DIN1(n9276), .DIN2(n6856), .DIN3(n6844), .Q(n9275) );
  nnd3s1 U10287 ( .DIN1(n6938), .DIN2(n6853), .DIN3(n9277), .Q(n9276) );
  nnd3s1 U10288 ( .DIN1(n9278), .DIN2(n7085), .DIN3(n7073), .Q(n9277) );
  nnd3s1 U10289 ( .DIN1(n7134), .DIN2(n7082), .DIN3(n9279), .Q(n9278) );
  nnd3s1 U10290 ( .DIN1(n9280), .DIN2(n7262), .DIN3(n7250), .Q(n9279) );
  nnd3s1 U10291 ( .DIN1(n7383), .DIN2(n7259), .DIN3(n9281), .Q(n9280) );
  nnd3s1 U10292 ( .DIN1(n9282), .DIN2(n7510), .DIN3(n7498), .Q(n9281) );
  nnd3s1 U10293 ( .DIN1(n7632), .DIN2(n7507), .DIN3(n9283), .Q(n9282) );
  nnd3s1 U10294 ( .DIN1(n9284), .DIN2(n7752), .DIN3(n7740), .Q(n9283) );
  nnd3s1 U10295 ( .DIN1(n7862), .DIN2(n7749), .DIN3(n9285), .Q(n9284) );
  nnd3s1 U10296 ( .DIN1(n9286), .DIN2(n7987), .DIN3(n7975), .Q(n9285) );
  nnd3s1 U10297 ( .DIN1(n8098), .DIN2(n7984), .DIN3(n9287), .Q(n9286) );
  nnd3s1 U10298 ( .DIN1(n9288), .DIN2(n8224), .DIN3(n8212), .Q(n9287) );
  nnd3s1 U10299 ( .DIN1(n8357), .DIN2(n8221), .DIN3(n9289), .Q(n9288) );
  nnd3s1 U10300 ( .DIN1(n9290), .DIN2(n8495), .DIN3(n8483), .Q(n9289) );
  nnd3s1 U10301 ( .DIN1(n8612), .DIN2(n8492), .DIN3(n9291), .Q(n9290) );
  nnd4s1 U10302 ( .DIN1(n8739), .DIN2(n9292), .DIN3(n9293), .DIN4(n211), 
        .Q(n9291) );
  or2s1 U10303 ( .DIN1(n7106), .DIN2(n432), .Q(n9293) );
  nor2s1 U10304 ( .DIN1(n5353), .DIN2(n331), .Q(n7106) );
  nnd2s1 U10305 ( .DIN1(n715), .DIN2(n331), .Q(n9292) );
  hi1s1 U10306 ( .DIN(n8736), .Q(n8739) );
  nnd2s1 U10307 ( .DIN1(n9252), .DIN2(n9458), .Q(n9257) );
  and2s1 U10308 ( .DIN1(n9262), .DIN2(n9294), .Q(n9252) );
  nnd2s1 U10309 ( .DIN1(n9295), .DIN2(n9259), .Q(n9294) );
  nnd2s1 U10310 ( .DIN1(n5387), .DIN2(n9296), .Q(n9295) );
  nnd3s1 U10311 ( .DIN1(n9297), .DIN2(n5463), .DIN3(n5454), .Q(n9296) );
  nnd3s1 U10312 ( .DIN1(n9298), .DIN2(n5466), .DIN3(n5623), .Q(n9297) );
  nnd3s1 U10313 ( .DIN1(n9299), .DIN2(n5765), .DIN3(n5756), .Q(n9298) );
  nnd3s1 U10314 ( .DIN1(n9300), .DIN2(n5768), .DIN3(n5855), .Q(n9299) );
  nnd3s1 U10315 ( .DIN1(n9301), .DIN2(n5989), .DIN3(n5980), .Q(n9300) );
  nnd3s1 U10316 ( .DIN1(n9302), .DIN2(n5992), .DIN3(n6077), .Q(n9301) );
  nnd3s1 U10317 ( .DIN1(n9303), .DIN2(n6206), .DIN3(n6197), .Q(n9302) );
  nnd3s1 U10318 ( .DIN1(n9304), .DIN2(n6209), .DIN3(n6286), .Q(n9303) );
  nnd3s1 U10319 ( .DIN1(n9305), .DIN2(n6424), .DIN3(n6415), .Q(n9304) );
  nnd3s1 U10320 ( .DIN1(n9306), .DIN2(n6427), .DIN3(n6507), .Q(n9305) );
  nnd3s1 U10321 ( .DIN1(n9307), .DIN2(n6633), .DIN3(n6624), .Q(n9306) );
  nnd3s1 U10322 ( .DIN1(n9308), .DIN2(n6636), .DIN3(n6715), .Q(n9307) );
  nnd3s1 U10323 ( .DIN1(n9309), .DIN2(n6853), .DIN3(n6844), .Q(n9308) );
  nnd3s1 U10324 ( .DIN1(n9310), .DIN2(n6856), .DIN3(n6940), .Q(n9309) );
  nnd3s1 U10325 ( .DIN1(n9311), .DIN2(n7082), .DIN3(n7073), .Q(n9310) );
  nnd3s1 U10326 ( .DIN1(n9312), .DIN2(n7085), .DIN3(n7136), .Q(n9311) );
  nnd3s1 U10327 ( .DIN1(n9313), .DIN2(n7259), .DIN3(n7250), .Q(n9312) );
  nnd3s1 U10328 ( .DIN1(n9314), .DIN2(n7262), .DIN3(n7385), .Q(n9313) );
  nnd3s1 U10329 ( .DIN1(n9315), .DIN2(n7507), .DIN3(n7498), .Q(n9314) );
  nnd3s1 U10330 ( .DIN1(n9316), .DIN2(n7510), .DIN3(n7634), .Q(n9315) );
  nnd3s1 U10331 ( .DIN1(n9317), .DIN2(n7749), .DIN3(n7740), .Q(n9316) );
  nnd3s1 U10332 ( .DIN1(n9318), .DIN2(n7752), .DIN3(n7864), .Q(n9317) );
  nnd3s1 U10333 ( .DIN1(n9319), .DIN2(n7984), .DIN3(n7975), .Q(n9318) );
  nnd3s1 U10334 ( .DIN1(n9320), .DIN2(n7987), .DIN3(n8100), .Q(n9319) );
  nnd3s1 U10335 ( .DIN1(n9321), .DIN2(n8221), .DIN3(n8212), .Q(n9320) );
  nnd3s1 U10336 ( .DIN1(n9322), .DIN2(n8224), .DIN3(n8359), .Q(n9321) );
  nnd3s1 U10337 ( .DIN1(n9323), .DIN2(n8492), .DIN3(n8483), .Q(n9322) );
  nnd3s1 U10338 ( .DIN1(n9324), .DIN2(n8495), .DIN3(n8614), .Q(n9323) );
  hi1s1 U10339 ( .DIN(n8743), .Q(n9324) );
  nor2s1 U10340 ( .DIN1(n8615), .DIN2(n8736), .Q(n8743) );
  nnd2s1 U10341 ( .DIN1(n9325), .DIN2(n9326), .Q(n8615) );
  nnd2s1 U10342 ( .DIN1(n9327), .DIN2(n714), .Q(n9326) );
  nnd2s1 U10343 ( .DIN1(n8878), .DIN2(n330), .Q(n9327) );
  nnd2s1 U10344 ( .DIN1(n432), .DIN2(n8873), .Q(n9325) );
  nnd2s1 U10345 ( .DIN1(n9233), .DIN2(n9328), .Q(n9255) );
  nor2s1 U10346 ( .DIN1(n2), .DIN2(n9458), .Q(n9233) );
  nnd2s1 U10347 ( .DIN1(n9329), .DIN2(n9237), .Q(n9254) );
  nor2s1 U10348 ( .DIN1(n2), .DIN2(n19), .Q(n9237) );
  hi1s1 U10349 ( .DIN(n9328), .Q(n9329) );
  nnd2s1 U10350 ( .DIN1(n9330), .DIN2(n9331), .Q(n9328) );
  nor4s1 U10351 ( .DIN1(n9332), .DIN2(n9333), .DIN3(n9334), .DIN4(n9335), 
        .Q(n9331) );
  nnd4s1 U10352 ( .DIN1(n7073), .DIN2(n6929), .DIN3(n6844), .DIN4(n6704), 
        .Q(n9335) );
  hi1s1 U10353 ( .DIN(n6701), .Q(n6704) );
  nnd2s1 U10354 ( .DIN1(n6633), .DIN2(n6636), .Q(n6701) );
  nnd2s1 U10355 ( .DIN1(reg_out_B[19]), .DIN2(n37), .Q(n6636) );
  nnd2s1 U10356 ( .DIN1(n414), .DIN2(n144), .Q(n6633) );
  hi1s1 U10357 ( .DIN(n6841), .Q(n6844) );
  nnd2s1 U10358 ( .DIN1(n6713), .DIN2(n6715), .Q(n6841) );
  nnd2s1 U10359 ( .DIN1(reg_out_B[18]), .DIN2(n70), .Q(n6715) );
  nnd2s1 U10360 ( .DIN1(n415), .DIN2(n45), .Q(n6713) );
  hi1s1 U10361 ( .DIN(n6926), .Q(n6929) );
  nnd2s1 U10362 ( .DIN1(n6853), .DIN2(n6856), .Q(n6926) );
  nnd2s1 U10363 ( .DIN1(reg_out_B[17]), .DIN2(n82), .Q(n6856) );
  nnd2s1 U10364 ( .DIN1(n416), .DIN2(n135), .Q(n6853) );
  hi1s1 U10365 ( .DIN(n7070), .Q(n7073) );
  nnd2s1 U10366 ( .DIN1(n6938), .DIN2(n6940), .Q(n7070) );
  nnd2s1 U10367 ( .DIN1(reg_out_B[16]), .DIN2(n71), .Q(n6940) );
  nnd2s1 U10368 ( .DIN1(n417), .DIN2(n21), .Q(n6938) );
  nnd4s1 U10369 ( .DIN1(n6624), .DIN2(n6496), .DIN3(n6415), .DIN4(n6275), 
        .Q(n9334) );
  hi1s1 U10370 ( .DIN(n6272), .Q(n6275) );
  nnd2s1 U10371 ( .DIN1(n6206), .DIN2(n6209), .Q(n6272) );
  nnd2s1 U10372 ( .DIN1(reg_out_B[23]), .DIN2(n68), .Q(n6209) );
  nnd2s1 U10373 ( .DIN1(n410), .DIN2(n53), .Q(n6206) );
  hi1s1 U10374 ( .DIN(n6412), .Q(n6415) );
  nnd2s1 U10375 ( .DIN1(n6284), .DIN2(n6286), .Q(n6412) );
  nnd2s1 U10376 ( .DIN1(reg_out_B[22]), .DIN2(n67), .Q(n6286) );
  nnd2s1 U10377 ( .DIN1(n411), .DIN2(n3), .Q(n6284) );
  hi1s1 U10378 ( .DIN(n6493), .Q(n6496) );
  nnd2s1 U10379 ( .DIN1(n6424), .DIN2(n6427), .Q(n6493) );
  nnd2s1 U10380 ( .DIN1(reg_out_B[21]), .DIN2(n78), .Q(n6427) );
  nnd2s1 U10381 ( .DIN1(n412), .DIN2(n23), .Q(n6424) );
  hi1s1 U10382 ( .DIN(n6621), .Q(n6624) );
  nnd2s1 U10383 ( .DIN1(n6505), .DIN2(n6507), .Q(n6621) );
  nnd2s1 U10384 ( .DIN1(reg_out_B[20]), .DIN2(n69), .Q(n6507) );
  nnd2s1 U10385 ( .DIN1(n413), .DIN2(n52), .Q(n6505) );
  nnd4s1 U10386 ( .DIN1(n6197), .DIN2(n6066), .DIN3(n5980), .DIN4(n5844), 
        .Q(n9333) );
  hi1s1 U10387 ( .DIN(n5841), .Q(n5844) );
  nnd2s1 U10388 ( .DIN1(n5765), .DIN2(n5768), .Q(n5841) );
  nnd2s1 U10389 ( .DIN1(reg_out_B[27]), .DIN2(n38), .Q(n5768) );
  nnd2s1 U10390 ( .DIN1(n407), .DIN2(n134), .Q(n5765) );
  hi1s1 U10391 ( .DIN(n5977), .Q(n5980) );
  nnd2s1 U10392 ( .DIN1(n5853), .DIN2(n5855), .Q(n5977) );
  nnd2s1 U10393 ( .DIN1(reg_out_B[26]), .DIN2(n336), .Q(n5855) );
  nnd2s1 U10394 ( .DIN1(n435), .DIN2(n20), .Q(n5853) );
  hi1s1 U10395 ( .DIN(n6063), .Q(n6066) );
  nnd2s1 U10396 ( .DIN1(n5989), .DIN2(n5992), .Q(n6063) );
  nnd2s1 U10397 ( .DIN1(reg_out_B[25]), .DIN2(n83), .Q(n5992) );
  nnd2s1 U10398 ( .DIN1(n408), .DIN2(n25), .Q(n5989) );
  hi1s1 U10399 ( .DIN(n6194), .Q(n6197) );
  nnd2s1 U10400 ( .DIN1(n6075), .DIN2(n6077), .Q(n6194) );
  nnd2s1 U10401 ( .DIN1(reg_out_B[24]), .DIN2(n30), .Q(n6077) );
  nnd2s1 U10402 ( .DIN1(n409), .DIN2(n145), .Q(n6075) );
  nnd4s1 U10403 ( .DIN1(n5756), .DIN2(n5612), .DIN3(n5454), .DIN4(n5377), 
        .Q(n9332) );
  hi1s1 U10404 ( .DIN(n5370), .Q(n5377) );
  nnd2s1 U10405 ( .DIN1(n9259), .DIN2(n9262), .Q(n5370) );
  nnd2s1 U10406 ( .DIN1(n734), .DIN2(n133), .Q(n9262) );
  nnd2s1 U10407 ( .DIN1(reg_out_B[31]), .DIN2(n62), .Q(n9259) );
  hi1s1 U10408 ( .DIN(n5450), .Q(n5454) );
  nnd2s1 U10409 ( .DIN1(n5387), .DIN2(n5390), .Q(n5450) );
  nnd2s1 U10410 ( .DIN1(n718), .DIN2(n18), .Q(n5390) );
  nnd2s1 U10411 ( .DIN1(reg_out_B[30]), .DIN2(n717), .Q(n5387) );
  hi1s1 U10412 ( .DIN(n5609), .Q(n5612) );
  nnd2s1 U10413 ( .DIN1(n5463), .DIN2(n5466), .Q(n5609) );
  nnd2s1 U10414 ( .DIN1(reg_out_B[29]), .DIN2(n79), .Q(n5466) );
  nnd2s1 U10415 ( .DIN1(n406), .DIN2(n43), .Q(n5463) );
  hi1s1 U10416 ( .DIN(n5753), .Q(n5756) );
  nnd2s1 U10417 ( .DIN1(n5621), .DIN2(n5623), .Q(n5753) );
  nnd2s1 U10418 ( .DIN1(reg_out_B[28]), .DIN2(n335), .Q(n5623) );
  nnd2s1 U10419 ( .DIN1(n12), .DIN2(n44), .Q(n5621) );
  nor4s1 U10420 ( .DIN1(n9336), .DIN2(n9337), .DIN3(n9338), .DIN4(n9339), 
        .Q(n9330) );
  or4s1 U10421 ( .DIN1(n8869), .DIN2(n9246), .DIN3(n8736), .DIN4(n8600), 
        .Q(n9339) );
  nnd2s1 U10422 ( .DIN1(n8492), .DIN2(n8495), .Q(n8600) );
  nnd2s1 U10423 ( .DIN1(n438), .DIN2(n77), .Q(n8495) );
  nnd2s1 U10424 ( .DIN1(n431), .DIN2(n337), .Q(n8492) );
  nnd2s1 U10425 ( .DIN1(n8612), .DIN2(n8614), .Q(n8736) );
  nnd2s1 U10426 ( .DIN1(n742), .DIN2(n80), .Q(n8614) );
  nnd2s1 U10427 ( .DIN1(n426), .DIN2(n5490), .Q(n8612) );
  nnd2s1 U10428 ( .DIN1(n8873), .DIN2(n9340), .Q(n9246) );
  nnd2s1 U10429 ( .DIN1(n430), .DIN2(n1), .Q(n9340) );
  hi1s1 U10430 ( .DIN(n8878), .Q(n8873) );
  nor2s1 U10431 ( .DIN1(n1), .DIN2(n33), .Q(n8878) );
  xnr2s1 U10432 ( .DIN1(reg_out_B[1]), .DIN2(n330), .Q(n8869) );
  nnd4s1 U10433 ( .DIN1(n8483), .DIN2(n8348), .DIN3(n8212), .DIN4(n8089), 
        .Q(n9338) );
  hi1s1 U10434 ( .DIN(n8086), .Q(n8089) );
  nnd2s1 U10435 ( .DIN1(n7984), .DIN2(n7987), .Q(n8086) );
  nnd2s1 U10436 ( .DIN1(reg_out_B[7]), .DIN2(n63), .Q(n7987) );
  nnd2s1 U10437 ( .DIN1(n429), .DIN2(n51), .Q(n7984) );
  hi1s1 U10438 ( .DIN(n8209), .Q(n8212) );
  nnd2s1 U10439 ( .DIN1(n8098), .DIN2(n8100), .Q(n8209) );
  nnd2s1 U10440 ( .DIN1(reg_out_B[6]), .DIN2(n333), .Q(n8100) );
  nnd2s1 U10441 ( .DIN1(n34), .DIN2(n143), .Q(n8098) );
  hi1s1 U10442 ( .DIN(n8345), .Q(n8348) );
  nnd2s1 U10443 ( .DIN1(n8221), .DIN2(n8224), .Q(n8345) );
  nnd2s1 U10444 ( .DIN1(n716), .DIN2(n81), .Q(n8224) );
  nnd2s1 U10445 ( .DIN1(n428), .DIN2(n5337), .Q(n8221) );
  hi1s1 U10446 ( .DIN(n8480), .Q(n8483) );
  nnd2s1 U10447 ( .DIN1(n8357), .DIN2(n8359), .Q(n8480) );
  nnd2s1 U10448 ( .DIN1(n753), .DIN2(n334), .Q(n8359) );
  nnd2s1 U10449 ( .DIN1(n10), .DIN2(n808), .Q(n8357) );
  nnd4s1 U10450 ( .DIN1(n7975), .DIN2(n7853), .DIN3(n7740), .DIN4(n7623), 
        .Q(n9337) );
  hi1s1 U10451 ( .DIN(n7620), .Q(n7623) );
  nnd2s1 U10452 ( .DIN1(n7507), .DIN2(n7510), .Q(n7620) );
  nnd2s1 U10453 ( .DIN1(reg_out_B[11]), .DIN2(n84), .Q(n7510) );
  nnd2s1 U10454 ( .DIN1(n422), .DIN2(n136), .Q(n7507) );
  hi1s1 U10455 ( .DIN(n7737), .Q(n7740) );
  nnd2s1 U10456 ( .DIN1(n7632), .DIN2(n7634), .Q(n7737) );
  nnd2s1 U10457 ( .DIN1(reg_out_B[10]), .DIN2(n65), .Q(n7634) );
  nnd2s1 U10458 ( .DIN1(n423), .DIN2(n22), .Q(n7632) );
  hi1s1 U10459 ( .DIN(n7850), .Q(n7853) );
  nnd2s1 U10460 ( .DIN1(n7749), .DIN2(n7752), .Q(n7850) );
  nnd2s1 U10461 ( .DIN1(reg_out_B[9]), .DIN2(n66), .Q(n7752) );
  nnd2s1 U10462 ( .DIN1(n424), .DIN2(n4), .Q(n7749) );
  hi1s1 U10463 ( .DIN(n7972), .Q(n7975) );
  nnd2s1 U10464 ( .DIN1(n7862), .DIN2(n7864), .Q(n7972) );
  nnd2s1 U10465 ( .DIN1(reg_out_B[8]), .DIN2(n332), .Q(n7864) );
  nnd2s1 U10466 ( .DIN1(n425), .DIN2(n24), .Q(n7862) );
  nnd4s1 U10467 ( .DIN1(n7498), .DIN2(n7374), .DIN3(n7250), .DIN4(n7125), 
        .Q(n9336) );
  hi1s1 U10468 ( .DIN(n7122), .Q(n7125) );
  nnd2s1 U10469 ( .DIN1(n7082), .DIN2(n7085), .Q(n7122) );
  nnd2s1 U10470 ( .DIN1(reg_out_B[15]), .DIN2(n85), .Q(n7085) );
  nnd2s1 U10471 ( .DIN1(n418), .DIN2(n26), .Q(n7082) );
  hi1s1 U10472 ( .DIN(n7247), .Q(n7250) );
  nnd2s1 U10473 ( .DIN1(n7134), .DIN2(n7136), .Q(n7247) );
  nnd2s1 U10474 ( .DIN1(reg_out_B[14]), .DIN2(n31), .Q(n7136) );
  nnd2s1 U10475 ( .DIN1(n419), .DIN2(n146), .Q(n7134) );
  hi1s1 U10476 ( .DIN(n7371), .Q(n7374) );
  nnd2s1 U10477 ( .DIN1(n7259), .DIN2(n7262), .Q(n7371) );
  nnd2s1 U10478 ( .DIN1(reg_out_B[13]), .DIN2(n86), .Q(n7262) );
  nnd2s1 U10479 ( .DIN1(n420), .DIN2(n54), .Q(n7259) );
  hi1s1 U10480 ( .DIN(n7495), .Q(n7498) );
  nnd2s1 U10481 ( .DIN1(n7383), .DIN2(n7385), .Q(n7495) );
  nnd2s1 U10482 ( .DIN1(reg_out_B[12]), .DIN2(n64), .Q(n7385) );
  nnd2s1 U10483 ( .DIN1(n421), .DIN2(n46), .Q(n7383) );
  and2s1 U10484 ( .DIN1(n9416), .DIN2(n377), .Q(n9217) );
  nnd2s1 U10485 ( .DIN1(n9341), .DIN2(n9241), .Q(n9222) );
  nnd2s1 U10486 ( .DIN1(n9342), .DIN2(n204), .Q(n9241) );
  nnd4s1 U10487 ( .DIN1(n9343), .DIN2(n9344), .DIN3(n9345), .DIN4(n9346), 
        .Q(n9342) );
  nnd2s1 U10488 ( .DIN1(n628), .DIN2(n9347), .Q(n9346) );
  nnd4s1 U10489 ( .DIN1(n9348), .DIN2(n9349), .DIN3(n9350), .DIN4(n9351), 
        .Q(n9347) );
  nnd2s1 U10490 ( .DIN1(n771), .DIN2(n80), .Q(n9351) );
  nnd2s1 U10491 ( .DIN1(n532), .DIN2(n77), .Q(n9350) );
  nnd2s1 U10492 ( .DIN1(n773), .DIN2(n330), .Q(n9349) );
  nnd2s1 U10493 ( .DIN1(n755), .DIN2(n331), .Q(n9348) );
  or2s1 U10494 ( .DIN1(n7526), .DIN2(n5359), .Q(n9345) );
  hi1s1 U10495 ( .DIN(n5876), .Q(n5359) );
  nnd4s1 U10496 ( .DIN1(n7514), .DIN2(n7269), .DIN3(n6876), .DIN4(n7104), 
        .Q(n7526) );
  nnd2s1 U10497 ( .DIN1(n772), .DIN2(n419), .Q(n7104) );
  nnd2s1 U10498 ( .DIN1(n531), .DIN2(n418), .Q(n6876) );
  nnd2s1 U10499 ( .DIN1(n774), .DIN2(n420), .Q(n7269) );
  nnd2s1 U10500 ( .DIN1(n754), .DIN2(n421), .Q(n7514) );
  or2s1 U10501 ( .DIN1(n8003), .DIN2(n208), .Q(n9344) );
  nnd4s1 U10502 ( .DIN1(n7991), .DIN2(n7757), .DIN3(n7270), .DIN4(n7517), 
        .Q(n8003) );
  nnd2s1 U10503 ( .DIN1(n771), .DIN2(n423), .Q(n7517) );
  nnd2s1 U10504 ( .DIN1(n532), .DIN2(n422), .Q(n7270) );
  nnd2s1 U10505 ( .DIN1(n773), .DIN2(n424), .Q(n7757) );
  nnd2s1 U10506 ( .DIN1(n755), .DIN2(n36), .Q(n7991) );
  or2s1 U10507 ( .DIN1(n8503), .DIN2(n140), .Q(n9343) );
  nnd4s1 U10508 ( .DIN1(n8509), .DIN2(n8228), .DIN3(n7758), .DIN4(n7994), 
        .Q(n8503) );
  nnd2s1 U10509 ( .DIN1(n772), .DIN2(n427), .Q(n7994) );
  nnd2s1 U10510 ( .DIN1(n531), .DIN2(n429), .Q(n7758) );
  nnd2s1 U10511 ( .DIN1(n774), .DIN2(n428), .Q(n8228) );
  nnd2s1 U10512 ( .DIN1(n754), .DIN2(n433), .Q(n8509) );
  nnd2s1 U10513 ( .DIN1(n5994), .DIN2(n9352), .Q(n9341) );
  nnd2s1 U10514 ( .DIN1(n386), .DIN2(n7086), .Q(n9352) );
  nnd4s1 U10515 ( .DIN1(n9353), .DIN2(n9354), .DIN3(n9355), .DIN4(n9356), 
        .Q(n7086) );
  nnd2s1 U10516 ( .DIN1(n5876), .DIN2(n7539), .Q(n9356) );
  nnd4s1 U10517 ( .DIN1(n5784), .DIN2(n5491), .DIN3(n9357), .DIN4(n9358), 
        .Q(n7539) );
  nnd2s1 U10518 ( .DIN1(n718), .DIN2(n772), .Q(n9358) );
  nnd2s1 U10519 ( .DIN1(n532), .DIN2(n734), .Q(n9357) );
  nnd2s1 U10520 ( .DIN1(n773), .DIN2(n406), .Q(n5491) );
  nnd2s1 U10521 ( .DIN1(n755), .DIN2(n434), .Q(n5784) );
  nor2s1 U10522 ( .DIN1(n337), .DIN2(n5490), .Q(n5876) );
  nnd2s1 U10523 ( .DIN1(n546), .DIN2(n7536), .Q(n9355) );
  nnd4s1 U10524 ( .DIN1(n6227), .DIN2(n6012), .DIN3(n5492), .DIN4(n5787), 
        .Q(n7536) );
  nnd2s1 U10525 ( .DIN1(n771), .DIN2(n6), .Q(n5787) );
  nnd2s1 U10526 ( .DIN1(n531), .DIN2(n407), .Q(n5492) );
  nnd2s1 U10527 ( .DIN1(n774), .DIN2(n408), .Q(n6012) );
  nnd2s1 U10528 ( .DIN1(n754), .DIN2(n409), .Q(n6227) );
  nnd2s1 U10529 ( .DIN1(n621), .DIN2(n7537), .Q(n9354) );
  nnd4s1 U10530 ( .DIN1(n6653), .DIN2(n6447), .DIN3(n9359), .DIN4(n9360), 
        .Q(n7537) );
  nnd2s1 U10531 ( .DIN1(n772), .DIN2(n411), .Q(n9360) );
  nnd2s1 U10532 ( .DIN1(n532), .DIN2(n410), .Q(n9359) );
  nnd2s1 U10533 ( .DIN1(n773), .DIN2(n412), .Q(n6447) );
  nnd2s1 U10534 ( .DIN1(n755), .DIN2(n413), .Q(n6653) );
  nnd2s1 U10535 ( .DIN1(n628), .DIN2(n7535), .Q(n9353) );
  nnd4s1 U10536 ( .DIN1(n7101), .DIN2(n6875), .DIN3(n6448), .DIN4(n6656), 
        .Q(n7535) );
  nnd2s1 U10537 ( .DIN1(n771), .DIN2(n415), .Q(n6656) );
  nnd2s1 U10538 ( .DIN1(n531), .DIN2(n414), .Q(n6448) );
  nnd2s1 U10539 ( .DIN1(n774), .DIN2(n416), .Q(n6875) );
  nnd2s1 U10540 ( .DIN1(n754), .DIN2(n417), .Q(n7101) );
  nnd2s1 U10541 ( .DIN1(n9361), .DIN2(n9236), .Q(n5994) );
  and2s1 U10542 ( .DIN1(n7108), .DIN2(n808), .Q(n9236) );
  nor2s1 U10543 ( .DIN1(n9244), .DIN2(reg_out_B[5]), .Q(n7108) );
  or4s1 U10544 ( .DIN1(n9362), .DIN2(n9363), .DIN3(n9364), .DIN4(n9365), 
        .Q(n9244) );
  nnd4s1 U10545 ( .DIN1(n134), .DIN2(n44), .DIN3(n20), .DIN4(n9366), .Q(n9365)
         );
  and3s1 U10546 ( .DIN1(n145), .DIN2(n25), .DIN3(n53), .Q(n9366) );
  nnd4s1 U10547 ( .DIN1(n18), .DIN2(n133), .DIN3(n43), .DIN4(n9367), .Q(n9364)
         );
  and4s1 U10548 ( .DIN1(n143), .DIN2(n51), .DIN3(n24), .DIN4(n4), .Q(n9367) );
  nnd4s1 U10549 ( .DIN1(n136), .DIN2(n46), .DIN3(n22), .DIN4(n9368), .Q(n9363)
         );
  and3s1 U10550 ( .DIN1(n146), .DIN2(n26), .DIN3(n54), .Q(n9368) );
  nnd4s1 U10551 ( .DIN1(n135), .DIN2(n45), .DIN3(n21), .DIN4(n9369), .Q(n9362)
         );
  and4s1 U10552 ( .DIN1(n144), .DIN2(n52), .DIN3(n23), .DIN4(n3), .Q(n9369) );
  hi1s1 U10553 ( .DIN(n9220), .Q(n9361) );
  nnd3s1 U10554 ( .DIN1(n9458), .DIN2(n2), .DIN3(n9238), .Q(n9220) );
  and4s1 U10555 ( .DIN1(n9416), .DIN2(n9454), .DIN3(n9456), .DIN4(n17), 
        .Q(n9238) );
  hi1s1 U10556 ( .DIN(n8728), .Q(n5324) );
  nnd4s1 U10557 ( .DIN1(n9370), .DIN2(n9022), .DIN3(n39), .DIN4(n117), 
        .Q(n8728) );
  nnd3s1 U10558 ( .DIN1(n9371), .DIN2(n9372), .DIN3(n9373), .Q(\EXinst/n1423 )
         );
  nnd3s1 U10559 ( .DIN1(n9370), .DIN2(IR_opcode_field[5]), .DIN3(n9053), 
        .Q(n9373) );
  and3s1 U10560 ( .DIN1(n760), .DIN2(n101), .DIN3(n550), .Q(n9370) );
  nnd2s1 U10561 ( .DIN1(word), .DIN2(n527), .Q(n9372) );
  nnd2s1 U10562 ( .DIN1(n9374), .DIN2(n550), .Q(n9371) );
  nnd2s1 U10563 ( .DIN1(n9375), .DIN2(n9376), .Q(\EXinst/n1387 ) );
  nnd2s1 U10564 ( .DIN1(n528), .DIN2(byte), .Q(n9376) );
  nnd3s1 U10565 ( .DIN1(n9022), .DIN2(n9035), .DIN3(n9453), .Q(n9375) );
  nnd2s1 U10566 ( .DIN1(n9377), .DIN2(n9378), .Q(n9035) );
  nnd3s1 U10567 ( .DIN1(n760), .DIN2(n101), .DIN3(IR_opcode_field[5]), 
        .Q(n9378) );
  nor2s1 U10568 ( .DIN1(n9415), .DIN2(n48), .Q(\EXinst/N1341 ) );
  nor2s1 U10569 ( .DIN1(n9414), .DIN2(n48), .Q(\EXinst/N1340 ) );
  and4s1 U10570 ( .DIN1(n9037), .DIN2(n551), .DIN3(n40), .DIN4(n760), 
        .Q(\EXinst/N1339 ) );
  nor2s1 U10571 ( .DIN1(n9413), .DIN2(n48), .Q(\EXinst/N1338 ) );
  and2s1 U10572 ( .DIN1(n551), .DIN2(reg_write), .Q(\EXinst/N1337 ) );
  nor2s1 U10573 ( .DIN1(n133), .DIN2(n9379), .Q(\EXinst/N1336 ) );
  nor2s1 U10574 ( .DIN1(n18), .DIN2(n9379), .Q(\EXinst/N1335 ) );
  nor2s1 U10575 ( .DIN1(n43), .DIN2(n9379), .Q(\EXinst/N1334 ) );
  nor2s1 U10576 ( .DIN1(n44), .DIN2(n9379), .Q(\EXinst/N1333 ) );
  nor2s1 U10577 ( .DIN1(n134), .DIN2(n9379), .Q(\EXinst/N1332 ) );
  nor2s1 U10578 ( .DIN1(n20), .DIN2(n9379), .Q(\EXinst/N1331 ) );
  nor2s1 U10579 ( .DIN1(n25), .DIN2(n9379), .Q(\EXinst/N1330 ) );
  nor2s1 U10580 ( .DIN1(n145), .DIN2(n9379), .Q(\EXinst/N1329 ) );
  nor2s1 U10581 ( .DIN1(n53), .DIN2(n9379), .Q(\EXinst/N1328 ) );
  nor2s1 U10582 ( .DIN1(n3), .DIN2(n9379), .Q(\EXinst/N1327 ) );
  nor2s1 U10583 ( .DIN1(n23), .DIN2(n9379), .Q(\EXinst/N1326 ) );
  nor2s1 U10584 ( .DIN1(n52), .DIN2(n9379), .Q(\EXinst/N1325 ) );
  nor2s1 U10585 ( .DIN1(n144), .DIN2(n9379), .Q(\EXinst/N1324 ) );
  nor2s1 U10586 ( .DIN1(n45), .DIN2(n9379), .Q(\EXinst/N1323 ) );
  nor2s1 U10587 ( .DIN1(n135), .DIN2(n9379), .Q(\EXinst/N1322 ) );
  nor2s1 U10588 ( .DIN1(n21), .DIN2(n9379), .Q(\EXinst/N1321 ) );
  nnd3s1 U10589 ( .DIN1(n9380), .DIN2(n9381), .DIN3(n9453), .Q(n9379) );
  nnd2s1 U10590 ( .DIN1(n9374), .DIN2(n11), .Q(n9380) );
  and3s1 U10591 ( .DIN1(n9037), .DIN2(IR_opcode_field[3]), .DIN3(n9053), 
        .Q(n9374) );
  nor2s1 U10592 ( .DIN1(n132), .DIN2(IR_opcode_field[1]), .Q(n9053) );
  nor2s1 U10593 ( .DIN1(n26), .DIN2(n9382), .Q(\EXinst/N1320 ) );
  nor2s1 U10594 ( .DIN1(n146), .DIN2(n9382), .Q(\EXinst/N1319 ) );
  nor2s1 U10595 ( .DIN1(n54), .DIN2(n9382), .Q(\EXinst/N1318 ) );
  nor2s1 U10596 ( .DIN1(n46), .DIN2(n9382), .Q(\EXinst/N1317 ) );
  nor2s1 U10597 ( .DIN1(n136), .DIN2(n9382), .Q(\EXinst/N1316 ) );
  nor2s1 U10598 ( .DIN1(n22), .DIN2(n9382), .Q(\EXinst/N1315 ) );
  nor2s1 U10599 ( .DIN1(n4), .DIN2(n9382), .Q(\EXinst/N1314 ) );
  nor2s1 U10600 ( .DIN1(n24), .DIN2(n9382), .Q(\EXinst/N1313 ) );
  nnd2s1 U10601 ( .DIN1(n551), .DIN2(n9381), .Q(n9382) );
  nnd4s1 U10602 ( .DIN1(n9037), .DIN2(n9022), .DIN3(IR_opcode_field[3]), 
        .DIN4(n11), .Q(n9381) );
  nor2s1 U10603 ( .DIN1(IR_opcode_field[0]), .DIN2(IR_opcode_field[1]), 
        .Q(n9022) );
  hi1s1 U10604 ( .DIN(n9377), .Q(n9037) );
  nnd3s1 U10605 ( .DIN1(n39), .DIN2(n101), .DIN3(IR_opcode_field[5]), 
        .Q(n9377) );
  nor2s1 U10606 ( .DIN1(n528), .DIN2(n51), .Q(\EXinst/N1312 ) );
  nor2s1 U10607 ( .DIN1(n48), .DIN2(n143), .Q(\EXinst/N1311 ) );
  nor2s1 U10608 ( .DIN1(n527), .DIN2(n5337), .Q(\EXinst/N1310 ) );
  hi1s1 U10609 ( .DIN(n716), .Q(n5337) );
  nor2s1 U10610 ( .DIN1(n527), .DIN2(n807), .Q(\EXinst/N1309 ) );
  nor2s1 U10611 ( .DIN1(n528), .DIN2(n337), .Q(\EXinst/N1308 ) );
  nor2s1 U10612 ( .DIN1(n528), .DIN2(n5490), .Q(\EXinst/N1307 ) );
  hi1s1 U10613 ( .DIN(n741), .Q(n5490) );
  nor2s1 U10614 ( .DIN1(n527), .DIN2(n714), .Q(\EXinst/N1306 ) );
  nor2s1 U10615 ( .DIN1(n527), .DIN2(n1), .Q(\EXinst/N1305 ) );
endmodule

