
module s35932 ( CK, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, 
        CRC_OUT_1_11, CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, 
        CRC_OUT_1_16, CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, 
        CRC_OUT_1_20, CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, 
        CRC_OUT_1_25, CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, 
        CRC_OUT_1_3, CRC_OUT_1_30, CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, 
        CRC_OUT_1_6, CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, 
        CRC_OUT_2_1, CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, 
        CRC_OUT_2_14, CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, 
        CRC_OUT_2_19, CRC_OUT_2_2, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, 
        CRC_OUT_2_23, CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, 
        CRC_OUT_2_28, CRC_OUT_2_29, CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, 
        CRC_OUT_2_4, CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, 
        CRC_OUT_2_9, CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, 
        CRC_OUT_3_12, CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, 
        CRC_OUT_3_17, CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, 
        CRC_OUT_3_21, CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, 
        CRC_OUT_3_26, CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, 
        CRC_OUT_3_30, CRC_OUT_3_31, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, 
        CRC_OUT_3_7, CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, 
        CRC_OUT_4_10, CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, 
        CRC_OUT_4_15, CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, 
        CRC_OUT_4_2, CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, 
        CRC_OUT_4_24, CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, 
        CRC_OUT_4_29, CRC_OUT_4_3, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, 
        CRC_OUT_4_5, CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, 
        CRC_OUT_5_0, CRC_OUT_5_1, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, 
        CRC_OUT_5_13, CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, 
        CRC_OUT_5_18, CRC_OUT_5_19, CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, 
        CRC_OUT_5_22, CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, 
        CRC_OUT_5_27, CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, 
        CRC_OUT_5_31, CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, 
        CRC_OUT_5_8, CRC_OUT_5_9, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, 
        CRC_OUT_6_11, CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, 
        CRC_OUT_6_16, CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, 
        CRC_OUT_6_20, CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, 
        CRC_OUT_6_25, CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, 
        CRC_OUT_6_3, CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, 
        CRC_OUT_6_6, CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, 
        CRC_OUT_7_1, CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, 
        CRC_OUT_7_14, CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, 
        CRC_OUT_7_19, CRC_OUT_7_2, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, 
        CRC_OUT_7_23, CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, 
        CRC_OUT_7_28, CRC_OUT_7_29, CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, 
        CRC_OUT_7_4, CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, 
        CRC_OUT_7_9, CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, 
        CRC_OUT_8_12, CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, 
        CRC_OUT_8_17, CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, 
        CRC_OUT_8_21, CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, 
        CRC_OUT_8_26, CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, 
        CRC_OUT_8_30, CRC_OUT_8_31, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, 
        CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, 
        CRC_OUT_9_10, CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, 
        CRC_OUT_9_15, CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, 
        CRC_OUT_9_2, CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, 
        CRC_OUT_9_24, CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, 
        CRC_OUT_9_29, CRC_OUT_9_3, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, 
        CRC_OUT_9_5, CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, 
        DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12, DATA_0_13, 
        DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18, DATA_0_19, 
        DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23, DATA_0_24, 
        DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29, DATA_0_3, 
        DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6, DATA_0_7, DATA_0_8, 
        DATA_0_9, DATA_9_0, DATA_9_1, DATA_9_10, DATA_9_11, DATA_9_12, 
        DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16, DATA_9_17, DATA_9_18, 
        DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21, DATA_9_22, DATA_9_23, 
        DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27, DATA_9_28, DATA_9_29, 
        DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4, DATA_9_5, DATA_9_6, DATA_9_7, 
        DATA_9_8, DATA_9_9, RESET, TM0, TM1 );
  input  CK, DATA_0_0, DATA_0_1, DATA_0_10, DATA_0_11, DATA_0_12,
         DATA_0_13, DATA_0_14, DATA_0_15, DATA_0_16, DATA_0_17, DATA_0_18,
         DATA_0_19, DATA_0_2, DATA_0_20, DATA_0_21, DATA_0_22, DATA_0_23,
         DATA_0_24, DATA_0_25, DATA_0_26, DATA_0_27, DATA_0_28, DATA_0_29,
         DATA_0_3, DATA_0_30, DATA_0_31, DATA_0_4, DATA_0_5, DATA_0_6,
         DATA_0_7, DATA_0_8, DATA_0_9, RESET, TM0, TM1;
  output CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12,
         CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17,
         CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_2, CRC_OUT_1_20, CRC_OUT_1_21,
         CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26,
         CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_3, CRC_OUT_1_30,
         CRC_OUT_1_31, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7,
         CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_10,
         CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15,
         CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_2,
         CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24,
         CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29,
         CRC_OUT_2_3, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_2_4, CRC_OUT_2_5,
         CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_3_0,
         CRC_OUT_3_1, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13,
         CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18,
         CRC_OUT_3_19, CRC_OUT_3_2, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22,
         CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27,
         CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_3, CRC_OUT_3_30, CRC_OUT_3_31,
         CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8,
         CRC_OUT_3_9, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_10, CRC_OUT_4_11,
         CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16,
         CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_2, CRC_OUT_4_20,
         CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25,
         CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_3,
         CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6,
         CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_5_0, CRC_OUT_5_1,
         CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14,
         CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19,
         CRC_OUT_5_2, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23,
         CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28,
         CRC_OUT_5_29, CRC_OUT_5_3, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_5_4,
         CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9,
         CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12,
         CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17,
         CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_2, CRC_OUT_6_20, CRC_OUT_6_21,
         CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26,
         CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_3, CRC_OUT_6_30,
         CRC_OUT_6_31, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7,
         CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_10,
         CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15,
         CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_2,
         CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24,
         CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29,
         CRC_OUT_7_3, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_7_4, CRC_OUT_7_5,
         CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_8_0,
         CRC_OUT_8_1, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13,
         CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18,
         CRC_OUT_8_19, CRC_OUT_8_2, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22,
         CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27,
         CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_3, CRC_OUT_8_30, CRC_OUT_8_31,
         CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8,
         CRC_OUT_8_9, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_10, CRC_OUT_9_11,
         CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16,
         CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_2, CRC_OUT_9_20,
         CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25,
         CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_3,
         CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6,
         CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, DATA_9_0, DATA_9_1, DATA_9_10,
         DATA_9_11, DATA_9_12, DATA_9_13, DATA_9_14, DATA_9_15, DATA_9_16,
         DATA_9_17, DATA_9_18, DATA_9_19, DATA_9_2, DATA_9_20, DATA_9_21,
         DATA_9_22, DATA_9_23, DATA_9_24, DATA_9_25, DATA_9_26, DATA_9_27,
         DATA_9_28, DATA_9_29, DATA_9_3, DATA_9_30, DATA_9_31, DATA_9_4,
         DATA_9_5, DATA_9_6, DATA_9_7, DATA_9_8, DATA_9_9;
  wire   WX485, WX484, WX487, WX486, WX489, WX488, WX491, WX490, WX493, WX492,
         WX495, WX494, WX497, WX496, WX499, WX498, WX501, WX500, WX503, WX502,
         WX505, WX504, WX507, WX506, WX509, WX508, WX511, WX510, WX513, WX512,
         WX515, WX514, WX517, WX516, WX519, WX518, WX521, WX520, WX523, WX522,
         WX525, WX524, WX527, WX526, WX529, WX528, WX531, WX530, WX533, WX532,
         WX535, WX534, WX537, WX536, WX539, WX538, WX541, WX540, WX543, WX542,
         WX545, WX544, WX547, WX546, WX645, WX644, WX647, WX646, WX649, WX648,
         WX651, WX650, WX653, WX652, WX655, WX654, WX657, WX656, WX659, WX658,
         WX661, WX660, WX663, WX662, WX665, WX664, WX667, WX666, WX669, WX668,
         WX671, WX670, WX673, WX672, WX675, WX674, WX677, WX676, WX679, WX678,
         WX681, WX680, WX683, WX682, WX685, WX684, WX687, WX686, WX689, WX688,
         WX691, WX690, WX693, WX692, WX695, WX694, WX697, WX696, WX699, WX698,
         WX701, WX700, WX703, WX702, WX705, WX704, WX707, WX706, WX709, WX708,
         WX711, WX710, WX713, WX712, WX715, WX714, WX717, WX716, WX719, WX718,
         WX721, WX720, WX723, WX722, WX725, WX724, WX727, WX726, WX729, WX728,
         WX731, WX730, WX733, WX732, WX735, WX734, WX737, WX736, WX739, WX738,
         WX741, WX740, WX743, WX742, WX745, WX744, WX747, WX746, WX749, WX748,
         WX751, WX750, WX753, WX752, WX755, WX754, WX757, WX756, WX759, WX758,
         WX761, WX760, WX763, WX762, WX765, WX764, WX767, WX766, WX769, WX768,
         WX771, WX770, WX773, WX772, WX775, WX774, WX777, WX776, WX779, WX778,
         WX781, WX780, WX783, WX782, WX785, WX784, WX787, WX786, WX789, WX788,
         WX791, WX790, WX793, WX792, WX795, WX794, WX797, WX796, WX799, WX798,
         WX801, WX800, WX803, WX802, WX805, WX804, WX807, WX806, WX809, WX808,
         WX811, WX810, WX813, WX812, WX815, WX814, WX817, WX816, WX819, WX818,
         WX821, WX820, WX823, WX822, WX825, WX824, WX827, WX826, WX829, WX828,
         WX831, WX830, WX833, WX832, WX835, WX834, WX837, WX836, WX839, WX838,
         WX841, WX840, WX843, WX842, WX845, WX844, WX847, WX846, WX849, WX848,
         WX851, WX850, WX853, WX852, WX855, WX854, WX857, WX856, WX859, WX858,
         WX861, WX860, WX863, WX862, WX865, WX864, WX867, WX866, WX869, WX868,
         WX871, WX870, WX873, WX872, WX875, WX874, WX877, WX876, WX879, WX878,
         WX881, WX880, WX883, WX882, WX885, WX884, WX887, WX886, WX889, WX888,
         WX891, WX890, WX893, WX892, WX895, WX894, WX897, WX896, WX899, WX898,
         WX1264, WX1266, WX1268, WX1270, WX1272, WX1274, WX1276, WX1278,
         WX1280, WX1282, WX1284, WX1286, WX1288, WX1290, WX1292, WX1294,
         WX1296, WX1298, WX1300, WX1302, WX1304, WX1306, WX1308, WX1310,
         WX1312, WX1314, WX1316, WX1318, WX1320, WX1322, WX1324, WX1326,
         WX1778, WX1777, WX1780, WX1779, WX1782, WX1781, WX1784, WX1783,
         WX1786, WX1785, WX1788, WX1787, WX1790, WX1789, WX1792, WX1791,
         WX1794, WX1793, WX1796, WX1795, WX1798, WX1797, WX1800, WX1799,
         WX1802, WX1801, WX1804, WX1803, WX1806, WX1805, WX1808, WX1807,
         WX1810, WX1809, WX1812, WX1811, WX1814, WX1813, WX1816, WX1815,
         WX1818, WX1817, WX1820, WX1819, WX1822, WX1821, WX1824, WX1823,
         WX1826, WX1825, WX1828, WX1827, WX1830, WX1829, WX1832, WX1831,
         WX1834, WX1833, WX1836, WX1835, WX1838, WX1837, WX1840, WX1839,
         WX1938, WX1937, WX1940, WX1939, WX1942, WX1941, WX1944, WX1943,
         WX1946, WX1945, WX1948, WX1947, WX1950, WX1949, WX1952, WX1951,
         WX1954, WX1953, WX1956, WX1955, WX1958, WX1957, WX1960, WX1959,
         WX1962, WX1961, WX1964, WX1963, WX1966, WX1965, WX1968, WX1967,
         WX1970, WX1969, WX1972, WX1971, WX1974, WX1973, WX1976, WX1975,
         WX1978, WX1977, WX1980, WX1979, WX1982, WX1981, WX1984, WX1983,
         WX1986, WX1985, WX1988, WX1987, WX1990, WX1989, WX1992, WX1991,
         WX1994, WX1993, WX1996, WX1995, WX1998, WX1997, WX2000, WX1999,
         WX2001, WX2003, WX2005, WX2007, WX2009, WX2011, WX2013, WX2015,
         WX2017, WX2019, WX2021, WX2023, WX2025, WX2027, WX2029, WX2031,
         WX2033, WX2035, WX2037, WX2039, WX2041, WX2043, WX2045, WX2047,
         WX2049, WX2051, WX2053, WX2055, WX2057, WX2059, WX2061, WX2063,
         WX2066, WX2065, WX2068, WX2067, WX2070, WX2069, WX2072, WX2071,
         WX2074, WX2073, WX2076, WX2075, WX2078, WX2077, WX2080, WX2079,
         WX2082, WX2081, WX2084, WX2083, WX2086, WX2085, WX2088, WX2087,
         WX2090, WX2089, WX2092, WX2091, WX2094, WX2093, WX2096, WX2095,
         WX2098, WX2097, WX2100, WX2099, WX2102, WX2101, WX2104, WX2103,
         WX2106, WX2105, WX2108, WX2107, WX2110, WX2109, WX2112, WX2111,
         WX2114, WX2113, WX2116, WX2115, WX2118, WX2117, WX2120, WX2119,
         WX2122, WX2121, WX2124, WX2123, WX2126, WX2125, WX2128, WX2127,
         WX2130, WX2129, WX2132, WX2131, WX2134, WX2133, WX2136, WX2135,
         WX2138, WX2137, WX2140, WX2139, WX2142, WX2141, WX2144, WX2143,
         WX2146, WX2145, WX2148, WX2147, WX2150, WX2149, WX2152, WX2151,
         WX2154, WX2153, WX2156, WX2155, WX2158, WX2157, WX2160, WX2159,
         WX2162, WX2161, WX2164, WX2163, WX2166, WX2165, WX2168, WX2167,
         WX2170, WX2169, WX2172, WX2171, WX2174, WX2173, WX2176, WX2175,
         WX2178, WX2177, WX2180, WX2179, WX2182, WX2181, WX2184, WX2183,
         WX2186, WX2185, WX2188, WX2187, WX2190, WX2189, WX2192, WX2191,
         WX2557, WX2559, WX2561, WX2563, WX2565, WX2567, WX2569, WX2571,
         WX2573, WX2575, WX2577, WX2579, WX2581, WX2583, WX2585, WX2587,
         WX2589, WX2591, WX2593, WX2595, WX2597, WX2599, WX2601, WX2603,
         WX2605, WX2607, WX2609, WX2611, WX2613, WX2615, WX2617, WX2619,
         WX3071, WX3070, WX3073, WX3072, WX3075, WX3074, WX3077, WX3076,
         WX3079, WX3078, WX3081, WX3080, WX3083, WX3082, WX3085, WX3084,
         WX3087, WX3086, WX3089, WX3088, WX3091, WX3090, WX3093, WX3092,
         WX3095, WX3094, WX3097, WX3096, WX3099, WX3098, WX3101, WX3100,
         WX3103, WX3102, WX3105, WX3104, WX3107, WX3106, WX3109, WX3108,
         WX3111, WX3110, WX3113, WX3112, WX3115, WX3114, WX3117, WX3116,
         WX3119, WX3118, WX3121, WX3120, WX3123, WX3122, WX3125, WX3124,
         WX3127, WX3126, WX3129, WX3128, WX3131, WX3130, WX3133, WX3132,
         WX3231, WX3230, WX3233, WX3232, WX3235, WX3234, WX3237, WX3236,
         WX3239, WX3238, WX3241, WX3240, WX3243, WX3242, WX3245, WX3244,
         WX3247, WX3246, WX3249, WX3248, WX3251, WX3250, WX3253, WX3252,
         WX3255, WX3254, WX3257, WX3256, WX3259, WX3258, WX3261, WX3260,
         WX3262, WX3264, WX3266, WX3268, WX3270, WX3272, WX3274, WX3276,
         WX3278, WX3280, WX3282, WX3284, WX3286, WX3288, WX3290, WX3292,
         WX3294, WX3296, WX3298, WX3300, WX3302, WX3304, WX3306, WX3308,
         WX3310, WX3312, WX3314, WX3316, WX3318, WX3320, WX3322, WX3324,
         WX3327, WX3326, WX3329, WX3328, WX3331, WX3330, WX3333, WX3332,
         WX3335, WX3334, WX3337, WX3336, WX3339, WX3338, WX3341, WX3340,
         WX3343, WX3342, WX3345, WX3344, WX3347, WX3346, WX3349, WX3348,
         WX3351, WX3350, WX3353, WX3352, WX3355, WX3354, WX3357, WX3356,
         WX3359, WX3358, WX3361, WX3360, WX3363, WX3362, WX3365, WX3364,
         WX3367, WX3366, WX3369, WX3368, WX3371, WX3370, WX3373, WX3372,
         WX3375, WX3374, WX3377, WX3376, WX3379, WX3378, WX3381, WX3380,
         WX3383, WX3382, WX3385, WX3384, WX3387, WX3386, WX3389, WX3388,
         WX3391, WX3390, WX3393, WX3392, WX3395, WX3394, WX3397, WX3396,
         WX3399, WX3398, WX3401, WX3400, WX3403, WX3402, WX3405, WX3404,
         WX3407, WX3406, WX3409, WX3408, WX3411, WX3410, WX3413, WX3412,
         WX3415, WX3414, WX3417, WX3416, WX3419, WX3418, WX3421, WX3420,
         WX3423, WX3422, WX3425, WX3424, WX3427, WX3426, WX3429, WX3428,
         WX3431, WX3430, WX3433, WX3432, WX3435, WX3434, WX3437, WX3436,
         WX3439, WX3438, WX3441, WX3440, WX3443, WX3442, WX3445, WX3444,
         WX3447, WX3446, WX3449, WX3448, WX3451, WX3450, WX3453, WX3452,
         WX3455, WX3454, WX3457, WX3456, WX3459, WX3458, WX3461, WX3460,
         WX3463, WX3462, WX3465, WX3464, WX3467, WX3466, WX3469, WX3468,
         WX3471, WX3470, WX3473, WX3472, WX3475, WX3474, WX3477, WX3476,
         WX3479, WX3478, WX3481, WX3480, WX3483, WX3482, WX3485, WX3484,
         WX3850, WX3852, WX3854, WX3856, WX3858, WX3860, WX3862, WX3864,
         WX3866, WX3868, WX3870, WX3872, WX3874, WX3876, WX3878, WX3880,
         WX3882, WX3884, WX3886, WX3888, WX3890, WX3892, WX3894, WX3896,
         WX3898, WX3900, WX3902, WX3904, WX3906, WX3908, WX3910, WX3912,
         WX4364, WX4363, WX4366, WX4365, WX4368, WX4367, WX4370, WX4369,
         WX4372, WX4371, WX4374, WX4373, WX4376, WX4375, WX4378, WX4377,
         WX4380, WX4379, WX4382, WX4381, WX4384, WX4383, WX4386, WX4385,
         WX4388, WX4387, WX4390, WX4389, WX4392, WX4391, WX4394, WX4393,
         WX4396, WX4395, WX4398, WX4397, WX4400, WX4399, WX4402, WX4401,
         WX4404, WX4403, WX4406, WX4405, WX4408, WX4407, WX4410, WX4409,
         WX4412, WX4411, WX4414, WX4413, WX4416, WX4415, WX4418, WX4417,
         WX4420, WX4419, WX4422, WX4421, WX4424, WX4423, WX4426, WX4425,
         WX4524, WX4523, WX4526, WX4525, WX4528, WX4527, WX4530, WX4529,
         WX4532, WX4531, WX4534, WX4533, WX4536, WX4535, WX4538, WX4537,
         WX4540, WX4539, WX4542, WX4541, WX4544, WX4543, WX4546, WX4545,
         WX4548, WX4547, WX4550, WX4549, WX4552, WX4551, WX4554, WX4553,
         WX4555, WX4557, WX4559, WX4561, WX4563, WX4565, WX4567, WX4569,
         WX4571, WX4573, WX4575, WX4577, WX4579, WX4581, WX4583, WX4585,
         WX4587, WX4589, WX4591, WX4593, WX4595, WX4597, WX4599, WX4601,
         WX4603, WX4605, WX4607, WX4609, WX4611, WX4613, WX4615, WX4617,
         WX4620, WX4619, WX4622, WX4621, WX4624, WX4623, WX4626, WX4625,
         WX4628, WX4627, WX4630, WX4629, WX4632, WX4631, WX4634, WX4633,
         WX4636, WX4635, WX4638, WX4637, WX4640, WX4639, WX4642, WX4641,
         WX4644, WX4643, WX4646, WX4645, WX4648, WX4647, WX4650, WX4649,
         WX4652, WX4651, WX4654, WX4653, WX4656, WX4655, WX4658, WX4657,
         WX4660, WX4659, WX4662, WX4661, WX4664, WX4663, WX4666, WX4665,
         WX4668, WX4667, WX4670, WX4669, WX4672, WX4671, WX4674, WX4673,
         WX4676, WX4675, WX4678, WX4677, WX4680, WX4679, WX4682, WX4681,
         WX4684, WX4683, WX4686, WX4685, WX4688, WX4687, WX4690, WX4689,
         WX4692, WX4691, WX4694, WX4693, WX4696, WX4695, WX4698, WX4697,
         WX4700, WX4699, WX4702, WX4701, WX4704, WX4703, WX4706, WX4705,
         WX4708, WX4707, WX4710, WX4709, WX4712, WX4711, WX4714, WX4713,
         WX4716, WX4715, WX4718, WX4717, WX4720, WX4719, WX4722, WX4721,
         WX4724, WX4723, WX4726, WX4725, WX4728, WX4727, WX4730, WX4729,
         WX4732, WX4731, WX4734, WX4733, WX4736, WX4735, WX4738, WX4737,
         WX4740, WX4739, WX4742, WX4741, WX4744, WX4743, WX4746, WX4745,
         WX4748, WX4747, WX4750, WX4749, WX4752, WX4751, WX4754, WX4753,
         WX4756, WX4755, WX4758, WX4757, WX4760, WX4759, WX4762, WX4761,
         WX4764, WX4763, WX4766, WX4765, WX4768, WX4767, WX4770, WX4769,
         WX4772, WX4771, WX4774, WX4773, WX4776, WX4775, WX4778, WX4777,
         WX5143, WX5145, WX5147, WX5149, WX5151, WX5153, WX5155, WX5157,
         WX5159, WX5161, WX5163, WX5165, WX5167, WX5169, WX5171, WX5173,
         WX5175, WX5177, WX5179, WX5181, WX5183, WX5185, WX5187, WX5189,
         WX5191, WX5193, WX5195, WX5197, WX5199, WX5201, WX5203, WX5205,
         WX5657, WX5656, WX5659, WX5658, WX5661, WX5660, WX5663, WX5662,
         WX5665, WX5664, WX5667, WX5666, WX5669, WX5668, WX5671, WX5670,
         WX5673, WX5672, WX5675, WX5674, WX5677, WX5676, WX5679, WX5678,
         WX5681, WX5680, WX5683, WX5682, WX5685, WX5684, WX5687, WX5686,
         WX5689, WX5688, WX5691, WX5690, WX5693, WX5692, WX5695, WX5694,
         WX5697, WX5696, WX5699, WX5698, WX5701, WX5700, WX5703, WX5702,
         WX5705, WX5704, WX5707, WX5706, WX5709, WX5708, WX5711, WX5710,
         WX5713, WX5712, WX5715, WX5714, WX5717, WX5716, WX5719, WX5718,
         WX5817, WX5816, WX5819, WX5818, WX5821, WX5820, WX5823, WX5822,
         WX5825, WX5824, WX5827, WX5826, WX5829, WX5828, WX5831, WX5830,
         WX5833, WX5832, WX5835, WX5834, WX5837, WX5836, WX5839, WX5838,
         WX5841, WX5840, WX5843, WX5842, WX5845, WX5844, WX5847, WX5846,
         WX5848, WX5850, WX5852, WX5854, WX5856, WX5858, WX5860, WX5862,
         WX5864, WX5866, WX5868, WX5870, WX5872, WX5874, WX5876, WX5878,
         WX5880, WX5882, WX5884, WX5886, WX5888, WX5890, WX5892, WX5894,
         WX5896, WX5898, WX5900, WX5902, WX5904, WX5906, WX5908, WX5910,
         WX5913, WX5912, WX5915, WX5914, WX5917, WX5916, WX5919, WX5918,
         WX5921, WX5920, WX5923, WX5922, WX5925, WX5924, WX5927, WX5926,
         WX5929, WX5928, WX5931, WX5930, WX5933, WX5932, WX5935, WX5934,
         WX5937, WX5936, WX5939, WX5938, WX5941, WX5940, WX5943, WX5942,
         WX5945, WX5944, WX5947, WX5946, WX5949, WX5948, WX5951, WX5950,
         WX5953, WX5952, WX5955, WX5954, WX5957, WX5956, WX5959, WX5958,
         WX5961, WX5960, WX5963, WX5962, WX5965, WX5964, WX5967, WX5966,
         WX5969, WX5968, WX5971, WX5970, WX5973, WX5972, WX5975, WX5974,
         WX5977, WX5976, WX5979, WX5978, WX5981, WX5980, WX5983, WX5982,
         WX5985, WX5984, WX5987, WX5986, WX5989, WX5988, WX5991, WX5990,
         WX5993, WX5992, WX5995, WX5994, WX5997, WX5996, WX5999, WX5998,
         WX6001, WX6000, WX6003, WX6002, WX6005, WX6004, WX6007, WX6006,
         WX6009, WX6008, WX6011, WX6010, WX6013, WX6012, WX6015, WX6014,
         WX6017, WX6016, WX6019, WX6018, WX6021, WX6020, WX6023, WX6022,
         WX6025, WX6024, WX6027, WX6026, WX6029, WX6028, WX6031, WX6030,
         WX6033, WX6032, WX6035, WX6034, WX6037, WX6036, WX6039, WX6038,
         WX6041, WX6040, WX6043, WX6042, WX6045, WX6044, WX6047, WX6046,
         WX6049, WX6048, WX6051, WX6050, WX6053, WX6052, WX6055, WX6054,
         WX6057, WX6056, WX6059, WX6058, WX6061, WX6060, WX6063, WX6062,
         WX6065, WX6064, WX6067, WX6066, WX6069, WX6068, WX6071, WX6070,
         WX6436, WX6438, WX6440, WX6442, WX6444, WX6446, WX6448, WX6450,
         WX6452, WX6454, WX6456, WX6458, WX6460, WX6462, WX6464, WX6466,
         WX6468, WX6470, WX6472, WX6474, WX6476, WX6478, WX6480, WX6482,
         WX6484, WX6486, WX6488, WX6490, WX6492, WX6494, WX6496, WX6498,
         WX6950, WX6949, WX6952, WX6951, WX6954, WX6953, WX6956, WX6955,
         WX6958, WX6957, WX6960, WX6959, WX6962, WX6961, WX6964, WX6963,
         WX6966, WX6965, WX6968, WX6967, WX6970, WX6969, WX6972, WX6971,
         WX6974, WX6973, WX6976, WX6975, WX6978, WX6977, WX6980, WX6979,
         WX6982, WX6981, WX6984, WX6983, WX6986, WX6985, WX6988, WX6987,
         WX6990, WX6989, WX6992, WX6991, WX6994, WX6993, WX6996, WX6995,
         WX6998, WX6997, WX7000, WX6999, WX7002, WX7001, WX7004, WX7003,
         WX7006, WX7005, WX7008, WX7007, WX7010, WX7009, WX7012, WX7011,
         WX7110, WX7109, WX7112, WX7111, WX7114, WX7113, WX7116, WX7115,
         WX7118, WX7117, WX7120, WX7119, WX7122, WX7121, WX7124, WX7123,
         WX7126, WX7125, WX7128, WX7127, WX7130, WX7129, WX7132, WX7131,
         WX7134, WX7133, WX7136, WX7135, WX7138, WX7137, WX7140, WX7139,
         WX7141, WX7143, WX7145, WX7147, WX7149, WX7151, WX7153, WX7155,
         WX7157, WX7159, WX7161, WX7163, WX7165, WX7167, WX7169, WX7171,
         WX7173, WX7175, WX7177, WX7179, WX7181, WX7183, WX7185, WX7187,
         WX7189, WX7191, WX7193, WX7195, WX7197, WX7199, WX7201, WX7203,
         WX7206, WX7205, WX7208, WX7207, WX7210, WX7209, WX7212, WX7211,
         WX7214, WX7213, WX7216, WX7215, WX7218, WX7217, WX7220, WX7219,
         WX7222, WX7221, WX7224, WX7223, WX7226, WX7225, WX7228, WX7227,
         WX7230, WX7229, WX7232, WX7231, WX7234, WX7233, WX7236, WX7235,
         WX7238, WX7237, WX7240, WX7239, WX7242, WX7241, WX7244, WX7243,
         WX7246, WX7245, WX7248, WX7247, WX7250, WX7249, WX7252, WX7251,
         WX7254, WX7253, WX7256, WX7255, WX7258, WX7257, WX7260, WX7259,
         WX7262, WX7261, WX7264, WX7263, WX7266, WX7265, WX7268, WX7267,
         WX7270, WX7269, WX7272, WX7271, WX7274, WX7273, WX7276, WX7275,
         WX7278, WX7277, WX7280, WX7279, WX7282, WX7281, WX7284, WX7283,
         WX7286, WX7285, WX7288, WX7287, WX7290, WX7289, WX7292, WX7291,
         WX7294, WX7293, WX7296, WX7295, WX7298, WX7297, WX7300, WX7299,
         WX7302, WX7301, WX7304, WX7303, WX7306, WX7305, WX7308, WX7307,
         WX7310, WX7309, WX7312, WX7311, WX7314, WX7313, WX7316, WX7315,
         WX7318, WX7317, WX7320, WX7319, WX7322, WX7321, WX7324, WX7323,
         WX7326, WX7325, WX7328, WX7327, WX7330, WX7329, WX7332, WX7331,
         WX7334, WX7333, WX7336, WX7335, WX7338, WX7337, WX7340, WX7339,
         WX7342, WX7341, WX7344, WX7343, WX7346, WX7345, WX7348, WX7347,
         WX7350, WX7349, WX7352, WX7351, WX7354, WX7353, WX7356, WX7355,
         WX7358, WX7357, WX7360, WX7359, WX7362, WX7361, WX7364, WX7363,
         WX7729, WX7731, WX7733, WX7735, WX7737, WX7739, WX7741, WX7743,
         WX7745, WX7747, WX7749, WX7751, WX7753, WX7755, WX7757, WX7759,
         WX7761, WX7763, WX7765, WX7767, WX7769, WX7771, WX7773, WX7775,
         WX7777, WX7779, WX7781, WX7783, WX7785, WX7787, WX7789, WX7791,
         WX8243, WX8242, WX8245, WX8244, WX8247, WX8246, WX8249, WX8248,
         WX8251, WX8250, WX8253, WX8252, WX8255, WX8254, WX8257, WX8256,
         WX8259, WX8258, WX8261, WX8260, WX8263, WX8262, WX8265, WX8264,
         WX8267, WX8266, WX8269, WX8268, WX8271, WX8270, WX8273, WX8272,
         WX8275, WX8274, WX8277, WX8276, WX8279, WX8278, WX8281, WX8280,
         WX8283, WX8282, WX8285, WX8284, WX8287, WX8286, WX8289, WX8288,
         WX8291, WX8290, WX8293, WX8292, WX8295, WX8294, WX8297, WX8296,
         WX8299, WX8298, WX8301, WX8300, WX8303, WX8302, WX8305, WX8304,
         WX8403, WX8402, WX8405, WX8404, WX8407, WX8406, WX8409, WX8408,
         WX8411, WX8410, WX8413, WX8412, WX8415, WX8414, WX8417, WX8416,
         WX8419, WX8418, WX8421, WX8420, WX8423, WX8422, WX8425, WX8424,
         WX8427, WX8426, WX8429, WX8428, WX8431, WX8430, WX8433, WX8432,
         WX8434, WX8436, WX8438, WX8440, WX8442, WX8444, WX8446, WX8448,
         WX8450, WX8452, WX8454, WX8456, WX8458, WX8460, WX8462, WX8464,
         WX8466, WX8468, WX8470, WX8472, WX8474, WX8476, WX8478, WX8480,
         WX8482, WX8484, WX8486, WX8488, WX8490, WX8492, WX8494, WX8496,
         WX8499, WX8498, WX8501, WX8500, WX8503, WX8502, WX8505, WX8504,
         WX8507, WX8506, WX8509, WX8508, WX8511, WX8510, WX8513, WX8512,
         WX8515, WX8514, WX8517, WX8516, WX8519, WX8518, WX8521, WX8520,
         WX8523, WX8522, WX8525, WX8524, WX8527, WX8526, WX8529, WX8528,
         WX8531, WX8530, WX8533, WX8532, WX8535, WX8534, WX8537, WX8536,
         WX8539, WX8538, WX8541, WX8540, WX8543, WX8542, WX8545, WX8544,
         WX8547, WX8546, WX8549, WX8548, WX8551, WX8550, WX8553, WX8552,
         WX8555, WX8554, WX8557, WX8556, WX8559, WX8558, WX8561, WX8560,
         WX8563, WX8562, WX8565, WX8564, WX8567, WX8566, WX8569, WX8568,
         WX8571, WX8570, WX8573, WX8572, WX8575, WX8574, WX8577, WX8576,
         WX8579, WX8578, WX8581, WX8580, WX8583, WX8582, WX8585, WX8584,
         WX8587, WX8586, WX8589, WX8588, WX8591, WX8590, WX8593, WX8592,
         WX8595, WX8594, WX8597, WX8596, WX8599, WX8598, WX8601, WX8600,
         WX8603, WX8602, WX8605, WX8604, WX8607, WX8606, WX8609, WX8608,
         WX8611, WX8610, WX8613, WX8612, WX8615, WX8614, WX8617, WX8616,
         WX8619, WX8618, WX8621, WX8620, WX8623, WX8622, WX8625, WX8624,
         WX8627, WX8626, WX8629, WX8628, WX8631, WX8630, WX8633, WX8632,
         WX8635, WX8634, WX8637, WX8636, WX8639, WX8638, WX8641, WX8640,
         WX8643, WX8642, WX8645, WX8644, WX8647, WX8646, WX8649, WX8648,
         WX8651, WX8650, WX8653, WX8652, WX8655, WX8654, WX8657, WX8656,
         WX9022, WX9024, WX9026, WX9028, WX9030, WX9032, WX9034, WX9036,
         WX9038, WX9040, WX9042, WX9044, WX9046, WX9048, WX9050, WX9052,
         WX9054, WX9056, WX9058, WX9060, WX9062, WX9064, WX9066, WX9068,
         WX9070, WX9072, WX9074, WX9076, WX9078, WX9080, WX9082, WX9084,
         WX9536, WX9535, WX9538, WX9537, WX9540, WX9539, WX9542, WX9541,
         WX9544, WX9543, WX9546, WX9545, WX9548, WX9547, WX9550, WX9549,
         WX9552, WX9551, WX9554, WX9553, WX9556, WX9555, WX9558, WX9557,
         WX9560, WX9559, WX9562, WX9561, WX9564, WX9563, WX9566, WX9565,
         WX9568, WX9567, WX9570, WX9569, WX9572, WX9571, WX9574, WX9573,
         WX9576, WX9575, WX9578, WX9577, WX9580, WX9579, WX9582, WX9581,
         WX9584, WX9583, WX9586, WX9585, WX9588, WX9587, WX9590, WX9589,
         WX9592, WX9591, WX9594, WX9593, WX9596, WX9595, WX9598, WX9597,
         WX9696, WX9695, WX9698, WX9697, WX9700, WX9699, WX9702, WX9701,
         WX9704, WX9703, WX9706, WX9705, WX9708, WX9707, WX9710, WX9709,
         WX9712, WX9711, WX9714, WX9713, WX9716, WX9715, WX9718, WX9717,
         WX9720, WX9719, WX9722, WX9721, WX9724, WX9723, WX9726, WX9725,
         WX9727, WX9729, WX9731, WX9733, WX9735, WX9737, WX9739, WX9741,
         WX9743, WX9745, WX9747, WX9749, WX9751, WX9753, WX9755, WX9757,
         WX9759, WX9761, WX9763, WX9765, WX9767, WX9769, WX9771, WX9773,
         WX9775, WX9777, WX9779, WX9781, WX9783, WX9785, WX9787, WX9789,
         WX9792, WX9791, WX9794, WX9793, WX9796, WX9795, WX9798, WX9797,
         WX9800, WX9799, WX9802, WX9801, WX9804, WX9803, WX9806, WX9805,
         WX9808, WX9807, WX9810, WX9809, WX9812, WX9811, WX9814, WX9813,
         WX9816, WX9815, WX9818, WX9817, WX9820, WX9819, WX9822, WX9821,
         WX9824, WX9823, WX9826, WX9825, WX9828, WX9827, WX9830, WX9829,
         WX9832, WX9831, WX9834, WX9833, WX9836, WX9835, WX9838, WX9837,
         WX9840, WX9839, WX9842, WX9841, WX9844, WX9843, WX9846, WX9845,
         WX9848, WX9847, WX9850, WX9849, WX9852, WX9851, WX9854, WX9853,
         WX9856, WX9855, WX9858, WX9857, WX9860, WX9859, WX9862, WX9861,
         WX9864, WX9863, WX9866, WX9865, WX9868, WX9867, WX9870, WX9869,
         WX9872, WX9871, WX9874, WX9873, WX9876, WX9875, WX9878, WX9877,
         WX9880, WX9879, WX9882, WX9881, WX9884, WX9883, WX9886, WX9885,
         WX9888, WX9887, WX9890, WX9889, WX9892, WX9891, WX9894, WX9893,
         WX9896, WX9895, WX9898, WX9897, WX9900, WX9899, WX9902, WX9901,
         WX9904, WX9903, WX9906, WX9905, WX9908, WX9907, WX9910, WX9909,
         WX9912, WX9911, WX9914, WX9913, WX9916, WX9915, WX9918, WX9917,
         WX9920, WX9919, WX9922, WX9921, WX9924, WX9923, WX9926, WX9925,
         WX9928, WX9927, WX9930, WX9929, WX9932, WX9931, WX9934, WX9933,
         WX9936, WX9935, WX9938, WX9937, WX9940, WX9939, WX9942, WX9941,
         WX9944, WX9943, WX9946, WX9945, WX9948, WX9947, WX9950, WX9949,
         WX10315, WX10317, WX10319, WX10321, WX10323, WX10325, WX10327,
         WX10329, WX10331, WX10333, WX10335, WX10337, WX10339, WX10341,
         WX10343, WX10345, WX10347, WX10349, WX10351, WX10353, WX10355,
         WX10357, WX10359, WX10361, WX10363, WX10365, WX10367, WX10369,
         WX10371, WX10373, WX10375, WX10377, WX10829, WX10828, WX10831,
         WX10830, WX10833, WX10832, WX10835, WX10834, WX10837, WX10836,
         WX10839, WX10838, WX10841, WX10840, WX10843, WX10842, WX10845,
         WX10844, WX10847, WX10846, WX10849, WX10848, WX10851, WX10850,
         WX10853, WX10852, WX10855, WX10854, WX10857, WX10856, WX10859,
         WX10858, WX10861, WX10860, WX10863, WX10862, WX10865, WX10864,
         WX10867, WX10866, WX10869, WX10868, WX10871, WX10870, WX10873,
         WX10872, WX10875, WX10874, WX10877, WX10876, WX10879, WX10878,
         WX10881, WX10880, WX10883, WX10882, WX10885, WX10884, WX10887,
         WX10886, WX10889, WX10888, WX10891, WX10890, WX10989, WX10988,
         WX10991, WX10990, WX10993, WX10992, WX10995, WX10994, WX10997,
         WX10996, WX10999, WX10998, WX11001, WX11000, WX11003, WX11002,
         WX11005, WX11004, WX11007, WX11006, WX11009, WX11008, WX11011,
         WX11010, WX11013, WX11012, WX11015, WX11014, WX11017, WX11016,
         WX11019, WX11018, WX11021, WX11020, WX11023, WX11022, WX11025,
         WX11024, WX11027, WX11026, WX11029, WX11028, WX11031, WX11030,
         WX11033, WX11032, WX11035, WX11034, WX11037, WX11036, WX11039,
         WX11038, WX11041, WX11040, WX11043, WX11042, WX11045, WX11044,
         WX11047, WX11046, WX11049, WX11048, WX11051, WX11050, WX11052,
         WX11054, WX11056, WX11058, WX11060, WX11062, WX11064, WX11066,
         WX11068, WX11070, WX11072, WX11074, WX11076, WX11078, WX11080,
         WX11082, WX11084, WX11086, WX11088, WX11090, WX11092, WX11094,
         WX11096, WX11098, WX11100, WX11102, WX11104, WX11106, WX11108,
         WX11110, WX11112, WX11114, WX11117, WX11116, WX11119, WX11118,
         WX11121, WX11120, WX11123, WX11122, WX11125, WX11124, WX11127,
         WX11126, WX11129, WX11128, WX11131, WX11130, WX11133, WX11132,
         WX11135, WX11134, WX11137, WX11136, WX11139, WX11138, WX11141,
         WX11140, WX11143, WX11142, WX11145, WX11144, WX11147, WX11146,
         WX11149, WX11148, WX11151, WX11150, WX11153, WX11152, WX11155,
         WX11154, WX11157, WX11156, WX11159, WX11158, WX11161, WX11160,
         WX11163, WX11162, WX11165, WX11164, WX11167, WX11166, WX11169,
         WX11168, WX11171, WX11170, WX11173, WX11172, WX11175, WX11174,
         WX11177, WX11176, WX11179, WX11178, WX11181, WX11180, WX11183,
         WX11182, WX11185, WX11184, WX11187, WX11186, WX11189, WX11188,
         WX11191, WX11190, WX11193, WX11192, WX11195, WX11194, WX11197,
         WX11196, WX11199, WX11198, WX11201, WX11200, WX11203, WX11202,
         WX11205, WX11204, WX11207, WX11206, WX11209, WX11208, WX11211,
         WX11210, WX11213, WX11212, WX11215, WX11214, WX11217, WX11216,
         WX11219, WX11218, WX11221, WX11220, WX11223, WX11222, WX11225,
         WX11224, WX11227, WX11226, WX11229, WX11228, WX11231, WX11230,
         WX11233, WX11232, WX11235, WX11234, WX11237, WX11236, WX11239,
         WX11238, WX11241, WX11240, WX11243, WX11242, WX11608, WX11610,
         WX11612, WX11614, WX11616, WX11618, WX11620, WX11622, WX11624,
         WX11626, WX11628, WX11630, WX11632, WX11634, WX11636, WX11638,
         WX11640, WX11642, WX11644, WX11646, WX11648, WX11650, WX11652,
         WX11654, WX11656, WX11658, WX11660, WX11662, WX11664, WX11666,
         WX11668, WX11670, WX1010, WX1017, WX1024, WX1031, WX1038, WX1045,
         WX1052, WX1059, WX1066, WX1073, WX1080, WX1087, WX1094, WX1101,
         WX1108, WX1115, WX1122, WX1129, WX1136, WX1143, WX1150, WX1157,
         WX1164, WX1171, WX1178, WX1185, WX1192, WX1199, WX1206, WX1213,
         WX1220, WX1227, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148;
  assign DATA_9_31 = WX1010;
  assign DATA_9_30 = WX1017;
  assign DATA_9_29 = WX1024;
  assign DATA_9_28 = WX1031;
  assign DATA_9_27 = WX1038;
  assign DATA_9_26 = WX1045;
  assign DATA_9_25 = WX1052;
  assign DATA_9_24 = WX1059;
  assign DATA_9_23 = WX1066;
  assign DATA_9_22 = WX1073;
  assign DATA_9_21 = WX1080;
  assign DATA_9_20 = WX1087;
  assign DATA_9_19 = WX1094;
  assign DATA_9_18 = WX1101;
  assign DATA_9_17 = WX1108;
  assign DATA_9_16 = WX1115;
  assign DATA_9_15 = WX1122;
  assign DATA_9_14 = WX1129;
  assign DATA_9_13 = WX1136;
  assign DATA_9_12 = WX1143;
  assign DATA_9_11 = WX1150;
  assign DATA_9_10 = WX1157;
  assign DATA_9_9 = WX1164;
  assign DATA_9_8 = WX1171;
  assign DATA_9_7 = WX1178;
  assign DATA_9_6 = WX1185;
  assign DATA_9_5 = WX1192;
  assign DATA_9_4 = WX1199;
  assign DATA_9_3 = WX1206;
  assign DATA_9_2 = WX1213;
  assign DATA_9_1 = WX1220;
  assign DATA_9_0 = WX1227;

  hi1s1 U4709 ( .Q(n3333), .DIN(n4001) );
  hi1s1 U4710 ( .Q(n3334), .DIN(n3333) );
  hi1s1 U4711 ( .Q(n3335), .DIN(n3993) );
  hi1s1 U4712 ( .Q(n3336), .DIN(n3335) );
  hi1s1 U4713 ( .Q(n3337), .DIN(n4009) );
  hi1s1 U4714 ( .Q(n3338), .DIN(n3337) );
  hi1s1 U4715 ( .Q(n3339), .DIN(n3985) );
  hi1s1 U4716 ( .Q(n3340), .DIN(n3339) );
  hi1s1 U4717 ( .Q(n3341), .DIN(n4017) );
  hi1s1 U4718 ( .Q(n3342), .DIN(n3341) );
  hi1s1 U4719 ( .Q(n3343), .DIN(n3977) );
  hi1s1 U4720 ( .Q(n3344), .DIN(n3343) );
  hi1s1 U4721 ( .Q(n3345), .DIN(n4025) );
  hi1s1 U4722 ( .Q(n3346), .DIN(n3345) );
  hi1s1 U4723 ( .Q(n3347), .DIN(n3969) );
  hi1s1 U4724 ( .Q(n3348), .DIN(n3347) );
  hi1s1 U4725 ( .Q(n3349), .DIN(n4033) );
  hi1s1 U4726 ( .Q(n3350), .DIN(n3349) );
  hi1s1 U4727 ( .Q(n3351), .DIN(n3961) );
  hi1s1 U4728 ( .Q(n3352), .DIN(n3351) );
  hi1s1 U4729 ( .Q(n3353), .DIN(n4041) );
  hi1s1 U4730 ( .Q(n3354), .DIN(n3353) );
  hi1s1 U4731 ( .Q(n3355), .DIN(n3953) );
  hi1s1 U4732 ( .Q(n3356), .DIN(n3355) );
  hi1s1 U4733 ( .Q(n3357), .DIN(n6147) );
  hi1s1 U4734 ( .Q(n3358), .DIN(n3357) );
  hi1s1 U4735 ( .Q(n3359), .DIN(n3945) );
  hi1s1 U4736 ( .Q(n3360), .DIN(n3359) );
  hi1s1 U4737 ( .Q(n3362), .DIN(TM0) );
  hi1s1 U4738 ( .Q(n3361), .DIN(TM0) );
  hi1s1 U4739 ( .Q(n3363), .DIN(RESET) );
  hi1s1 U4740 ( .Q(n3364), .DIN(RESET) );
  hi1s1 U4741 ( .Q(n3365), .DIN(RESET) );
  hi1s1 U4742 ( .Q(n3366), .DIN(RESET) );
  hi1s1 U4743 ( .Q(n3367), .DIN(RESET) );
  hi1s1 U4744 ( .Q(n3368), .DIN(n3432) );
  hi1s1 U4745 ( .Q(n3369), .DIN(n3432) );
  hi1s1 U4746 ( .Q(n3370), .DIN(n3432) );
  hi1s1 U4747 ( .Q(n3371), .DIN(n3431) );
  hi1s1 U4748 ( .Q(n3372), .DIN(n3431) );
  hi1s1 U4749 ( .Q(n3373), .DIN(n3431) );
  hi1s1 U4750 ( .Q(n3374), .DIN(n3430) );
  hi1s1 U4751 ( .Q(n3375), .DIN(n3430) );
  hi1s1 U4752 ( .Q(n3376), .DIN(n3430) );
  hi1s1 U4753 ( .Q(n3377), .DIN(n3429) );
  hi1s1 U4754 ( .Q(n3378), .DIN(n3429) );
  hi1s1 U4755 ( .Q(n3379), .DIN(n3429) );
  hi1s1 U4756 ( .Q(n3380), .DIN(n3428) );
  hi1s1 U4757 ( .Q(n3381), .DIN(n3428) );
  hi1s1 U4758 ( .Q(n3382), .DIN(n3428) );
  hi1s1 U4759 ( .Q(n3383), .DIN(n3427) );
  hi1s1 U4760 ( .Q(n3384), .DIN(n3427) );
  hi1s1 U4761 ( .Q(n3385), .DIN(n3427) );
  hi1s1 U4762 ( .Q(n3386), .DIN(n3426) );
  hi1s1 U4763 ( .Q(n3387), .DIN(n3426) );
  hi1s1 U4764 ( .Q(n3388), .DIN(n3426) );
  hi1s1 U4765 ( .Q(n3389), .DIN(n3425) );
  hi1s1 U4766 ( .Q(n3390), .DIN(n3425) );
  hi1s1 U4767 ( .Q(n3391), .DIN(n3425) );
  hi1s1 U4768 ( .Q(n3392), .DIN(n3424) );
  hi1s1 U4769 ( .Q(n3393), .DIN(n3424) );
  hi1s1 U4770 ( .Q(n3394), .DIN(n3424) );
  hi1s1 U4771 ( .Q(n3395), .DIN(n3423) );
  hi1s1 U4772 ( .Q(n3396), .DIN(n3423) );
  hi1s1 U4773 ( .Q(n3397), .DIN(n3423) );
  hi1s1 U4774 ( .Q(n3398), .DIN(RESET) );
  hi1s1 U4775 ( .Q(n3399), .DIN(RESET) );
  hi1s1 U4776 ( .Q(n3400), .DIN(RESET) );
  hi1s1 U4777 ( .Q(n3401), .DIN(RESET) );
  hi1s1 U4778 ( .Q(n3402), .DIN(RESET) );
  hi1s1 U4779 ( .Q(n3403), .DIN(RESET) );
  hi1s1 U4780 ( .Q(n3404), .DIN(RESET) );
  hi1s1 U4781 ( .Q(n3405), .DIN(RESET) );
  hi1s1 U4782 ( .Q(n3406), .DIN(RESET) );
  hi1s1 U4783 ( .Q(n3407), .DIN(n3422) );
  hi1s1 U4784 ( .Q(n3408), .DIN(n3422) );
  hi1s1 U4785 ( .Q(n3409), .DIN(n3422) );
  hi1s1 U4786 ( .Q(n3410), .DIN(n3421) );
  hi1s1 U4787 ( .Q(n3411), .DIN(n3421) );
  hi1s1 U4788 ( .Q(n3412), .DIN(n3421) );
  hi1s1 U4789 ( .Q(n3413), .DIN(n3420) );
  hi1s1 U4790 ( .Q(n3414), .DIN(n3420) );
  hi1s1 U4791 ( .Q(n3415), .DIN(n3420) );
  hi1s1 U4792 ( .Q(n3416), .DIN(n3419) );
  hi1s1 U4793 ( .Q(n3417), .DIN(n3419) );
  hi1s1 U4794 ( .Q(n3418), .DIN(n3419) );
  hi1s1 U4795 ( .Q(n3419), .DIN(n3587) );
  hi1s1 U4796 ( .Q(n3420), .DIN(n3587) );
  hi1s1 U4797 ( .Q(n3421), .DIN(n3587) );
  hi1s1 U4798 ( .Q(n3422), .DIN(n3587) );
  hi1s1 U4799 ( .Q(n3423), .DIN(n3587) );
  hi1s1 U4800 ( .Q(n3424), .DIN(n3587) );
  hi1s1 U4801 ( .Q(n3425), .DIN(n3587) );
  hi1s1 U4802 ( .Q(n3426), .DIN(n3587) );
  hi1s1 U4803 ( .Q(n3427), .DIN(n3587) );
  hi1s1 U4804 ( .Q(n3428), .DIN(n3587) );
  hi1s1 U4805 ( .Q(n3429), .DIN(n3587) );
  hi1s1 U4806 ( .Q(n3430), .DIN(n3587) );
  hi1s1 U4807 ( .Q(n3431), .DIN(n3587) );
  hi1s1 U4808 ( .Q(n3432), .DIN(n3587) );
  hi1s1 U4809 ( .Q(n3433), .DIN(n3463) );
  hi1s1 U4810 ( .Q(n3434), .DIN(n3463) );
  hi1s1 U4811 ( .Q(n3435), .DIN(n3462) );
  hi1s1 U4812 ( .Q(n3436), .DIN(n3462) );
  hi1s1 U4813 ( .Q(n3437), .DIN(n3462) );
  hi1s1 U4814 ( .Q(n3438), .DIN(n3461) );
  hi1s1 U4815 ( .Q(n3439), .DIN(n3461) );
  hi1s1 U4816 ( .Q(n3440), .DIN(n3461) );
  hi1s1 U4817 ( .Q(n3441), .DIN(n3460) );
  hi1s1 U4818 ( .Q(n3442), .DIN(n3460) );
  hi1s1 U4819 ( .Q(n3443), .DIN(n3460) );
  hi1s1 U4820 ( .Q(n3444), .DIN(n3459) );
  hi1s1 U4821 ( .Q(n3445), .DIN(n3459) );
  hi1s1 U4822 ( .Q(n3446), .DIN(n3459) );
  hi1s1 U4823 ( .Q(n3447), .DIN(n3458) );
  hi1s1 U4824 ( .Q(n3448), .DIN(n3458) );
  hi1s1 U4825 ( .Q(n3449), .DIN(n3458) );
  hi1s1 U4826 ( .Q(n3450), .DIN(n3457) );
  hi1s1 U4827 ( .Q(n3451), .DIN(n3457) );
  hi1s1 U4828 ( .Q(n3452), .DIN(n3457) );
  hi1s1 U4829 ( .Q(n3453), .DIN(n3456) );
  hi1s1 U4830 ( .Q(n3454), .DIN(n3456) );
  hi1s1 U4831 ( .Q(n3455), .DIN(n3456) );
  hi1s1 U4832 ( .Q(n3456), .DIN(n3592) );
  hi1s1 U4833 ( .Q(n3457), .DIN(n3592) );
  hi1s1 U4834 ( .Q(n3458), .DIN(n3592) );
  hi1s1 U4835 ( .Q(n3459), .DIN(n3592) );
  hi1s1 U4836 ( .Q(n3460), .DIN(n3592) );
  hi1s1 U4837 ( .Q(n3461), .DIN(n3592) );
  hi1s1 U4838 ( .Q(n3462), .DIN(n3592) );
  hi1s1 U4839 ( .Q(n3463), .DIN(n3592) );
  hi1s1 U4840 ( .Q(n3464), .DIN(n3494) );
  hi1s1 U4841 ( .Q(n3465), .DIN(n3494) );
  hi1s1 U4842 ( .Q(n3466), .DIN(n3493) );
  hi1s1 U4843 ( .Q(n3467), .DIN(n3493) );
  hi1s1 U4844 ( .Q(n3468), .DIN(n3493) );
  hi1s1 U4845 ( .Q(n3469), .DIN(n3492) );
  hi1s1 U4846 ( .Q(n3470), .DIN(n3492) );
  hi1s1 U4847 ( .Q(n3471), .DIN(n3492) );
  hi1s1 U4848 ( .Q(n3472), .DIN(n3491) );
  hi1s1 U4849 ( .Q(n3473), .DIN(n3491) );
  hi1s1 U4850 ( .Q(n3474), .DIN(n3491) );
  hi1s1 U4851 ( .Q(n3475), .DIN(n3490) );
  hi1s1 U4852 ( .Q(n3476), .DIN(n3490) );
  hi1s1 U4853 ( .Q(n3477), .DIN(n3490) );
  hi1s1 U4854 ( .Q(n3478), .DIN(n3489) );
  hi1s1 U4855 ( .Q(n3479), .DIN(n3489) );
  hi1s1 U4856 ( .Q(n3480), .DIN(n3489) );
  hi1s1 U4857 ( .Q(n3481), .DIN(n3488) );
  hi1s1 U4858 ( .Q(n3482), .DIN(n3488) );
  hi1s1 U4859 ( .Q(n3483), .DIN(n3488) );
  hi1s1 U4860 ( .Q(n3484), .DIN(n3487) );
  hi1s1 U4861 ( .Q(n3485), .DIN(n3487) );
  hi1s1 U4862 ( .Q(n3486), .DIN(n3487) );
  hi1s1 U4863 ( .Q(n3487), .DIN(n3594) );
  hi1s1 U4864 ( .Q(n3488), .DIN(n3594) );
  hi1s1 U4865 ( .Q(n3489), .DIN(n3594) );
  hi1s1 U4866 ( .Q(n3490), .DIN(n3594) );
  hi1s1 U4867 ( .Q(n3491), .DIN(n3594) );
  hi1s1 U4868 ( .Q(n3492), .DIN(n3594) );
  hi1s1 U4869 ( .Q(n3493), .DIN(n3594) );
  hi1s1 U4870 ( .Q(n3494), .DIN(n3594) );
  hi1s1 U4871 ( .Q(n3495), .DIN(n3526) );
  hi1s1 U4872 ( .Q(n3496), .DIN(n3526) );
  hi1s1 U4873 ( .Q(n3497), .DIN(n3526) );
  hi1s1 U4874 ( .Q(n3498), .DIN(n3525) );
  hi1s1 U4875 ( .Q(n3499), .DIN(n3525) );
  hi1s1 U4876 ( .Q(n3500), .DIN(n3525) );
  hi1s1 U4877 ( .Q(n3501), .DIN(n3524) );
  hi1s1 U4878 ( .Q(n3502), .DIN(n3524) );
  hi1s1 U4879 ( .Q(n3503), .DIN(n3524) );
  hi1s1 U4880 ( .Q(n3504), .DIN(n3523) );
  hi1s1 U4881 ( .Q(n3505), .DIN(n3523) );
  hi1s1 U4882 ( .Q(n3506), .DIN(n3523) );
  hi1s1 U4883 ( .Q(n3507), .DIN(n3522) );
  hi1s1 U4884 ( .Q(n3508), .DIN(n3522) );
  hi1s1 U4885 ( .Q(n3509), .DIN(n3522) );
  hi1s1 U4886 ( .Q(n3510), .DIN(n3521) );
  hi1s1 U4887 ( .Q(n3511), .DIN(n3521) );
  hi1s1 U4888 ( .Q(n3512), .DIN(n3521) );
  hi1s1 U4889 ( .Q(n3513), .DIN(n3520) );
  hi1s1 U4890 ( .Q(n3514), .DIN(n3520) );
  hi1s1 U4891 ( .Q(n3515), .DIN(n3520) );
  hi1s1 U4892 ( .Q(n3516), .DIN(n3519) );
  hi1s1 U4893 ( .Q(n3517), .DIN(n3519) );
  hi1s1 U4894 ( .Q(n3518), .DIN(n3519) );
  hi1s1 U4895 ( .Q(n3519), .DIN(n3596) );
  hi1s1 U4896 ( .Q(n3520), .DIN(n3596) );
  hi1s1 U4897 ( .Q(n3521), .DIN(n3596) );
  hi1s1 U4898 ( .Q(n3522), .DIN(n3596) );
  hi1s1 U4899 ( .Q(n3523), .DIN(n3596) );
  hi1s1 U4900 ( .Q(n3524), .DIN(n3596) );
  hi1s1 U4901 ( .Q(n3525), .DIN(n3596) );
  hi1s1 U4902 ( .Q(n3526), .DIN(n3596) );
  hi1s1 U4903 ( .Q(n3527), .DIN(n3558) );
  hi1s1 U4904 ( .Q(n3528), .DIN(n3558) );
  hi1s1 U4905 ( .Q(n3529), .DIN(n3558) );
  hi1s1 U4906 ( .Q(n3530), .DIN(n3557) );
  hi1s1 U4907 ( .Q(n3531), .DIN(n3557) );
  hi1s1 U4908 ( .Q(n3532), .DIN(n3557) );
  hi1s1 U4909 ( .Q(n3533), .DIN(n3556) );
  hi1s1 U4910 ( .Q(n3534), .DIN(n3556) );
  hi1s1 U4911 ( .Q(n3535), .DIN(n3556) );
  hi1s1 U4912 ( .Q(n3536), .DIN(n3555) );
  hi1s1 U4913 ( .Q(n3537), .DIN(n3555) );
  hi1s1 U4914 ( .Q(n3538), .DIN(n3555) );
  hi1s1 U4915 ( .Q(n3539), .DIN(n3554) );
  hi1s1 U4916 ( .Q(n3540), .DIN(n3554) );
  hi1s1 U4917 ( .Q(n3541), .DIN(n3554) );
  hi1s1 U4918 ( .Q(n3542), .DIN(n3553) );
  hi1s1 U4919 ( .Q(n3543), .DIN(n3553) );
  hi1s1 U4920 ( .Q(n3544), .DIN(n3553) );
  hi1s1 U4921 ( .Q(n3545), .DIN(n3552) );
  hi1s1 U4922 ( .Q(n3546), .DIN(n3552) );
  hi1s1 U4923 ( .Q(n3547), .DIN(n3552) );
  hi1s1 U4924 ( .Q(n3548), .DIN(n3551) );
  hi1s1 U4925 ( .Q(n3549), .DIN(n3551) );
  hi1s1 U4926 ( .Q(n3550), .DIN(n3551) );
  hi1s1 U4927 ( .Q(n3551), .DIN(n3597) );
  hi1s1 U4928 ( .Q(n3552), .DIN(n3597) );
  hi1s1 U4929 ( .Q(n3553), .DIN(n3597) );
  hi1s1 U4930 ( .Q(n3554), .DIN(n3597) );
  hi1s1 U4931 ( .Q(n3555), .DIN(n3597) );
  hi1s1 U4932 ( .Q(n3556), .DIN(n3597) );
  hi1s1 U4933 ( .Q(n3557), .DIN(n3597) );
  hi1s1 U4934 ( .Q(n3558), .DIN(n3597) );
  hi1s1 U4935 ( .Q(n3559), .DIN(n3586) );
  hi1s1 U4936 ( .Q(n3560), .DIN(n3586) );
  hi1s1 U4937 ( .Q(n3561), .DIN(n3586) );
  hi1s1 U4938 ( .Q(n3562), .DIN(n3585) );
  hi1s1 U4939 ( .Q(n3563), .DIN(n3585) );
  hi1s1 U4940 ( .Q(n3564), .DIN(n3585) );
  hi1s1 U4941 ( .Q(n3565), .DIN(n3584) );
  hi1s1 U4942 ( .Q(n3566), .DIN(n3584) );
  hi1s1 U4943 ( .Q(n3567), .DIN(n3584) );
  hi1s1 U4944 ( .Q(n3568), .DIN(n3583) );
  hi1s1 U4945 ( .Q(n3569), .DIN(n3583) );
  hi1s1 U4946 ( .Q(n3570), .DIN(n3583) );
  hi1s1 U4947 ( .Q(n3571), .DIN(n3582) );
  hi1s1 U4948 ( .Q(n3572), .DIN(n3582) );
  hi1s1 U4949 ( .Q(n3573), .DIN(n3582) );
  hi1s1 U4950 ( .Q(n3574), .DIN(n3581) );
  hi1s1 U4951 ( .Q(n3575), .DIN(n3581) );
  hi1s1 U4952 ( .Q(n3576), .DIN(n3581) );
  hi1s1 U4953 ( .Q(n3577), .DIN(n3580) );
  hi1s1 U4954 ( .Q(n3578), .DIN(n3580) );
  hi1s1 U4955 ( .Q(n3579), .DIN(n3580) );
  hi1s1 U4956 ( .Q(n3580), .DIN(n3937) );
  hi1s1 U4957 ( .Q(n3581), .DIN(n3937) );
  hi1s1 U4958 ( .Q(n3582), .DIN(n3937) );
  hi1s1 U4959 ( .Q(n3583), .DIN(n3937) );
  hi1s1 U4960 ( .Q(n3584), .DIN(n3937) );
  hi1s1 U4961 ( .Q(n3585), .DIN(n3937) );
  hi1s1 U4962 ( .Q(n3586), .DIN(n3937) );
  and2s1 U4963 ( .Q(WX9949), .DIN1(RESET), .DIN2(WX9886) );
  and2s1 U4964 ( .Q(WX9947), .DIN1(RESET), .DIN2(WX9884) );
  and2s1 U4965 ( .Q(WX9945), .DIN1(RESET), .DIN2(WX9882) );
  and2s1 U4966 ( .Q(WX9943), .DIN1(RESET), .DIN2(WX9880) );
  and2s1 U4967 ( .Q(WX9941), .DIN1(RESET), .DIN2(WX9878) );
  and2s1 U4968 ( .Q(WX9939), .DIN1(RESET), .DIN2(WX9876) );
  and2s1 U4969 ( .Q(WX9937), .DIN1(RESET), .DIN2(WX9874) );
  and2s1 U4970 ( .Q(WX9935), .DIN1(RESET), .DIN2(WX9872) );
  and2s1 U4971 ( .Q(WX9933), .DIN1(RESET), .DIN2(WX9870) );
  and2s1 U4972 ( .Q(WX9931), .DIN1(RESET), .DIN2(WX9868) );
  and2s1 U4973 ( .Q(WX9929), .DIN1(RESET), .DIN2(WX9866) );
  and2s1 U4974 ( .Q(WX9927), .DIN1(RESET), .DIN2(WX9864) );
  and2s1 U4975 ( .Q(WX9925), .DIN1(RESET), .DIN2(WX9862) );
  and2s1 U4976 ( .Q(WX9923), .DIN1(RESET), .DIN2(WX9860) );
  and2s1 U4977 ( .Q(WX9921), .DIN1(RESET), .DIN2(WX9858) );
  and2s1 U4978 ( .Q(WX9919), .DIN1(RESET), .DIN2(WX9856) );
  and2s1 U4979 ( .Q(WX9917), .DIN1(RESET), .DIN2(WX9854) );
  and2s1 U4980 ( .Q(WX9915), .DIN1(RESET), .DIN2(WX9852) );
  and2s1 U4981 ( .Q(WX9913), .DIN1(RESET), .DIN2(WX9850) );
  and2s1 U4982 ( .Q(WX9911), .DIN1(RESET), .DIN2(WX9848) );
  and2s1 U4983 ( .Q(WX9909), .DIN1(RESET), .DIN2(WX9846) );
  and2s1 U4984 ( .Q(WX9907), .DIN1(RESET), .DIN2(WX9844) );
  and2s1 U4985 ( .Q(WX9905), .DIN1(RESET), .DIN2(WX9842) );
  and2s1 U4986 ( .Q(WX9903), .DIN1(RESET), .DIN2(WX9840) );
  and2s1 U4987 ( .Q(WX9901), .DIN1(RESET), .DIN2(WX9838) );
  and2s1 U4988 ( .Q(WX9899), .DIN1(RESET), .DIN2(WX9836) );
  and2s1 U4989 ( .Q(WX9897), .DIN1(RESET), .DIN2(WX9834) );
  and2s1 U4990 ( .Q(WX9895), .DIN1(RESET), .DIN2(WX9832) );
  and2s1 U4991 ( .Q(WX9893), .DIN1(RESET), .DIN2(WX9830) );
  and2s1 U4992 ( .Q(WX9891), .DIN1(RESET), .DIN2(WX9828) );
  and2s1 U4993 ( .Q(WX9889), .DIN1(RESET), .DIN2(WX9826) );
  and2s1 U4994 ( .Q(WX9887), .DIN1(RESET), .DIN2(WX9824) );
  and2s1 U4995 ( .Q(WX9885), .DIN1(RESET), .DIN2(WX9822) );
  and2s1 U4996 ( .Q(WX9883), .DIN1(RESET), .DIN2(WX9820) );
  and2s1 U4997 ( .Q(WX9881), .DIN1(RESET), .DIN2(WX9818) );
  and2s1 U4998 ( .Q(WX9879), .DIN1(RESET), .DIN2(WX9816) );
  and2s1 U4999 ( .Q(WX9877), .DIN1(RESET), .DIN2(WX9814) );
  and2s1 U5000 ( .Q(WX9875), .DIN1(RESET), .DIN2(WX9812) );
  and2s1 U5001 ( .Q(WX9873), .DIN1(RESET), .DIN2(WX9810) );
  and2s1 U5002 ( .Q(WX9871), .DIN1(RESET), .DIN2(WX9808) );
  and2s1 U5003 ( .Q(WX9869), .DIN1(RESET), .DIN2(WX9806) );
  and2s1 U5004 ( .Q(WX9867), .DIN1(RESET), .DIN2(WX9804) );
  and2s1 U5005 ( .Q(WX9865), .DIN1(RESET), .DIN2(WX9802) );
  and2s1 U5006 ( .Q(WX9863), .DIN1(RESET), .DIN2(WX9800) );
  and2s1 U5007 ( .Q(WX9861), .DIN1(RESET), .DIN2(WX9798) );
  and2s1 U5008 ( .Q(WX9859), .DIN1(RESET), .DIN2(WX9796) );
  and2s1 U5009 ( .Q(WX9857), .DIN1(RESET), .DIN2(WX9794) );
  and2s1 U5010 ( .Q(WX9855), .DIN1(RESET), .DIN2(WX9792) );
  nor2s1 U5011 ( .Q(WX9853), .DIN1(n3390), .DIN2(n2949) );
  nor2s1 U5012 ( .Q(WX9851), .DIN1(n3383), .DIN2(n2950) );
  nor2s1 U5013 ( .Q(WX9849), .DIN1(n3377), .DIN2(n2951) );
  nor2s1 U5014 ( .Q(WX9847), .DIN1(n3377), .DIN2(n2952) );
  nor2s1 U5015 ( .Q(WX9845), .DIN1(n3377), .DIN2(n2953) );
  nor2s1 U5016 ( .Q(WX9843), .DIN1(n3377), .DIN2(n2954) );
  nor2s1 U5017 ( .Q(WX9841), .DIN1(n3377), .DIN2(n2955) );
  nor2s1 U5018 ( .Q(WX9839), .DIN1(n3377), .DIN2(n2956) );
  nor2s1 U5019 ( .Q(WX9837), .DIN1(n3377), .DIN2(n2957) );
  nor2s1 U5020 ( .Q(WX9835), .DIN1(n3377), .DIN2(n2958) );
  nor2s1 U5021 ( .Q(WX9833), .DIN1(n3378), .DIN2(n2959) );
  nor2s1 U5022 ( .Q(WX9831), .DIN1(n3378), .DIN2(n2960) );
  nor2s1 U5023 ( .Q(WX9829), .DIN1(n3378), .DIN2(n2961) );
  nor2s1 U5024 ( .Q(WX9827), .DIN1(n3378), .DIN2(n2962) );
  nor2s1 U5025 ( .Q(WX9825), .DIN1(n3378), .DIN2(n2963) );
  nor2s1 U5026 ( .Q(WX9823), .DIN1(n3378), .DIN2(n2964) );
  nor2s1 U5027 ( .Q(WX9821), .DIN1(n3378), .DIN2(n3109) );
  nor2s1 U5028 ( .Q(WX9819), .DIN1(n3378), .DIN2(n3110) );
  nor2s1 U5029 ( .Q(WX9817), .DIN1(n3378), .DIN2(n3111) );
  nor2s1 U5030 ( .Q(WX9815), .DIN1(n3378), .DIN2(n3112) );
  nor2s1 U5031 ( .Q(WX9813), .DIN1(n3379), .DIN2(n3113) );
  nor2s1 U5032 ( .Q(WX9811), .DIN1(n3379), .DIN2(n3114) );
  nor2s1 U5033 ( .Q(WX9809), .DIN1(n3379), .DIN2(n3115) );
  nor2s1 U5034 ( .Q(WX9807), .DIN1(n3379), .DIN2(n3116) );
  nor2s1 U5035 ( .Q(WX9805), .DIN1(n3379), .DIN2(n3117) );
  nor2s1 U5036 ( .Q(WX9803), .DIN1(n3379), .DIN2(n3118) );
  nor2s1 U5037 ( .Q(WX9801), .DIN1(n3379), .DIN2(n3119) );
  nor2s1 U5038 ( .Q(WX9799), .DIN1(n3379), .DIN2(n3120) );
  nor2s1 U5039 ( .Q(WX9797), .DIN1(n3379), .DIN2(n3121) );
  nor2s1 U5040 ( .Q(WX9795), .DIN1(n3379), .DIN2(n3122) );
  nor2s1 U5041 ( .Q(WX9793), .DIN1(n3380), .DIN2(n3123) );
  nor2s1 U5042 ( .Q(WX9791), .DIN1(n3380), .DIN2(n3124) );
  and2s1 U5043 ( .Q(WX9789), .DIN1(RESET), .DIN2(WX9726) );
  and2s1 U5044 ( .Q(WX9787), .DIN1(RESET), .DIN2(WX9724) );
  and2s1 U5045 ( .Q(WX9785), .DIN1(RESET), .DIN2(WX9722) );
  and2s1 U5046 ( .Q(WX9783), .DIN1(RESET), .DIN2(WX9720) );
  and2s1 U5047 ( .Q(WX9781), .DIN1(RESET), .DIN2(WX9718) );
  and2s1 U5048 ( .Q(WX9779), .DIN1(RESET), .DIN2(WX9716) );
  and2s1 U5049 ( .Q(WX9777), .DIN1(RESET), .DIN2(WX9714) );
  and2s1 U5050 ( .Q(WX9775), .DIN1(RESET), .DIN2(WX9712) );
  and2s1 U5051 ( .Q(WX9773), .DIN1(RESET), .DIN2(WX9710) );
  and2s1 U5052 ( .Q(WX9771), .DIN1(RESET), .DIN2(WX9708) );
  and2s1 U5053 ( .Q(WX9769), .DIN1(RESET), .DIN2(WX9706) );
  and2s1 U5054 ( .Q(WX9767), .DIN1(RESET), .DIN2(WX9704) );
  and2s1 U5055 ( .Q(WX9765), .DIN1(RESET), .DIN2(WX9702) );
  and2s1 U5056 ( .Q(WX9763), .DIN1(RESET), .DIN2(WX9700) );
  and2s1 U5057 ( .Q(WX9761), .DIN1(RESET), .DIN2(WX9698) );
  and2s1 U5058 ( .Q(WX9759), .DIN1(RESET), .DIN2(WX9696) );
  nnd4s1 U5059 ( .Q(WX9757), .DIN1(n3588), .DIN2(n3589), .DIN3(n3590), .DIN4(
        n3591) );
  nnd2s1 U5060 ( .Q(n3591), .DIN1(n3455), .DIN2(n3593) );
  nnd2s1 U5061 ( .Q(n3590), .DIN1(n3464), .DIN2(n3595) );
  nnd2s1 U5062 ( .Q(n3589), .DIN1(WX9598), .DIN2(n3518) );
  nnd2s1 U5063 ( .Q(n3588), .DIN1(CRC_OUT_2_0), .DIN2(n3550) );
  nnd4s1 U5064 ( .Q(WX9755), .DIN1(n3598), .DIN2(n3599), .DIN3(n3600), .DIN4(
        n3601) );
  nnd2s1 U5065 ( .Q(n3601), .DIN1(n3455), .DIN2(n3602) );
  nnd2s1 U5066 ( .Q(n3600), .DIN1(n3464), .DIN2(n3603) );
  nnd2s1 U5067 ( .Q(n3599), .DIN1(WX9596), .DIN2(n3518) );
  nnd2s1 U5068 ( .Q(n3598), .DIN1(CRC_OUT_2_1), .DIN2(n3550) );
  nnd4s1 U5069 ( .Q(WX9753), .DIN1(n3604), .DIN2(n3605), .DIN3(n3606), .DIN4(
        n3607) );
  nnd2s1 U5070 ( .Q(n3607), .DIN1(n3454), .DIN2(n3608) );
  nnd2s1 U5071 ( .Q(n3606), .DIN1(n3464), .DIN2(n3609) );
  nnd2s1 U5072 ( .Q(n3605), .DIN1(WX9594), .DIN2(n3518) );
  nnd2s1 U5073 ( .Q(n3604), .DIN1(CRC_OUT_2_2), .DIN2(n3550) );
  nnd4s1 U5074 ( .Q(WX9751), .DIN1(n3610), .DIN2(n3611), .DIN3(n3612), .DIN4(
        n3613) );
  nnd2s1 U5075 ( .Q(n3613), .DIN1(n3454), .DIN2(n3614) );
  nnd2s1 U5076 ( .Q(n3612), .DIN1(n3464), .DIN2(n3615) );
  nnd2s1 U5077 ( .Q(n3611), .DIN1(WX9592), .DIN2(n3518) );
  nnd2s1 U5078 ( .Q(n3610), .DIN1(CRC_OUT_2_3), .DIN2(n3550) );
  nnd4s1 U5079 ( .Q(WX9749), .DIN1(n3616), .DIN2(n3617), .DIN3(n3618), .DIN4(
        n3619) );
  nnd2s1 U5080 ( .Q(n3619), .DIN1(n3454), .DIN2(n3620) );
  nnd2s1 U5081 ( .Q(n3618), .DIN1(n3464), .DIN2(n3621) );
  nnd2s1 U5082 ( .Q(n3617), .DIN1(WX9590), .DIN2(n3518) );
  nnd2s1 U5083 ( .Q(n3616), .DIN1(CRC_OUT_2_4), .DIN2(n3550) );
  nnd4s1 U5084 ( .Q(WX9747), .DIN1(n3622), .DIN2(n3623), .DIN3(n3624), .DIN4(
        n3625) );
  nnd2s1 U5085 ( .Q(n3625), .DIN1(n3454), .DIN2(n3626) );
  nnd2s1 U5086 ( .Q(n3624), .DIN1(n3464), .DIN2(n3627) );
  nnd2s1 U5087 ( .Q(n3623), .DIN1(WX9588), .DIN2(n3518) );
  nnd2s1 U5088 ( .Q(n3622), .DIN1(CRC_OUT_2_5), .DIN2(n3550) );
  nnd4s1 U5089 ( .Q(WX9745), .DIN1(n3628), .DIN2(n3629), .DIN3(n3630), .DIN4(
        n3631) );
  nnd2s1 U5090 ( .Q(n3631), .DIN1(n3454), .DIN2(n3632) );
  nnd2s1 U5091 ( .Q(n3630), .DIN1(n3464), .DIN2(n3633) );
  nnd2s1 U5092 ( .Q(n3629), .DIN1(WX9586), .DIN2(n3518) );
  nnd2s1 U5093 ( .Q(n3628), .DIN1(CRC_OUT_2_6), .DIN2(n3550) );
  nnd4s1 U5094 ( .Q(WX9743), .DIN1(n3634), .DIN2(n3635), .DIN3(n3636), .DIN4(
        n3637) );
  nnd2s1 U5095 ( .Q(n3637), .DIN1(n3454), .DIN2(n3638) );
  nnd2s1 U5096 ( .Q(n3636), .DIN1(n3464), .DIN2(n3639) );
  nnd2s1 U5097 ( .Q(n3635), .DIN1(WX9584), .DIN2(n3518) );
  nnd2s1 U5098 ( .Q(n3634), .DIN1(CRC_OUT_2_7), .DIN2(n3550) );
  nnd4s1 U5099 ( .Q(WX9741), .DIN1(n3640), .DIN2(n3641), .DIN3(n3642), .DIN4(
        n3643) );
  nnd2s1 U5100 ( .Q(n3643), .DIN1(n3454), .DIN2(n3644) );
  nnd2s1 U5101 ( .Q(n3642), .DIN1(n3464), .DIN2(n3645) );
  nnd2s1 U5102 ( .Q(n3641), .DIN1(WX9582), .DIN2(n3518) );
  nnd2s1 U5103 ( .Q(n3640), .DIN1(CRC_OUT_2_8), .DIN2(n3550) );
  nnd4s1 U5104 ( .Q(WX9739), .DIN1(n3646), .DIN2(n3647), .DIN3(n3648), .DIN4(
        n3649) );
  nnd2s1 U5105 ( .Q(n3649), .DIN1(n3454), .DIN2(n3650) );
  nnd2s1 U5106 ( .Q(n3648), .DIN1(n3464), .DIN2(n3651) );
  nnd2s1 U5107 ( .Q(n3647), .DIN1(WX9580), .DIN2(n3518) );
  nnd2s1 U5108 ( .Q(n3646), .DIN1(CRC_OUT_2_9), .DIN2(n3550) );
  nnd4s1 U5109 ( .Q(WX9737), .DIN1(n3652), .DIN2(n3653), .DIN3(n3654), .DIN4(
        n3655) );
  nnd2s1 U5110 ( .Q(n3655), .DIN1(n3454), .DIN2(n3656) );
  nnd2s1 U5111 ( .Q(n3654), .DIN1(n3464), .DIN2(n3657) );
  nnd2s1 U5112 ( .Q(n3653), .DIN1(WX9578), .DIN2(n3518) );
  nnd2s1 U5113 ( .Q(n3652), .DIN1(CRC_OUT_2_10), .DIN2(n3550) );
  nnd4s1 U5114 ( .Q(WX9735), .DIN1(n3658), .DIN2(n3659), .DIN3(n3660), .DIN4(
        n3661) );
  nnd2s1 U5115 ( .Q(n3661), .DIN1(n3454), .DIN2(n3662) );
  nnd2s1 U5116 ( .Q(n3660), .DIN1(n3464), .DIN2(n3663) );
  nnd2s1 U5117 ( .Q(n3659), .DIN1(WX9576), .DIN2(n3518) );
  nnd2s1 U5118 ( .Q(n3658), .DIN1(CRC_OUT_2_11), .DIN2(n3550) );
  nnd4s1 U5119 ( .Q(WX9733), .DIN1(n3664), .DIN2(n3665), .DIN3(n3666), .DIN4(
        n3667) );
  nnd2s1 U5120 ( .Q(n3667), .DIN1(n3454), .DIN2(n3668) );
  nnd2s1 U5121 ( .Q(n3666), .DIN1(n3464), .DIN2(n3669) );
  nnd2s1 U5122 ( .Q(n3665), .DIN1(WX9574), .DIN2(n3517) );
  nnd2s1 U5123 ( .Q(n3664), .DIN1(CRC_OUT_2_12), .DIN2(n3549) );
  nnd4s1 U5124 ( .Q(WX9731), .DIN1(n3670), .DIN2(n3671), .DIN3(n3672), .DIN4(
        n3673) );
  nnd2s1 U5125 ( .Q(n3673), .DIN1(n3454), .DIN2(n3674) );
  nnd2s1 U5126 ( .Q(n3672), .DIN1(n3465), .DIN2(n3675) );
  nnd2s1 U5127 ( .Q(n3671), .DIN1(WX9572), .DIN2(n3517) );
  nnd2s1 U5128 ( .Q(n3670), .DIN1(CRC_OUT_2_13), .DIN2(n3549) );
  nnd4s1 U5129 ( .Q(WX9729), .DIN1(n3676), .DIN2(n3677), .DIN3(n3678), .DIN4(
        n3679) );
  nnd2s1 U5130 ( .Q(n3679), .DIN1(n3454), .DIN2(n3680) );
  nnd2s1 U5131 ( .Q(n3678), .DIN1(n3465), .DIN2(n3681) );
  nnd2s1 U5132 ( .Q(n3677), .DIN1(WX9570), .DIN2(n3517) );
  nnd2s1 U5133 ( .Q(n3676), .DIN1(CRC_OUT_2_14), .DIN2(n3549) );
  nnd4s1 U5134 ( .Q(WX9727), .DIN1(n3682), .DIN2(n3683), .DIN3(n3684), .DIN4(
        n3685) );
  nnd2s1 U5135 ( .Q(n3685), .DIN1(n3453), .DIN2(n3686) );
  nnd2s1 U5136 ( .Q(n3684), .DIN1(n3465), .DIN2(n3687) );
  nnd2s1 U5137 ( .Q(n3683), .DIN1(WX9568), .DIN2(n3517) );
  nnd2s1 U5138 ( .Q(n3682), .DIN1(CRC_OUT_2_15), .DIN2(n3549) );
  nnd4s1 U5139 ( .Q(WX9725), .DIN1(n3688), .DIN2(n3689), .DIN3(n3690), .DIN4(
        n3691) );
  nnd2s1 U5140 ( .Q(n3691), .DIN1(n3453), .DIN2(n3692) );
  nnd2s1 U5141 ( .Q(n3690), .DIN1(n3465), .DIN2(n3693) );
  nnd2s1 U5142 ( .Q(n3689), .DIN1(WX9566), .DIN2(n3517) );
  nnd2s1 U5143 ( .Q(n3688), .DIN1(CRC_OUT_2_16), .DIN2(n3549) );
  nnd4s1 U5144 ( .Q(WX9723), .DIN1(n3694), .DIN2(n3695), .DIN3(n3696), .DIN4(
        n3697) );
  nnd2s1 U5145 ( .Q(n3697), .DIN1(n3453), .DIN2(n3698) );
  nnd2s1 U5146 ( .Q(n3696), .DIN1(n3465), .DIN2(n3699) );
  nnd2s1 U5147 ( .Q(n3695), .DIN1(WX9564), .DIN2(n3517) );
  nnd2s1 U5148 ( .Q(n3694), .DIN1(CRC_OUT_2_17), .DIN2(n3549) );
  nnd4s1 U5149 ( .Q(WX9721), .DIN1(n3700), .DIN2(n3701), .DIN3(n3702), .DIN4(
        n3703) );
  nnd2s1 U5150 ( .Q(n3703), .DIN1(n3453), .DIN2(n3704) );
  nnd2s1 U5151 ( .Q(n3702), .DIN1(n3465), .DIN2(n3705) );
  nnd2s1 U5152 ( .Q(n3701), .DIN1(WX9562), .DIN2(n3517) );
  nnd2s1 U5153 ( .Q(n3700), .DIN1(CRC_OUT_2_18), .DIN2(n3549) );
  nnd4s1 U5154 ( .Q(WX9719), .DIN1(n3706), .DIN2(n3707), .DIN3(n3708), .DIN4(
        n3709) );
  nnd2s1 U5155 ( .Q(n3709), .DIN1(n3453), .DIN2(n3710) );
  nnd2s1 U5156 ( .Q(n3708), .DIN1(n3465), .DIN2(n3711) );
  nnd2s1 U5157 ( .Q(n3707), .DIN1(WX9560), .DIN2(n3517) );
  nnd2s1 U5158 ( .Q(n3706), .DIN1(CRC_OUT_2_19), .DIN2(n3549) );
  nnd4s1 U5159 ( .Q(WX9717), .DIN1(n3712), .DIN2(n3713), .DIN3(n3714), .DIN4(
        n3715) );
  nnd2s1 U5160 ( .Q(n3715), .DIN1(n3453), .DIN2(n3716) );
  nnd2s1 U5161 ( .Q(n3714), .DIN1(n3465), .DIN2(n3717) );
  nnd2s1 U5162 ( .Q(n3713), .DIN1(WX9558), .DIN2(n3517) );
  nnd2s1 U5163 ( .Q(n3712), .DIN1(CRC_OUT_2_20), .DIN2(n3549) );
  nnd4s1 U5164 ( .Q(WX9715), .DIN1(n3718), .DIN2(n3719), .DIN3(n3720), .DIN4(
        n3721) );
  nnd2s1 U5165 ( .Q(n3721), .DIN1(n3453), .DIN2(n3722) );
  nnd2s1 U5166 ( .Q(n3720), .DIN1(n3465), .DIN2(n3723) );
  nnd2s1 U5167 ( .Q(n3719), .DIN1(WX9556), .DIN2(n3517) );
  nnd2s1 U5168 ( .Q(n3718), .DIN1(CRC_OUT_2_21), .DIN2(n3549) );
  nnd4s1 U5169 ( .Q(WX9713), .DIN1(n3724), .DIN2(n3725), .DIN3(n3726), .DIN4(
        n3727) );
  nnd2s1 U5170 ( .Q(n3727), .DIN1(n3453), .DIN2(n3728) );
  nnd2s1 U5171 ( .Q(n3726), .DIN1(n3465), .DIN2(n3729) );
  nnd2s1 U5172 ( .Q(n3725), .DIN1(WX9554), .DIN2(n3517) );
  nnd2s1 U5173 ( .Q(n3724), .DIN1(CRC_OUT_2_22), .DIN2(n3549) );
  nnd4s1 U5174 ( .Q(WX9711), .DIN1(n3730), .DIN2(n3731), .DIN3(n3732), .DIN4(
        n3733) );
  nnd2s1 U5175 ( .Q(n3733), .DIN1(n3453), .DIN2(n3734) );
  nnd2s1 U5176 ( .Q(n3732), .DIN1(n3465), .DIN2(n3735) );
  nnd2s1 U5177 ( .Q(n3731), .DIN1(WX9552), .DIN2(n3517) );
  nnd2s1 U5178 ( .Q(n3730), .DIN1(CRC_OUT_2_23), .DIN2(n3549) );
  nnd4s1 U5179 ( .Q(WX9709), .DIN1(n3736), .DIN2(n3737), .DIN3(n3738), .DIN4(
        n3739) );
  nnd2s1 U5180 ( .Q(n3739), .DIN1(n3453), .DIN2(n3740) );
  nnd2s1 U5181 ( .Q(n3738), .DIN1(n3465), .DIN2(n3741) );
  nnd2s1 U5182 ( .Q(n3737), .DIN1(WX9550), .DIN2(n3516) );
  nnd2s1 U5183 ( .Q(n3736), .DIN1(CRC_OUT_2_24), .DIN2(n3548) );
  nnd4s1 U5184 ( .Q(WX9707), .DIN1(n3742), .DIN2(n3743), .DIN3(n3744), .DIN4(
        n3745) );
  nnd2s1 U5185 ( .Q(n3745), .DIN1(n3453), .DIN2(n3746) );
  nnd2s1 U5186 ( .Q(n3744), .DIN1(n3465), .DIN2(n3747) );
  nnd2s1 U5187 ( .Q(n3743), .DIN1(WX9548), .DIN2(n3516) );
  nnd2s1 U5188 ( .Q(n3742), .DIN1(CRC_OUT_2_25), .DIN2(n3548) );
  nnd4s1 U5189 ( .Q(WX9705), .DIN1(n3748), .DIN2(n3749), .DIN3(n3750), .DIN4(
        n3751) );
  nnd2s1 U5190 ( .Q(n3751), .DIN1(n3453), .DIN2(n3752) );
  nnd2s1 U5191 ( .Q(n3750), .DIN1(n3466), .DIN2(n3753) );
  nnd2s1 U5192 ( .Q(n3749), .DIN1(WX9546), .DIN2(n3516) );
  nnd2s1 U5193 ( .Q(n3748), .DIN1(CRC_OUT_2_26), .DIN2(n3548) );
  nnd4s1 U5194 ( .Q(WX9703), .DIN1(n3754), .DIN2(n3755), .DIN3(n3756), .DIN4(
        n3757) );
  nnd2s1 U5195 ( .Q(n3757), .DIN1(n3453), .DIN2(n3758) );
  nnd2s1 U5196 ( .Q(n3756), .DIN1(n3466), .DIN2(n3759) );
  nnd2s1 U5197 ( .Q(n3755), .DIN1(WX9544), .DIN2(n3516) );
  nnd2s1 U5198 ( .Q(n3754), .DIN1(CRC_OUT_2_27), .DIN2(n3548) );
  nnd4s1 U5199 ( .Q(WX9701), .DIN1(n3760), .DIN2(n3761), .DIN3(n3762), .DIN4(
        n3763) );
  nnd2s1 U5200 ( .Q(n3763), .DIN1(n3452), .DIN2(n3764) );
  nnd2s1 U5201 ( .Q(n3762), .DIN1(n3466), .DIN2(n3765) );
  nnd2s1 U5202 ( .Q(n3761), .DIN1(WX9542), .DIN2(n3516) );
  nnd2s1 U5203 ( .Q(n3760), .DIN1(CRC_OUT_2_28), .DIN2(n3548) );
  nnd4s1 U5204 ( .Q(WX9699), .DIN1(n3766), .DIN2(n3767), .DIN3(n3768), .DIN4(
        n3769) );
  nnd2s1 U5205 ( .Q(n3769), .DIN1(n3452), .DIN2(n3770) );
  nnd2s1 U5206 ( .Q(n3768), .DIN1(n3466), .DIN2(n3771) );
  nnd2s1 U5207 ( .Q(n3767), .DIN1(WX9540), .DIN2(n3516) );
  nnd2s1 U5208 ( .Q(n3766), .DIN1(CRC_OUT_2_29), .DIN2(n3548) );
  nnd4s1 U5209 ( .Q(WX9697), .DIN1(n3772), .DIN2(n3773), .DIN3(n3774), .DIN4(
        n3775) );
  nnd2s1 U5210 ( .Q(n3775), .DIN1(n3452), .DIN2(n3776) );
  nnd2s1 U5211 ( .Q(n3774), .DIN1(n3466), .DIN2(n3777) );
  nnd2s1 U5212 ( .Q(n3773), .DIN1(WX9538), .DIN2(n3516) );
  nnd2s1 U5213 ( .Q(n3772), .DIN1(CRC_OUT_2_30), .DIN2(n3548) );
  nnd4s1 U5214 ( .Q(WX9695), .DIN1(n3778), .DIN2(n3779), .DIN3(n3780), .DIN4(
        n3781) );
  nnd2s1 U5215 ( .Q(n3781), .DIN1(n3452), .DIN2(n3782) );
  nnd2s1 U5216 ( .Q(n3780), .DIN1(WX9536), .DIN2(n3516) );
  nnd2s1 U5217 ( .Q(n3779), .DIN1(n3466), .DIN2(n3783) );
  nnd2s1 U5218 ( .Q(n3778), .DIN1(CRC_OUT_2_31), .DIN2(n3548) );
  nor2s1 U5219 ( .Q(WX9597), .DIN1(WX9536), .DIN2(n3363) );
  and2s1 U5220 ( .Q(WX9595), .DIN1(RESET), .DIN2(WX9598) );
  and2s1 U5221 ( .Q(WX9593), .DIN1(RESET), .DIN2(WX9596) );
  and2s1 U5222 ( .Q(WX9591), .DIN1(RESET), .DIN2(WX9594) );
  and2s1 U5223 ( .Q(WX9589), .DIN1(RESET), .DIN2(WX9592) );
  and2s1 U5224 ( .Q(WX9587), .DIN1(RESET), .DIN2(WX9590) );
  and2s1 U5225 ( .Q(WX9585), .DIN1(RESET), .DIN2(WX9588) );
  and2s1 U5226 ( .Q(WX9583), .DIN1(RESET), .DIN2(WX9586) );
  and2s1 U5227 ( .Q(WX9581), .DIN1(RESET), .DIN2(WX9584) );
  and2s1 U5228 ( .Q(WX9579), .DIN1(RESET), .DIN2(WX9582) );
  and2s1 U5229 ( .Q(WX9577), .DIN1(RESET), .DIN2(WX9580) );
  and2s1 U5230 ( .Q(WX9575), .DIN1(RESET), .DIN2(WX9578) );
  and2s1 U5231 ( .Q(WX9573), .DIN1(RESET), .DIN2(WX9576) );
  and2s1 U5232 ( .Q(WX9571), .DIN1(RESET), .DIN2(WX9574) );
  and2s1 U5233 ( .Q(WX9569), .DIN1(RESET), .DIN2(WX9572) );
  and2s1 U5234 ( .Q(WX9567), .DIN1(RESET), .DIN2(WX9570) );
  and2s1 U5235 ( .Q(WX9565), .DIN1(RESET), .DIN2(WX9568) );
  and2s1 U5236 ( .Q(WX9563), .DIN1(RESET), .DIN2(WX9566) );
  and2s1 U5237 ( .Q(WX9561), .DIN1(RESET), .DIN2(WX9564) );
  and2s1 U5238 ( .Q(WX9559), .DIN1(RESET), .DIN2(WX9562) );
  and2s1 U5239 ( .Q(WX9557), .DIN1(RESET), .DIN2(WX9560) );
  and2s1 U5240 ( .Q(WX9555), .DIN1(RESET), .DIN2(WX9558) );
  and2s1 U5241 ( .Q(WX9553), .DIN1(RESET), .DIN2(WX9556) );
  and2s1 U5242 ( .Q(WX9551), .DIN1(RESET), .DIN2(WX9554) );
  and2s1 U5243 ( .Q(WX9549), .DIN1(RESET), .DIN2(WX9552) );
  and2s1 U5244 ( .Q(WX9547), .DIN1(RESET), .DIN2(WX9550) );
  and2s1 U5245 ( .Q(WX9545), .DIN1(RESET), .DIN2(WX9548) );
  and2s1 U5246 ( .Q(WX9543), .DIN1(RESET), .DIN2(WX9546) );
  and2s1 U5247 ( .Q(WX9541), .DIN1(RESET), .DIN2(WX9544) );
  and2s1 U5248 ( .Q(WX9539), .DIN1(RESET), .DIN2(WX9542) );
  and2s1 U5249 ( .Q(WX9537), .DIN1(RESET), .DIN2(WX9540) );
  and2s1 U5250 ( .Q(WX9535), .DIN1(RESET), .DIN2(WX9538) );
  nor2s1 U5251 ( .Q(WX9084), .DIN1(n3380), .DIN2(n3784) );
  xor2s1 U5252 ( .Q(n3784), .DIN1(WX8595), .DIN2(CRC_OUT_3_30) );
  nor2s1 U5253 ( .Q(WX9082), .DIN1(n3380), .DIN2(n3785) );
  xor2s1 U5254 ( .Q(n3785), .DIN1(WX8597), .DIN2(CRC_OUT_3_29) );
  nor2s1 U5255 ( .Q(WX9080), .DIN1(n3380), .DIN2(n3786) );
  xor2s1 U5256 ( .Q(n3786), .DIN1(WX8599), .DIN2(CRC_OUT_3_28) );
  nor2s1 U5257 ( .Q(WX9078), .DIN1(n3380), .DIN2(n3787) );
  xor2s1 U5258 ( .Q(n3787), .DIN1(WX8601), .DIN2(CRC_OUT_3_27) );
  nor2s1 U5259 ( .Q(WX9076), .DIN1(n3380), .DIN2(n3788) );
  xor2s1 U5260 ( .Q(n3788), .DIN1(WX8603), .DIN2(CRC_OUT_3_26) );
  nor2s1 U5261 ( .Q(WX9074), .DIN1(n3380), .DIN2(n3789) );
  xor2s1 U5262 ( .Q(n3789), .DIN1(WX8605), .DIN2(CRC_OUT_3_25) );
  nor2s1 U5263 ( .Q(WX9072), .DIN1(n3380), .DIN2(n3790) );
  xor2s1 U5264 ( .Q(n3790), .DIN1(WX8607), .DIN2(CRC_OUT_3_24) );
  nor2s1 U5265 ( .Q(WX9070), .DIN1(n3380), .DIN2(n3791) );
  xor2s1 U5266 ( .Q(n3791), .DIN1(WX8609), .DIN2(CRC_OUT_3_23) );
  nor2s1 U5267 ( .Q(WX9068), .DIN1(n3381), .DIN2(n3792) );
  xor2s1 U5268 ( .Q(n3792), .DIN1(WX8611), .DIN2(CRC_OUT_3_22) );
  nor2s1 U5269 ( .Q(WX9066), .DIN1(n3381), .DIN2(n3793) );
  xor2s1 U5270 ( .Q(n3793), .DIN1(WX8613), .DIN2(CRC_OUT_3_21) );
  nor2s1 U5271 ( .Q(WX9064), .DIN1(n3381), .DIN2(n3794) );
  xor2s1 U5272 ( .Q(n3794), .DIN1(WX8615), .DIN2(CRC_OUT_3_20) );
  nor2s1 U5273 ( .Q(WX9062), .DIN1(n3381), .DIN2(n3795) );
  xor2s1 U5274 ( .Q(n3795), .DIN1(WX8617), .DIN2(CRC_OUT_3_19) );
  nor2s1 U5275 ( .Q(WX9060), .DIN1(n3381), .DIN2(n3796) );
  xor2s1 U5276 ( .Q(n3796), .DIN1(WX8619), .DIN2(CRC_OUT_3_18) );
  nor2s1 U5277 ( .Q(WX9058), .DIN1(n3381), .DIN2(n3797) );
  xor2s1 U5278 ( .Q(n3797), .DIN1(WX8621), .DIN2(CRC_OUT_3_17) );
  nor2s1 U5279 ( .Q(WX9056), .DIN1(n3381), .DIN2(n3798) );
  xor2s1 U5280 ( .Q(n3798), .DIN1(WX8623), .DIN2(CRC_OUT_3_16) );
  nor2s1 U5281 ( .Q(WX9054), .DIN1(n3381), .DIN2(n3799) );
  xor2s1 U5282 ( .Q(n3799), .DIN1(CRC_OUT_3_15), .DIN2(n3800) );
  xor2s1 U5283 ( .Q(n3800), .DIN1(WX8625), .DIN2(CRC_OUT_3_31) );
  nor2s1 U5284 ( .Q(WX9052), .DIN1(n3381), .DIN2(n3801) );
  xor2s1 U5285 ( .Q(n3801), .DIN1(WX8627), .DIN2(CRC_OUT_3_14) );
  nor2s1 U5286 ( .Q(WX9050), .DIN1(n3381), .DIN2(n3802) );
  xor2s1 U5287 ( .Q(n3802), .DIN1(WX8629), .DIN2(CRC_OUT_3_13) );
  nor2s1 U5288 ( .Q(WX9048), .DIN1(n3382), .DIN2(n3803) );
  xor2s1 U5289 ( .Q(n3803), .DIN1(WX8631), .DIN2(CRC_OUT_3_12) );
  nor2s1 U5290 ( .Q(WX9046), .DIN1(n3382), .DIN2(n3804) );
  xor2s1 U5291 ( .Q(n3804), .DIN1(WX8633), .DIN2(CRC_OUT_3_11) );
  nor2s1 U5292 ( .Q(WX9044), .DIN1(n3382), .DIN2(n3805) );
  xor2s1 U5293 ( .Q(n3805), .DIN1(CRC_OUT_3_10), .DIN2(n3806) );
  xor2s1 U5294 ( .Q(n3806), .DIN1(WX8635), .DIN2(CRC_OUT_3_31) );
  nor2s1 U5295 ( .Q(WX9042), .DIN1(n3382), .DIN2(n3807) );
  xor2s1 U5296 ( .Q(n3807), .DIN1(WX8637), .DIN2(CRC_OUT_3_9) );
  nor2s1 U5297 ( .Q(WX9040), .DIN1(n3382), .DIN2(n3808) );
  xor2s1 U5298 ( .Q(n3808), .DIN1(WX8639), .DIN2(CRC_OUT_3_8) );
  nor2s1 U5299 ( .Q(WX9038), .DIN1(n3382), .DIN2(n3809) );
  xor2s1 U5300 ( .Q(n3809), .DIN1(WX8641), .DIN2(CRC_OUT_3_7) );
  nor2s1 U5301 ( .Q(WX9036), .DIN1(n3382), .DIN2(n3810) );
  xor2s1 U5302 ( .Q(n3810), .DIN1(WX8643), .DIN2(CRC_OUT_3_6) );
  nor2s1 U5303 ( .Q(WX9034), .DIN1(n3382), .DIN2(n3811) );
  xor2s1 U5304 ( .Q(n3811), .DIN1(WX8645), .DIN2(CRC_OUT_3_5) );
  nor2s1 U5305 ( .Q(WX9032), .DIN1(n3382), .DIN2(n3812) );
  xor2s1 U5306 ( .Q(n3812), .DIN1(WX8647), .DIN2(CRC_OUT_3_4) );
  nor2s1 U5307 ( .Q(WX9030), .DIN1(n3382), .DIN2(n3813) );
  xor2s1 U5308 ( .Q(n3813), .DIN1(CRC_OUT_3_3), .DIN2(n3814) );
  xor2s1 U5309 ( .Q(n3814), .DIN1(WX8649), .DIN2(CRC_OUT_3_31) );
  nor2s1 U5310 ( .Q(WX9028), .DIN1(n3383), .DIN2(n3815) );
  xor2s1 U5311 ( .Q(n3815), .DIN1(WX8651), .DIN2(CRC_OUT_3_2) );
  nor2s1 U5312 ( .Q(WX9026), .DIN1(n3383), .DIN2(n3816) );
  xor2s1 U5313 ( .Q(n3816), .DIN1(WX8653), .DIN2(CRC_OUT_3_1) );
  nor2s1 U5314 ( .Q(WX9024), .DIN1(n3383), .DIN2(n3817) );
  xor2s1 U5315 ( .Q(n3817), .DIN1(WX8655), .DIN2(CRC_OUT_3_0) );
  nor2s1 U5316 ( .Q(WX9022), .DIN1(n3383), .DIN2(n3818) );
  xor2s1 U5317 ( .Q(n3818), .DIN1(WX8657), .DIN2(CRC_OUT_3_31) );
  and2s1 U5318 ( .Q(WX898), .DIN1(RESET), .DIN2(WX835) );
  and2s1 U5319 ( .Q(WX896), .DIN1(RESET), .DIN2(WX833) );
  and2s1 U5320 ( .Q(WX894), .DIN1(RESET), .DIN2(WX831) );
  and2s1 U5321 ( .Q(WX892), .DIN1(RESET), .DIN2(WX829) );
  and2s1 U5322 ( .Q(WX890), .DIN1(RESET), .DIN2(WX827) );
  and2s1 U5323 ( .Q(WX888), .DIN1(RESET), .DIN2(WX825) );
  and2s1 U5324 ( .Q(WX886), .DIN1(RESET), .DIN2(WX823) );
  and2s1 U5325 ( .Q(WX884), .DIN1(RESET), .DIN2(WX821) );
  and2s1 U5326 ( .Q(WX882), .DIN1(RESET), .DIN2(WX819) );
  and2s1 U5327 ( .Q(WX880), .DIN1(RESET), .DIN2(WX817) );
  and2s1 U5328 ( .Q(WX878), .DIN1(RESET), .DIN2(WX815) );
  and2s1 U5329 ( .Q(WX876), .DIN1(RESET), .DIN2(WX813) );
  and2s1 U5330 ( .Q(WX874), .DIN1(RESET), .DIN2(WX811) );
  and2s1 U5331 ( .Q(WX872), .DIN1(RESET), .DIN2(WX809) );
  and2s1 U5332 ( .Q(WX870), .DIN1(RESET), .DIN2(WX807) );
  and2s1 U5333 ( .Q(WX868), .DIN1(RESET), .DIN2(WX805) );
  and2s1 U5334 ( .Q(WX866), .DIN1(RESET), .DIN2(WX803) );
  and2s1 U5335 ( .Q(WX8656), .DIN1(RESET), .DIN2(WX8593) );
  and2s1 U5336 ( .Q(WX8654), .DIN1(RESET), .DIN2(WX8591) );
  and2s1 U5337 ( .Q(WX8652), .DIN1(RESET), .DIN2(WX8589) );
  and2s1 U5338 ( .Q(WX8650), .DIN1(RESET), .DIN2(WX8587) );
  and2s1 U5339 ( .Q(WX8648), .DIN1(RESET), .DIN2(WX8585) );
  and2s1 U5340 ( .Q(WX8646), .DIN1(RESET), .DIN2(WX8583) );
  and2s1 U5341 ( .Q(WX8644), .DIN1(RESET), .DIN2(WX8581) );
  and2s1 U5342 ( .Q(WX8642), .DIN1(RESET), .DIN2(WX8579) );
  and2s1 U5343 ( .Q(WX8640), .DIN1(RESET), .DIN2(WX8577) );
  and2s1 U5344 ( .Q(WX864), .DIN1(RESET), .DIN2(WX801) );
  and2s1 U5345 ( .Q(WX8638), .DIN1(RESET), .DIN2(WX8575) );
  and2s1 U5346 ( .Q(WX8636), .DIN1(RESET), .DIN2(WX8573) );
  and2s1 U5347 ( .Q(WX8634), .DIN1(RESET), .DIN2(WX8571) );
  and2s1 U5348 ( .Q(WX8632), .DIN1(RESET), .DIN2(WX8569) );
  and2s1 U5349 ( .Q(WX8630), .DIN1(RESET), .DIN2(WX8567) );
  and2s1 U5350 ( .Q(WX8628), .DIN1(RESET), .DIN2(WX8565) );
  and2s1 U5351 ( .Q(WX8626), .DIN1(RESET), .DIN2(WX8563) );
  and2s1 U5352 ( .Q(WX8624), .DIN1(RESET), .DIN2(WX8561) );
  and2s1 U5353 ( .Q(WX8622), .DIN1(RESET), .DIN2(WX8559) );
  and2s1 U5354 ( .Q(WX8620), .DIN1(RESET), .DIN2(WX8557) );
  and2s1 U5355 ( .Q(WX862), .DIN1(RESET), .DIN2(WX799) );
  and2s1 U5356 ( .Q(WX8618), .DIN1(RESET), .DIN2(WX8555) );
  and2s1 U5357 ( .Q(WX8616), .DIN1(RESET), .DIN2(WX8553) );
  and2s1 U5358 ( .Q(WX8614), .DIN1(RESET), .DIN2(WX8551) );
  and2s1 U5359 ( .Q(WX8612), .DIN1(RESET), .DIN2(WX8549) );
  and2s1 U5360 ( .Q(WX8610), .DIN1(RESET), .DIN2(WX8547) );
  and2s1 U5361 ( .Q(WX8608), .DIN1(RESET), .DIN2(WX8545) );
  and2s1 U5362 ( .Q(WX8606), .DIN1(RESET), .DIN2(WX8543) );
  and2s1 U5363 ( .Q(WX8604), .DIN1(RESET), .DIN2(WX8541) );
  and2s1 U5364 ( .Q(WX8602), .DIN1(RESET), .DIN2(WX8539) );
  and2s1 U5365 ( .Q(WX8600), .DIN1(RESET), .DIN2(WX8537) );
  and2s1 U5366 ( .Q(WX860), .DIN1(RESET), .DIN2(WX797) );
  and2s1 U5367 ( .Q(WX8598), .DIN1(RESET), .DIN2(WX8535) );
  and2s1 U5368 ( .Q(WX8596), .DIN1(RESET), .DIN2(WX8533) );
  and2s1 U5369 ( .Q(WX8594), .DIN1(RESET), .DIN2(WX8531) );
  and2s1 U5370 ( .Q(WX8592), .DIN1(RESET), .DIN2(WX8529) );
  and2s1 U5371 ( .Q(WX8590), .DIN1(RESET), .DIN2(WX8527) );
  and2s1 U5372 ( .Q(WX8588), .DIN1(RESET), .DIN2(WX8525) );
  and2s1 U5373 ( .Q(WX8586), .DIN1(RESET), .DIN2(WX8523) );
  and2s1 U5374 ( .Q(WX8584), .DIN1(RESET), .DIN2(WX8521) );
  and2s1 U5375 ( .Q(WX8582), .DIN1(RESET), .DIN2(WX8519) );
  and2s1 U5376 ( .Q(WX8580), .DIN1(RESET), .DIN2(WX8517) );
  and2s1 U5377 ( .Q(WX858), .DIN1(RESET), .DIN2(WX795) );
  and2s1 U5378 ( .Q(WX8578), .DIN1(RESET), .DIN2(WX8515) );
  and2s1 U5379 ( .Q(WX8576), .DIN1(RESET), .DIN2(WX8513) );
  and2s1 U5380 ( .Q(WX8574), .DIN1(RESET), .DIN2(WX8511) );
  and2s1 U5381 ( .Q(WX8572), .DIN1(RESET), .DIN2(WX8509) );
  and2s1 U5382 ( .Q(WX8570), .DIN1(RESET), .DIN2(WX8507) );
  and2s1 U5383 ( .Q(WX8568), .DIN1(RESET), .DIN2(WX8505) );
  and2s1 U5384 ( .Q(WX8566), .DIN1(RESET), .DIN2(WX8503) );
  and2s1 U5385 ( .Q(WX8564), .DIN1(RESET), .DIN2(WX8501) );
  and2s1 U5386 ( .Q(WX8562), .DIN1(RESET), .DIN2(WX8499) );
  nor2s1 U5387 ( .Q(WX8560), .DIN1(n3383), .DIN2(n2965) );
  and2s1 U5388 ( .Q(WX856), .DIN1(RESET), .DIN2(WX793) );
  nor2s1 U5389 ( .Q(WX8558), .DIN1(n3383), .DIN2(n2966) );
  nor2s1 U5390 ( .Q(WX8556), .DIN1(n3383), .DIN2(n2967) );
  nor2s1 U5391 ( .Q(WX8554), .DIN1(n3383), .DIN2(n2968) );
  nor2s1 U5392 ( .Q(WX8552), .DIN1(n3383), .DIN2(n2969) );
  nor2s1 U5393 ( .Q(WX8550), .DIN1(n3384), .DIN2(n2970) );
  nor2s1 U5394 ( .Q(WX8548), .DIN1(n3384), .DIN2(n2971) );
  nor2s1 U5395 ( .Q(WX8546), .DIN1(n3384), .DIN2(n2972) );
  nor2s1 U5396 ( .Q(WX8544), .DIN1(n3384), .DIN2(n2973) );
  nor2s1 U5397 ( .Q(WX8542), .DIN1(n3384), .DIN2(n2974) );
  nor2s1 U5398 ( .Q(WX8540), .DIN1(n3384), .DIN2(n2975) );
  and2s1 U5399 ( .Q(WX854), .DIN1(RESET), .DIN2(WX791) );
  nor2s1 U5400 ( .Q(WX8538), .DIN1(n3384), .DIN2(n2976) );
  nor2s1 U5401 ( .Q(WX8536), .DIN1(n3384), .DIN2(n2977) );
  nor2s1 U5402 ( .Q(WX8534), .DIN1(n3384), .DIN2(n2978) );
  nor2s1 U5403 ( .Q(WX8532), .DIN1(n3384), .DIN2(n2979) );
  nor2s1 U5404 ( .Q(WX8530), .DIN1(n3385), .DIN2(n2980) );
  nor2s1 U5405 ( .Q(WX8528), .DIN1(n3385), .DIN2(n3125) );
  nor2s1 U5406 ( .Q(WX8526), .DIN1(n3385), .DIN2(n3126) );
  nor2s1 U5407 ( .Q(WX8524), .DIN1(n3385), .DIN2(n3127) );
  nor2s1 U5408 ( .Q(WX8522), .DIN1(n3385), .DIN2(n3128) );
  nor2s1 U5409 ( .Q(WX8520), .DIN1(n3385), .DIN2(n3129) );
  and2s1 U5410 ( .Q(WX852), .DIN1(RESET), .DIN2(WX789) );
  nor2s1 U5411 ( .Q(WX8518), .DIN1(n3385), .DIN2(n3130) );
  nor2s1 U5412 ( .Q(WX8516), .DIN1(n3385), .DIN2(n3131) );
  nor2s1 U5413 ( .Q(WX8514), .DIN1(n3385), .DIN2(n3132) );
  nor2s1 U5414 ( .Q(WX8512), .DIN1(n3385), .DIN2(n3133) );
  nor2s1 U5415 ( .Q(WX8510), .DIN1(n3386), .DIN2(n3134) );
  nor2s1 U5416 ( .Q(WX8508), .DIN1(n3386), .DIN2(n3135) );
  nor2s1 U5417 ( .Q(WX8506), .DIN1(n3386), .DIN2(n3136) );
  nor2s1 U5418 ( .Q(WX8504), .DIN1(n3386), .DIN2(n3137) );
  nor2s1 U5419 ( .Q(WX8502), .DIN1(n3386), .DIN2(n3138) );
  nor2s1 U5420 ( .Q(WX8500), .DIN1(n3386), .DIN2(n3139) );
  and2s1 U5421 ( .Q(WX850), .DIN1(RESET), .DIN2(WX787) );
  nor2s1 U5422 ( .Q(WX8498), .DIN1(n3386), .DIN2(n3140) );
  and2s1 U5423 ( .Q(WX8496), .DIN1(RESET), .DIN2(WX8433) );
  and2s1 U5424 ( .Q(WX8494), .DIN1(RESET), .DIN2(WX8431) );
  and2s1 U5425 ( .Q(WX8492), .DIN1(RESET), .DIN2(WX8429) );
  and2s1 U5426 ( .Q(WX8490), .DIN1(RESET), .DIN2(WX8427) );
  and2s1 U5427 ( .Q(WX8488), .DIN1(RESET), .DIN2(WX8425) );
  and2s1 U5428 ( .Q(WX8486), .DIN1(RESET), .DIN2(WX8423) );
  and2s1 U5429 ( .Q(WX8484), .DIN1(RESET), .DIN2(WX8421) );
  and2s1 U5430 ( .Q(WX8482), .DIN1(RESET), .DIN2(WX8419) );
  and2s1 U5431 ( .Q(WX8480), .DIN1(RESET), .DIN2(WX8417) );
  and2s1 U5432 ( .Q(WX848), .DIN1(RESET), .DIN2(WX785) );
  and2s1 U5433 ( .Q(WX8478), .DIN1(RESET), .DIN2(WX8415) );
  and2s1 U5434 ( .Q(WX8476), .DIN1(RESET), .DIN2(WX8413) );
  and2s1 U5435 ( .Q(WX8474), .DIN1(RESET), .DIN2(WX8411) );
  and2s1 U5436 ( .Q(WX8472), .DIN1(RESET), .DIN2(WX8409) );
  and2s1 U5437 ( .Q(WX8470), .DIN1(RESET), .DIN2(WX8407) );
  and2s1 U5438 ( .Q(WX8468), .DIN1(RESET), .DIN2(WX8405) );
  and2s1 U5439 ( .Q(WX8466), .DIN1(RESET), .DIN2(WX8403) );
  nnd4s1 U5440 ( .Q(WX8464), .DIN1(n3819), .DIN2(n3820), .DIN3(n3821), .DIN4(
        n3822) );
  nnd2s1 U5441 ( .Q(n3822), .DIN1(n3466), .DIN2(n3593) );
  xor2s1 U5442 ( .Q(n3593), .DIN1(n3823), .DIN2(n3824) );
  xor2s1 U5443 ( .Q(n3824), .DIN1(WX9822), .DIN2(n3109) );
  xor2s1 U5444 ( .Q(n3823), .DIN1(n3205), .DIN2(WX9886) );
  nnd2s1 U5445 ( .Q(n3821), .DIN1(n3452), .DIN2(n3825) );
  nnd2s1 U5446 ( .Q(n3820), .DIN1(WX8305), .DIN2(n3516) );
  nnd2s1 U5447 ( .Q(n3819), .DIN1(CRC_OUT_3_0), .DIN2(n3548) );
  nnd4s1 U5448 ( .Q(WX8462), .DIN1(n3826), .DIN2(n3827), .DIN3(n3828), .DIN4(
        n3829) );
  nnd2s1 U5449 ( .Q(n3829), .DIN1(n3466), .DIN2(n3602) );
  xor2s1 U5450 ( .Q(n3602), .DIN1(n3830), .DIN2(n3831) );
  xor2s1 U5451 ( .Q(n3831), .DIN1(WX9820), .DIN2(n3110) );
  xor2s1 U5452 ( .Q(n3830), .DIN1(n3206), .DIN2(WX9884) );
  nnd2s1 U5453 ( .Q(n3828), .DIN1(n3452), .DIN2(n3832) );
  nnd2s1 U5454 ( .Q(n3827), .DIN1(WX8303), .DIN2(n3516) );
  nnd2s1 U5455 ( .Q(n3826), .DIN1(CRC_OUT_3_1), .DIN2(n3548) );
  nnd4s1 U5456 ( .Q(WX8460), .DIN1(n3833), .DIN2(n3834), .DIN3(n3835), .DIN4(
        n3836) );
  nnd2s1 U5457 ( .Q(n3836), .DIN1(n3466), .DIN2(n3608) );
  xor2s1 U5458 ( .Q(n3608), .DIN1(n3837), .DIN2(n3838) );
  xor2s1 U5459 ( .Q(n3838), .DIN1(WX9818), .DIN2(n3111) );
  xor2s1 U5460 ( .Q(n3837), .DIN1(n3207), .DIN2(WX9882) );
  nnd2s1 U5461 ( .Q(n3835), .DIN1(n3452), .DIN2(n3839) );
  nnd2s1 U5462 ( .Q(n3834), .DIN1(WX8301), .DIN2(n3516) );
  nnd2s1 U5463 ( .Q(n3833), .DIN1(CRC_OUT_3_2), .DIN2(n3548) );
  and2s1 U5464 ( .Q(WX846), .DIN1(RESET), .DIN2(WX783) );
  nnd4s1 U5465 ( .Q(WX8458), .DIN1(n3840), .DIN2(n3841), .DIN3(n3842), .DIN4(
        n3843) );
  nnd2s1 U5466 ( .Q(n3843), .DIN1(n3466), .DIN2(n3614) );
  xor2s1 U5467 ( .Q(n3614), .DIN1(n3844), .DIN2(n3845) );
  xor2s1 U5468 ( .Q(n3845), .DIN1(WX9816), .DIN2(n3112) );
  xor2s1 U5469 ( .Q(n3844), .DIN1(n3208), .DIN2(WX9880) );
  nnd2s1 U5470 ( .Q(n3842), .DIN1(n3452), .DIN2(n3846) );
  nnd2s1 U5471 ( .Q(n3841), .DIN1(WX8299), .DIN2(n3516) );
  nnd2s1 U5472 ( .Q(n3840), .DIN1(CRC_OUT_3_3), .DIN2(n3548) );
  nnd4s1 U5473 ( .Q(WX8456), .DIN1(n3847), .DIN2(n3848), .DIN3(n3849), .DIN4(
        n3850) );
  nnd2s1 U5474 ( .Q(n3850), .DIN1(n3466), .DIN2(n3620) );
  xor2s1 U5475 ( .Q(n3620), .DIN1(n3851), .DIN2(n3852) );
  xor2s1 U5476 ( .Q(n3852), .DIN1(WX9814), .DIN2(n3113) );
  xor2s1 U5477 ( .Q(n3851), .DIN1(n3209), .DIN2(WX9878) );
  nnd2s1 U5478 ( .Q(n3849), .DIN1(n3452), .DIN2(n3853) );
  nnd2s1 U5479 ( .Q(n3848), .DIN1(WX8297), .DIN2(n3515) );
  nnd2s1 U5480 ( .Q(n3847), .DIN1(CRC_OUT_3_4), .DIN2(n3547) );
  nnd4s1 U5481 ( .Q(WX8454), .DIN1(n3854), .DIN2(n3855), .DIN3(n3856), .DIN4(
        n3857) );
  nnd2s1 U5482 ( .Q(n3857), .DIN1(n3466), .DIN2(n3626) );
  xor2s1 U5483 ( .Q(n3626), .DIN1(n3858), .DIN2(n3859) );
  xor2s1 U5484 ( .Q(n3859), .DIN1(WX9812), .DIN2(n3114) );
  xor2s1 U5485 ( .Q(n3858), .DIN1(n3210), .DIN2(WX9876) );
  nnd2s1 U5486 ( .Q(n3856), .DIN1(n3452), .DIN2(n3860) );
  nnd2s1 U5487 ( .Q(n3855), .DIN1(WX8295), .DIN2(n3515) );
  nnd2s1 U5488 ( .Q(n3854), .DIN1(CRC_OUT_3_5), .DIN2(n3547) );
  nnd4s1 U5489 ( .Q(WX8452), .DIN1(n3861), .DIN2(n3862), .DIN3(n3863), .DIN4(
        n3864) );
  nnd2s1 U5490 ( .Q(n3864), .DIN1(n3466), .DIN2(n3632) );
  xor2s1 U5491 ( .Q(n3632), .DIN1(n3865), .DIN2(n3866) );
  xor2s1 U5492 ( .Q(n3866), .DIN1(WX9810), .DIN2(n3115) );
  xor2s1 U5493 ( .Q(n3865), .DIN1(n3211), .DIN2(WX9874) );
  nnd2s1 U5494 ( .Q(n3863), .DIN1(n3452), .DIN2(n3867) );
  nnd2s1 U5495 ( .Q(n3862), .DIN1(WX8293), .DIN2(n3515) );
  nnd2s1 U5496 ( .Q(n3861), .DIN1(CRC_OUT_3_6), .DIN2(n3547) );
  nnd4s1 U5497 ( .Q(WX8450), .DIN1(n3868), .DIN2(n3869), .DIN3(n3870), .DIN4(
        n3871) );
  nnd2s1 U5498 ( .Q(n3871), .DIN1(n3467), .DIN2(n3638) );
  xor2s1 U5499 ( .Q(n3638), .DIN1(n3872), .DIN2(n3873) );
  xor2s1 U5500 ( .Q(n3873), .DIN1(WX9808), .DIN2(n3116) );
  xor2s1 U5501 ( .Q(n3872), .DIN1(n3212), .DIN2(WX9872) );
  nnd2s1 U5502 ( .Q(n3870), .DIN1(n3452), .DIN2(n3874) );
  nnd2s1 U5503 ( .Q(n3869), .DIN1(WX8291), .DIN2(n3515) );
  nnd2s1 U5504 ( .Q(n3868), .DIN1(CRC_OUT_3_7), .DIN2(n3547) );
  nnd4s1 U5505 ( .Q(WX8448), .DIN1(n3875), .DIN2(n3876), .DIN3(n3877), .DIN4(
        n3878) );
  nnd2s1 U5506 ( .Q(n3878), .DIN1(n3467), .DIN2(n3644) );
  xor2s1 U5507 ( .Q(n3644), .DIN1(n3879), .DIN2(n3880) );
  xor2s1 U5508 ( .Q(n3880), .DIN1(WX9806), .DIN2(n3117) );
  xor2s1 U5509 ( .Q(n3879), .DIN1(n3213), .DIN2(WX9870) );
  nnd2s1 U5510 ( .Q(n3877), .DIN1(n3452), .DIN2(n3881) );
  nnd2s1 U5511 ( .Q(n3876), .DIN1(WX8289), .DIN2(n3515) );
  nnd2s1 U5512 ( .Q(n3875), .DIN1(CRC_OUT_3_8), .DIN2(n3547) );
  nnd4s1 U5513 ( .Q(WX8446), .DIN1(n3882), .DIN2(n3883), .DIN3(n3884), .DIN4(
        n3885) );
  nnd2s1 U5514 ( .Q(n3885), .DIN1(n3467), .DIN2(n3650) );
  xor2s1 U5515 ( .Q(n3650), .DIN1(n3886), .DIN2(n3887) );
  xor2s1 U5516 ( .Q(n3887), .DIN1(WX9804), .DIN2(n3118) );
  xor2s1 U5517 ( .Q(n3886), .DIN1(n3214), .DIN2(WX9868) );
  nnd2s1 U5518 ( .Q(n3884), .DIN1(n3451), .DIN2(n3888) );
  nnd2s1 U5519 ( .Q(n3883), .DIN1(WX8287), .DIN2(n3515) );
  nnd2s1 U5520 ( .Q(n3882), .DIN1(CRC_OUT_3_9), .DIN2(n3547) );
  nnd4s1 U5521 ( .Q(WX8444), .DIN1(n3889), .DIN2(n3890), .DIN3(n3891), .DIN4(
        n3892) );
  nnd2s1 U5522 ( .Q(n3892), .DIN1(n3467), .DIN2(n3656) );
  xor2s1 U5523 ( .Q(n3656), .DIN1(n3893), .DIN2(n3894) );
  xor2s1 U5524 ( .Q(n3894), .DIN1(WX9802), .DIN2(n3119) );
  xor2s1 U5525 ( .Q(n3893), .DIN1(n3215), .DIN2(WX9866) );
  nnd2s1 U5526 ( .Q(n3891), .DIN1(n3451), .DIN2(n3895) );
  nnd2s1 U5527 ( .Q(n3890), .DIN1(WX8285), .DIN2(n3515) );
  nnd2s1 U5528 ( .Q(n3889), .DIN1(CRC_OUT_3_10), .DIN2(n3547) );
  nnd4s1 U5529 ( .Q(WX8442), .DIN1(n3896), .DIN2(n3897), .DIN3(n3898), .DIN4(
        n3899) );
  nnd2s1 U5530 ( .Q(n3899), .DIN1(n3467), .DIN2(n3662) );
  xor2s1 U5531 ( .Q(n3662), .DIN1(n3900), .DIN2(n3901) );
  xor2s1 U5532 ( .Q(n3901), .DIN1(WX9800), .DIN2(n3120) );
  xor2s1 U5533 ( .Q(n3900), .DIN1(n3216), .DIN2(WX9864) );
  nnd2s1 U5534 ( .Q(n3898), .DIN1(n3451), .DIN2(n3902) );
  nnd2s1 U5535 ( .Q(n3897), .DIN1(WX8283), .DIN2(n3515) );
  nnd2s1 U5536 ( .Q(n3896), .DIN1(CRC_OUT_3_11), .DIN2(n3547) );
  nnd4s1 U5537 ( .Q(WX8440), .DIN1(n3903), .DIN2(n3904), .DIN3(n3905), .DIN4(
        n3906) );
  nnd2s1 U5538 ( .Q(n3906), .DIN1(n3467), .DIN2(n3668) );
  xor2s1 U5539 ( .Q(n3668), .DIN1(n3907), .DIN2(n3908) );
  xor2s1 U5540 ( .Q(n3908), .DIN1(WX9798), .DIN2(n3121) );
  xor2s1 U5541 ( .Q(n3907), .DIN1(n3217), .DIN2(WX9862) );
  nnd2s1 U5542 ( .Q(n3905), .DIN1(n3451), .DIN2(n3909) );
  nnd2s1 U5543 ( .Q(n3904), .DIN1(WX8281), .DIN2(n3515) );
  nnd2s1 U5544 ( .Q(n3903), .DIN1(CRC_OUT_3_12), .DIN2(n3547) );
  and2s1 U5545 ( .Q(WX844), .DIN1(RESET), .DIN2(WX781) );
  nnd4s1 U5546 ( .Q(WX8438), .DIN1(n3910), .DIN2(n3911), .DIN3(n3912), .DIN4(
        n3913) );
  nnd2s1 U5547 ( .Q(n3913), .DIN1(n3467), .DIN2(n3674) );
  xor2s1 U5548 ( .Q(n3674), .DIN1(n3914), .DIN2(n3915) );
  xor2s1 U5549 ( .Q(n3915), .DIN1(WX9796), .DIN2(n3122) );
  xor2s1 U5550 ( .Q(n3914), .DIN1(n3218), .DIN2(WX9860) );
  nnd2s1 U5551 ( .Q(n3912), .DIN1(n3451), .DIN2(n3916) );
  nnd2s1 U5552 ( .Q(n3911), .DIN1(WX8279), .DIN2(n3515) );
  nnd2s1 U5553 ( .Q(n3910), .DIN1(CRC_OUT_3_13), .DIN2(n3547) );
  nnd4s1 U5554 ( .Q(WX8436), .DIN1(n3917), .DIN2(n3918), .DIN3(n3919), .DIN4(
        n3920) );
  nnd2s1 U5555 ( .Q(n3920), .DIN1(n3467), .DIN2(n3680) );
  xor2s1 U5556 ( .Q(n3680), .DIN1(n3921), .DIN2(n3922) );
  xor2s1 U5557 ( .Q(n3922), .DIN1(WX9794), .DIN2(n3123) );
  xor2s1 U5558 ( .Q(n3921), .DIN1(n3219), .DIN2(WX9858) );
  nnd2s1 U5559 ( .Q(n3919), .DIN1(n3451), .DIN2(n3923) );
  nnd2s1 U5560 ( .Q(n3918), .DIN1(WX8277), .DIN2(n3515) );
  nnd2s1 U5561 ( .Q(n3917), .DIN1(CRC_OUT_3_14), .DIN2(n3547) );
  nnd4s1 U5562 ( .Q(WX8434), .DIN1(n3924), .DIN2(n3925), .DIN3(n3926), .DIN4(
        n3927) );
  nnd2s1 U5563 ( .Q(n3927), .DIN1(n3467), .DIN2(n3686) );
  xor2s1 U5564 ( .Q(n3686), .DIN1(n3928), .DIN2(n3929) );
  xor2s1 U5565 ( .Q(n3929), .DIN1(WX9792), .DIN2(n3124) );
  xor2s1 U5566 ( .Q(n3928), .DIN1(n3220), .DIN2(WX9856) );
  nnd2s1 U5567 ( .Q(n3926), .DIN1(n3451), .DIN2(n3930) );
  nnd2s1 U5568 ( .Q(n3925), .DIN1(WX8275), .DIN2(n3515) );
  nnd2s1 U5569 ( .Q(n3924), .DIN1(CRC_OUT_3_15), .DIN2(n3547) );
  nnd4s1 U5570 ( .Q(WX8432), .DIN1(n3931), .DIN2(n3932), .DIN3(n3933), .DIN4(
        n3934) );
  nnd2s1 U5571 ( .Q(n3934), .DIN1(n3467), .DIN2(n3692) );
  xor2s1 U5572 ( .Q(n3692), .DIN1(n3935), .DIN2(n3936) );
  xor2s1 U5573 ( .Q(n3936), .DIN1(n3569), .DIN2(WX9726) );
  xor2s1 U5574 ( .Q(n3935), .DIN1(n2949), .DIN2(n3938) );
  xor2s1 U5575 ( .Q(n3938), .DIN1(WX9918), .DIN2(WX9854) );
  nnd2s1 U5576 ( .Q(n3933), .DIN1(n3451), .DIN2(n3939) );
  nnd2s1 U5577 ( .Q(n3932), .DIN1(WX8273), .DIN2(n3514) );
  nnd2s1 U5578 ( .Q(n3931), .DIN1(CRC_OUT_3_16), .DIN2(n3546) );
  nnd4s1 U5579 ( .Q(WX8430), .DIN1(n3940), .DIN2(n3941), .DIN3(n3942), .DIN4(
        n3943) );
  nnd2s1 U5580 ( .Q(n3943), .DIN1(n3467), .DIN2(n3698) );
  xor2s1 U5581 ( .Q(n3698), .DIN1(n3944), .DIN2(n3360) );
  xor2s1 U5582 ( .Q(n3945), .DIN1(n3559), .DIN2(WX9724) );
  xor2s1 U5583 ( .Q(n3944), .DIN1(n2950), .DIN2(n3946) );
  xor2s1 U5584 ( .Q(n3946), .DIN1(WX9916), .DIN2(WX9852) );
  nnd2s1 U5585 ( .Q(n3942), .DIN1(n3451), .DIN2(n3947) );
  nnd2s1 U5586 ( .Q(n3941), .DIN1(WX8271), .DIN2(n3514) );
  nnd2s1 U5587 ( .Q(n3940), .DIN1(CRC_OUT_3_17), .DIN2(n3546) );
  nnd4s1 U5588 ( .Q(WX8428), .DIN1(n3948), .DIN2(n3949), .DIN3(n3950), .DIN4(
        n3951) );
  nnd2s1 U5589 ( .Q(n3951), .DIN1(n3467), .DIN2(n3704) );
  xor2s1 U5590 ( .Q(n3704), .DIN1(n3952), .DIN2(n3356) );
  xor2s1 U5591 ( .Q(n3953), .DIN1(n3559), .DIN2(WX9722) );
  xor2s1 U5592 ( .Q(n3952), .DIN1(n2951), .DIN2(n3954) );
  xor2s1 U5593 ( .Q(n3954), .DIN1(WX9914), .DIN2(WX9850) );
  nnd2s1 U5594 ( .Q(n3950), .DIN1(n3451), .DIN2(n3955) );
  nnd2s1 U5595 ( .Q(n3949), .DIN1(WX8269), .DIN2(n3514) );
  nnd2s1 U5596 ( .Q(n3948), .DIN1(CRC_OUT_3_18), .DIN2(n3546) );
  nnd4s1 U5597 ( .Q(WX8426), .DIN1(n3956), .DIN2(n3957), .DIN3(n3958), .DIN4(
        n3959) );
  nnd2s1 U5598 ( .Q(n3959), .DIN1(n3467), .DIN2(n3710) );
  xor2s1 U5599 ( .Q(n3710), .DIN1(n3960), .DIN2(n3352) );
  xor2s1 U5600 ( .Q(n3961), .DIN1(n3559), .DIN2(WX9720) );
  xor2s1 U5601 ( .Q(n3960), .DIN1(n2952), .DIN2(n3962) );
  xor2s1 U5602 ( .Q(n3962), .DIN1(WX9912), .DIN2(WX9848) );
  nnd2s1 U5603 ( .Q(n3958), .DIN1(n3451), .DIN2(n3963) );
  nnd2s1 U5604 ( .Q(n3957), .DIN1(WX8267), .DIN2(n3514) );
  nnd2s1 U5605 ( .Q(n3956), .DIN1(CRC_OUT_3_19), .DIN2(n3546) );
  nnd4s1 U5606 ( .Q(WX8424), .DIN1(n3964), .DIN2(n3965), .DIN3(n3966), .DIN4(
        n3967) );
  nnd2s1 U5607 ( .Q(n3967), .DIN1(n3468), .DIN2(n3716) );
  xor2s1 U5608 ( .Q(n3716), .DIN1(n3968), .DIN2(n3348) );
  xor2s1 U5609 ( .Q(n3969), .DIN1(n3559), .DIN2(WX9718) );
  xor2s1 U5610 ( .Q(n3968), .DIN1(n2953), .DIN2(n3970) );
  xor2s1 U5611 ( .Q(n3970), .DIN1(WX9910), .DIN2(WX9846) );
  nnd2s1 U5612 ( .Q(n3966), .DIN1(n3451), .DIN2(n3971) );
  nnd2s1 U5613 ( .Q(n3965), .DIN1(WX8265), .DIN2(n3514) );
  nnd2s1 U5614 ( .Q(n3964), .DIN1(CRC_OUT_3_20), .DIN2(n3546) );
  nnd4s1 U5615 ( .Q(WX8422), .DIN1(n3972), .DIN2(n3973), .DIN3(n3974), .DIN4(
        n3975) );
  nnd2s1 U5616 ( .Q(n3975), .DIN1(n3468), .DIN2(n3722) );
  xor2s1 U5617 ( .Q(n3722), .DIN1(n3976), .DIN2(n3344) );
  xor2s1 U5618 ( .Q(n3977), .DIN1(n3559), .DIN2(WX9716) );
  xor2s1 U5619 ( .Q(n3976), .DIN1(n2954), .DIN2(n3978) );
  xor2s1 U5620 ( .Q(n3978), .DIN1(WX9908), .DIN2(WX9844) );
  nnd2s1 U5621 ( .Q(n3974), .DIN1(n3451), .DIN2(n3979) );
  nnd2s1 U5622 ( .Q(n3973), .DIN1(WX8263), .DIN2(n3514) );
  nnd2s1 U5623 ( .Q(n3972), .DIN1(CRC_OUT_3_21), .DIN2(n3546) );
  nnd4s1 U5624 ( .Q(WX8420), .DIN1(n3980), .DIN2(n3981), .DIN3(n3982), .DIN4(
        n3983) );
  nnd2s1 U5625 ( .Q(n3983), .DIN1(n3468), .DIN2(n3728) );
  xor2s1 U5626 ( .Q(n3728), .DIN1(n3984), .DIN2(n3340) );
  xor2s1 U5627 ( .Q(n3985), .DIN1(n3559), .DIN2(WX9714) );
  xor2s1 U5628 ( .Q(n3984), .DIN1(n2955), .DIN2(n3986) );
  xor2s1 U5629 ( .Q(n3986), .DIN1(WX9906), .DIN2(WX9842) );
  nnd2s1 U5630 ( .Q(n3982), .DIN1(n3450), .DIN2(n3987) );
  nnd2s1 U5631 ( .Q(n3981), .DIN1(WX8261), .DIN2(n3514) );
  nnd2s1 U5632 ( .Q(n3980), .DIN1(CRC_OUT_3_22), .DIN2(n3546) );
  and2s1 U5633 ( .Q(WX842), .DIN1(RESET), .DIN2(WX779) );
  nnd4s1 U5634 ( .Q(WX8418), .DIN1(n3988), .DIN2(n3989), .DIN3(n3990), .DIN4(
        n3991) );
  nnd2s1 U5635 ( .Q(n3991), .DIN1(n3468), .DIN2(n3734) );
  xor2s1 U5636 ( .Q(n3734), .DIN1(n3992), .DIN2(n3336) );
  xor2s1 U5637 ( .Q(n3993), .DIN1(n3560), .DIN2(WX9712) );
  xor2s1 U5638 ( .Q(n3992), .DIN1(n2956), .DIN2(n3994) );
  xor2s1 U5639 ( .Q(n3994), .DIN1(WX9904), .DIN2(WX9840) );
  nnd2s1 U5640 ( .Q(n3990), .DIN1(n3450), .DIN2(n3995) );
  nnd2s1 U5641 ( .Q(n3989), .DIN1(WX8259), .DIN2(n3514) );
  nnd2s1 U5642 ( .Q(n3988), .DIN1(CRC_OUT_3_23), .DIN2(n3546) );
  nnd4s1 U5643 ( .Q(WX8416), .DIN1(n3996), .DIN2(n3997), .DIN3(n3998), .DIN4(
        n3999) );
  nnd2s1 U5644 ( .Q(n3999), .DIN1(n3468), .DIN2(n3740) );
  xor2s1 U5645 ( .Q(n3740), .DIN1(n4000), .DIN2(n3334) );
  xor2s1 U5646 ( .Q(n4001), .DIN1(n3560), .DIN2(WX9710) );
  xor2s1 U5647 ( .Q(n4000), .DIN1(n2957), .DIN2(n4002) );
  xor2s1 U5648 ( .Q(n4002), .DIN1(WX9902), .DIN2(WX9838) );
  nnd2s1 U5649 ( .Q(n3998), .DIN1(n3450), .DIN2(n4003) );
  nnd2s1 U5650 ( .Q(n3997), .DIN1(WX8257), .DIN2(n3514) );
  nnd2s1 U5651 ( .Q(n3996), .DIN1(CRC_OUT_3_24), .DIN2(n3546) );
  nnd4s1 U5652 ( .Q(WX8414), .DIN1(n4004), .DIN2(n4005), .DIN3(n4006), .DIN4(
        n4007) );
  nnd2s1 U5653 ( .Q(n4007), .DIN1(n3468), .DIN2(n3746) );
  xor2s1 U5654 ( .Q(n3746), .DIN1(n4008), .DIN2(n3338) );
  xor2s1 U5655 ( .Q(n4009), .DIN1(n3560), .DIN2(WX9708) );
  xor2s1 U5656 ( .Q(n4008), .DIN1(n2958), .DIN2(n4010) );
  xor2s1 U5657 ( .Q(n4010), .DIN1(WX9900), .DIN2(WX9836) );
  nnd2s1 U5658 ( .Q(n4006), .DIN1(n3450), .DIN2(n4011) );
  nnd2s1 U5659 ( .Q(n4005), .DIN1(WX8255), .DIN2(n3514) );
  nnd2s1 U5660 ( .Q(n4004), .DIN1(CRC_OUT_3_25), .DIN2(n3546) );
  nnd4s1 U5661 ( .Q(WX8412), .DIN1(n4012), .DIN2(n4013), .DIN3(n4014), .DIN4(
        n4015) );
  nnd2s1 U5662 ( .Q(n4015), .DIN1(n3468), .DIN2(n3752) );
  xor2s1 U5663 ( .Q(n3752), .DIN1(n4016), .DIN2(n3342) );
  xor2s1 U5664 ( .Q(n4017), .DIN1(n3560), .DIN2(WX9706) );
  xor2s1 U5665 ( .Q(n4016), .DIN1(n2959), .DIN2(n4018) );
  xor2s1 U5666 ( .Q(n4018), .DIN1(WX9898), .DIN2(WX9834) );
  nnd2s1 U5667 ( .Q(n4014), .DIN1(n3450), .DIN2(n4019) );
  nnd2s1 U5668 ( .Q(n4013), .DIN1(WX8253), .DIN2(n3514) );
  nnd2s1 U5669 ( .Q(n4012), .DIN1(CRC_OUT_3_26), .DIN2(n3546) );
  nnd4s1 U5670 ( .Q(WX8410), .DIN1(n4020), .DIN2(n4021), .DIN3(n4022), .DIN4(
        n4023) );
  nnd2s1 U5671 ( .Q(n4023), .DIN1(n3468), .DIN2(n3758) );
  xor2s1 U5672 ( .Q(n3758), .DIN1(n4024), .DIN2(n3346) );
  xor2s1 U5673 ( .Q(n4025), .DIN1(n3560), .DIN2(WX9704) );
  xor2s1 U5674 ( .Q(n4024), .DIN1(n2960), .DIN2(n4026) );
  xor2s1 U5675 ( .Q(n4026), .DIN1(WX9896), .DIN2(WX9832) );
  nnd2s1 U5676 ( .Q(n4022), .DIN1(n3450), .DIN2(n4027) );
  nnd2s1 U5677 ( .Q(n4021), .DIN1(WX8251), .DIN2(n3514) );
  nnd2s1 U5678 ( .Q(n4020), .DIN1(CRC_OUT_3_27), .DIN2(n3546) );
  nnd4s1 U5679 ( .Q(WX8408), .DIN1(n4028), .DIN2(n4029), .DIN3(n4030), .DIN4(
        n4031) );
  nnd2s1 U5680 ( .Q(n4031), .DIN1(n3468), .DIN2(n3764) );
  xor2s1 U5681 ( .Q(n3764), .DIN1(n4032), .DIN2(n3350) );
  xor2s1 U5682 ( .Q(n4033), .DIN1(n3560), .DIN2(WX9702) );
  xor2s1 U5683 ( .Q(n4032), .DIN1(n2961), .DIN2(n4034) );
  xor2s1 U5684 ( .Q(n4034), .DIN1(WX9894), .DIN2(WX9830) );
  nnd2s1 U5685 ( .Q(n4030), .DIN1(n3450), .DIN2(n4035) );
  nnd2s1 U5686 ( .Q(n4029), .DIN1(WX8249), .DIN2(n3513) );
  nnd2s1 U5687 ( .Q(n4028), .DIN1(CRC_OUT_3_28), .DIN2(n3545) );
  nnd4s1 U5688 ( .Q(WX8406), .DIN1(n4036), .DIN2(n4037), .DIN3(n4038), .DIN4(
        n4039) );
  nnd2s1 U5689 ( .Q(n4039), .DIN1(n3468), .DIN2(n3770) );
  xor2s1 U5690 ( .Q(n3770), .DIN1(n4040), .DIN2(n3354) );
  xor2s1 U5691 ( .Q(n4041), .DIN1(n3560), .DIN2(WX9700) );
  xor2s1 U5692 ( .Q(n4040), .DIN1(n2962), .DIN2(n4042) );
  xor2s1 U5693 ( .Q(n4042), .DIN1(WX9892), .DIN2(WX9828) );
  nnd2s1 U5694 ( .Q(n4038), .DIN1(n3450), .DIN2(n4043) );
  nnd2s1 U5695 ( .Q(n4037), .DIN1(WX8247), .DIN2(n3513) );
  nnd2s1 U5696 ( .Q(n4036), .DIN1(CRC_OUT_3_29), .DIN2(n3545) );
  nnd4s1 U5697 ( .Q(WX8404), .DIN1(n4044), .DIN2(n4045), .DIN3(n4046), .DIN4(
        n4047) );
  nnd2s1 U5698 ( .Q(n4047), .DIN1(n3468), .DIN2(n3776) );
  xor2s1 U5699 ( .Q(n3776), .DIN1(n4048), .DIN2(n4049) );
  xor2s1 U5700 ( .Q(n4049), .DIN1(n3561), .DIN2(WX9698) );
  xor2s1 U5701 ( .Q(n4048), .DIN1(n2963), .DIN2(n4050) );
  xor2s1 U5702 ( .Q(n4050), .DIN1(WX9890), .DIN2(WX9826) );
  nnd2s1 U5703 ( .Q(n4046), .DIN1(n3450), .DIN2(n4051) );
  nnd2s1 U5704 ( .Q(n4045), .DIN1(WX8245), .DIN2(n3513) );
  nnd2s1 U5705 ( .Q(n4044), .DIN1(CRC_OUT_3_30), .DIN2(n3545) );
  nnd4s1 U5706 ( .Q(WX8402), .DIN1(n4052), .DIN2(n4053), .DIN3(n4054), .DIN4(
        n4055) );
  nnd2s1 U5707 ( .Q(n4055), .DIN1(n3468), .DIN2(n3782) );
  xor2s1 U5708 ( .Q(n3782), .DIN1(n4056), .DIN2(n4057) );
  xor2s1 U5709 ( .Q(n4057), .DIN1(n3561), .DIN2(WX9696) );
  xor2s1 U5710 ( .Q(n4056), .DIN1(n2964), .DIN2(n4058) );
  xor2s1 U5711 ( .Q(n4058), .DIN1(WX9888), .DIN2(WX9824) );
  nnd2s1 U5712 ( .Q(n4054), .DIN1(n3450), .DIN2(n4059) );
  nnd2s1 U5713 ( .Q(n4053), .DIN1(WX8243), .DIN2(n3513) );
  nnd2s1 U5714 ( .Q(n4052), .DIN1(CRC_OUT_3_31), .DIN2(n3545) );
  and2s1 U5715 ( .Q(WX840), .DIN1(RESET), .DIN2(WX777) );
  and2s1 U5716 ( .Q(WX838), .DIN1(RESET), .DIN2(WX775) );
  and2s1 U5717 ( .Q(WX836), .DIN1(RESET), .DIN2(WX773) );
  and2s1 U5718 ( .Q(WX834), .DIN1(RESET), .DIN2(WX771) );
  and2s1 U5719 ( .Q(WX832), .DIN1(RESET), .DIN2(WX769) );
  nor2s1 U5720 ( .Q(WX8304), .DIN1(WX8243), .DIN2(n3363) );
  and2s1 U5721 ( .Q(WX8302), .DIN1(RESET), .DIN2(WX8305) );
  and2s1 U5722 ( .Q(WX8300), .DIN1(RESET), .DIN2(WX8303) );
  and2s1 U5723 ( .Q(WX830), .DIN1(RESET), .DIN2(WX767) );
  and2s1 U5724 ( .Q(WX8298), .DIN1(RESET), .DIN2(WX8301) );
  and2s1 U5725 ( .Q(WX8296), .DIN1(RESET), .DIN2(WX8299) );
  and2s1 U5726 ( .Q(WX8294), .DIN1(RESET), .DIN2(WX8297) );
  and2s1 U5727 ( .Q(WX8292), .DIN1(RESET), .DIN2(WX8295) );
  and2s1 U5728 ( .Q(WX8290), .DIN1(RESET), .DIN2(WX8293) );
  and2s1 U5729 ( .Q(WX8288), .DIN1(RESET), .DIN2(WX8291) );
  and2s1 U5730 ( .Q(WX8286), .DIN1(RESET), .DIN2(WX8289) );
  and2s1 U5731 ( .Q(WX8284), .DIN1(RESET), .DIN2(WX8287) );
  and2s1 U5732 ( .Q(WX8282), .DIN1(RESET), .DIN2(WX8285) );
  and2s1 U5733 ( .Q(WX8280), .DIN1(RESET), .DIN2(WX8283) );
  and2s1 U5734 ( .Q(WX828), .DIN1(RESET), .DIN2(WX765) );
  and2s1 U5735 ( .Q(WX8278), .DIN1(RESET), .DIN2(WX8281) );
  and2s1 U5736 ( .Q(WX8276), .DIN1(RESET), .DIN2(WX8279) );
  and2s1 U5737 ( .Q(WX8274), .DIN1(RESET), .DIN2(WX8277) );
  and2s1 U5738 ( .Q(WX8272), .DIN1(RESET), .DIN2(WX8275) );
  and2s1 U5739 ( .Q(WX8270), .DIN1(RESET), .DIN2(WX8273) );
  and2s1 U5740 ( .Q(WX8268), .DIN1(RESET), .DIN2(WX8271) );
  and2s1 U5741 ( .Q(WX8266), .DIN1(RESET), .DIN2(WX8269) );
  and2s1 U5742 ( .Q(WX8264), .DIN1(RESET), .DIN2(WX8267) );
  and2s1 U5743 ( .Q(WX8262), .DIN1(RESET), .DIN2(WX8265) );
  and2s1 U5744 ( .Q(WX8260), .DIN1(RESET), .DIN2(WX8263) );
  and2s1 U5745 ( .Q(WX826), .DIN1(RESET), .DIN2(WX763) );
  and2s1 U5746 ( .Q(WX8258), .DIN1(RESET), .DIN2(WX8261) );
  and2s1 U5747 ( .Q(WX8256), .DIN1(RESET), .DIN2(WX8259) );
  and2s1 U5748 ( .Q(WX8254), .DIN1(RESET), .DIN2(WX8257) );
  and2s1 U5749 ( .Q(WX8252), .DIN1(RESET), .DIN2(WX8255) );
  and2s1 U5750 ( .Q(WX8250), .DIN1(RESET), .DIN2(WX8253) );
  and2s1 U5751 ( .Q(WX8248), .DIN1(RESET), .DIN2(WX8251) );
  and2s1 U5752 ( .Q(WX8246), .DIN1(RESET), .DIN2(WX8249) );
  and2s1 U5753 ( .Q(WX8244), .DIN1(RESET), .DIN2(WX8247) );
  and2s1 U5754 ( .Q(WX8242), .DIN1(RESET), .DIN2(WX8245) );
  and2s1 U5755 ( .Q(WX824), .DIN1(RESET), .DIN2(WX761) );
  and2s1 U5756 ( .Q(WX822), .DIN1(RESET), .DIN2(WX759) );
  and2s1 U5757 ( .Q(WX820), .DIN1(RESET), .DIN2(WX757) );
  and2s1 U5758 ( .Q(WX818), .DIN1(RESET), .DIN2(WX755) );
  and2s1 U5759 ( .Q(WX816), .DIN1(RESET), .DIN2(WX753) );
  and2s1 U5760 ( .Q(WX814), .DIN1(RESET), .DIN2(WX751) );
  and2s1 U5761 ( .Q(WX812), .DIN1(RESET), .DIN2(WX749) );
  and2s1 U5762 ( .Q(WX810), .DIN1(RESET), .DIN2(WX747) );
  and2s1 U5763 ( .Q(WX808), .DIN1(RESET), .DIN2(WX745) );
  and2s1 U5764 ( .Q(WX806), .DIN1(RESET), .DIN2(WX743) );
  and2s1 U5765 ( .Q(WX804), .DIN1(RESET), .DIN2(WX741) );
  and2s1 U5766 ( .Q(WX802), .DIN1(RESET), .DIN2(WX739) );
  and2s1 U5767 ( .Q(WX800), .DIN1(RESET), .DIN2(WX737) );
  and2s1 U5768 ( .Q(WX798), .DIN1(RESET), .DIN2(WX735) );
  and2s1 U5769 ( .Q(WX796), .DIN1(RESET), .DIN2(WX733) );
  and2s1 U5770 ( .Q(WX794), .DIN1(RESET), .DIN2(WX731) );
  and2s1 U5771 ( .Q(WX792), .DIN1(RESET), .DIN2(WX729) );
  and2s1 U5772 ( .Q(WX790), .DIN1(RESET), .DIN2(WX727) );
  and2s1 U5773 ( .Q(WX788), .DIN1(RESET), .DIN2(WX725) );
  and2s1 U5774 ( .Q(WX786), .DIN1(RESET), .DIN2(WX723) );
  and2s1 U5775 ( .Q(WX784), .DIN1(RESET), .DIN2(WX721) );
  and2s1 U5776 ( .Q(WX782), .DIN1(RESET), .DIN2(WX719) );
  and2s1 U5777 ( .Q(WX780), .DIN1(RESET), .DIN2(WX717) );
  nor2s1 U5778 ( .Q(WX7791), .DIN1(n3386), .DIN2(n4060) );
  xor2s1 U5779 ( .Q(n4060), .DIN1(WX7302), .DIN2(CRC_OUT_4_30) );
  nor2s1 U5780 ( .Q(WX7789), .DIN1(n3386), .DIN2(n4061) );
  xor2s1 U5781 ( .Q(n4061), .DIN1(WX7304), .DIN2(CRC_OUT_4_29) );
  nor2s1 U5782 ( .Q(WX7787), .DIN1(n3386), .DIN2(n4062) );
  xor2s1 U5783 ( .Q(n4062), .DIN1(WX7306), .DIN2(CRC_OUT_4_28) );
  nor2s1 U5784 ( .Q(WX7785), .DIN1(n3387), .DIN2(n4063) );
  xor2s1 U5785 ( .Q(n4063), .DIN1(WX7308), .DIN2(CRC_OUT_4_27) );
  nor2s1 U5786 ( .Q(WX7783), .DIN1(n3387), .DIN2(n4064) );
  xor2s1 U5787 ( .Q(n4064), .DIN1(WX7310), .DIN2(CRC_OUT_4_26) );
  nor2s1 U5788 ( .Q(WX7781), .DIN1(n3387), .DIN2(n4065) );
  xor2s1 U5789 ( .Q(n4065), .DIN1(WX7312), .DIN2(CRC_OUT_4_25) );
  and2s1 U5790 ( .Q(WX778), .DIN1(RESET), .DIN2(WX715) );
  nor2s1 U5791 ( .Q(WX7779), .DIN1(n3387), .DIN2(n4066) );
  xor2s1 U5792 ( .Q(n4066), .DIN1(WX7314), .DIN2(CRC_OUT_4_24) );
  nor2s1 U5793 ( .Q(WX7777), .DIN1(n3387), .DIN2(n4067) );
  xor2s1 U5794 ( .Q(n4067), .DIN1(WX7316), .DIN2(CRC_OUT_4_23) );
  nor2s1 U5795 ( .Q(WX7775), .DIN1(n3387), .DIN2(n4068) );
  xor2s1 U5796 ( .Q(n4068), .DIN1(WX7318), .DIN2(CRC_OUT_4_22) );
  nor2s1 U5797 ( .Q(WX7773), .DIN1(n3387), .DIN2(n4069) );
  xor2s1 U5798 ( .Q(n4069), .DIN1(WX7320), .DIN2(CRC_OUT_4_21) );
  nor2s1 U5799 ( .Q(WX7771), .DIN1(n3387), .DIN2(n4070) );
  xor2s1 U5800 ( .Q(n4070), .DIN1(WX7322), .DIN2(CRC_OUT_4_20) );
  nor2s1 U5801 ( .Q(WX7769), .DIN1(n3387), .DIN2(n4071) );
  xor2s1 U5802 ( .Q(n4071), .DIN1(WX7324), .DIN2(CRC_OUT_4_19) );
  nor2s1 U5803 ( .Q(WX7767), .DIN1(n3387), .DIN2(n4072) );
  xor2s1 U5804 ( .Q(n4072), .DIN1(WX7326), .DIN2(CRC_OUT_4_18) );
  nor2s1 U5805 ( .Q(WX7765), .DIN1(n3388), .DIN2(n4073) );
  xor2s1 U5806 ( .Q(n4073), .DIN1(WX7328), .DIN2(CRC_OUT_4_17) );
  nor2s1 U5807 ( .Q(WX7763), .DIN1(n3388), .DIN2(n4074) );
  xor2s1 U5808 ( .Q(n4074), .DIN1(WX7330), .DIN2(CRC_OUT_4_16) );
  nor2s1 U5809 ( .Q(WX7761), .DIN1(n3388), .DIN2(n4075) );
  xor2s1 U5810 ( .Q(n4075), .DIN1(CRC_OUT_4_15), .DIN2(n4076) );
  xor2s1 U5811 ( .Q(n4076), .DIN1(WX7332), .DIN2(CRC_OUT_4_31) );
  and2s1 U5812 ( .Q(WX776), .DIN1(RESET), .DIN2(WX713) );
  nor2s1 U5813 ( .Q(WX7759), .DIN1(n3388), .DIN2(n4077) );
  xor2s1 U5814 ( .Q(n4077), .DIN1(WX7334), .DIN2(CRC_OUT_4_14) );
  nor2s1 U5815 ( .Q(WX7757), .DIN1(n3388), .DIN2(n4078) );
  xor2s1 U5816 ( .Q(n4078), .DIN1(WX7336), .DIN2(CRC_OUT_4_13) );
  nor2s1 U5817 ( .Q(WX7755), .DIN1(n3388), .DIN2(n4079) );
  xor2s1 U5818 ( .Q(n4079), .DIN1(WX7338), .DIN2(CRC_OUT_4_12) );
  nor2s1 U5819 ( .Q(WX7753), .DIN1(n3388), .DIN2(n4080) );
  xor2s1 U5820 ( .Q(n4080), .DIN1(WX7340), .DIN2(CRC_OUT_4_11) );
  nor2s1 U5821 ( .Q(WX7751), .DIN1(n3388), .DIN2(n4081) );
  xor2s1 U5822 ( .Q(n4081), .DIN1(CRC_OUT_4_10), .DIN2(n4082) );
  xor2s1 U5823 ( .Q(n4082), .DIN1(WX7342), .DIN2(CRC_OUT_4_31) );
  nor2s1 U5824 ( .Q(WX7749), .DIN1(n3388), .DIN2(n4083) );
  xor2s1 U5825 ( .Q(n4083), .DIN1(WX7344), .DIN2(CRC_OUT_4_9) );
  nor2s1 U5826 ( .Q(WX7747), .DIN1(n3388), .DIN2(n4084) );
  xor2s1 U5827 ( .Q(n4084), .DIN1(WX7346), .DIN2(CRC_OUT_4_8) );
  nor2s1 U5828 ( .Q(WX7745), .DIN1(n3389), .DIN2(n4085) );
  xor2s1 U5829 ( .Q(n4085), .DIN1(WX7348), .DIN2(CRC_OUT_4_7) );
  nor2s1 U5830 ( .Q(WX7743), .DIN1(n3389), .DIN2(n4086) );
  xor2s1 U5831 ( .Q(n4086), .DIN1(WX7350), .DIN2(CRC_OUT_4_6) );
  nor2s1 U5832 ( .Q(WX7741), .DIN1(n3389), .DIN2(n4087) );
  xor2s1 U5833 ( .Q(n4087), .DIN1(WX7352), .DIN2(CRC_OUT_4_5) );
  and2s1 U5834 ( .Q(WX774), .DIN1(RESET), .DIN2(WX711) );
  nor2s1 U5835 ( .Q(WX7739), .DIN1(n3389), .DIN2(n4088) );
  xor2s1 U5836 ( .Q(n4088), .DIN1(WX7354), .DIN2(CRC_OUT_4_4) );
  nor2s1 U5837 ( .Q(WX7737), .DIN1(n3389), .DIN2(n4089) );
  xor2s1 U5838 ( .Q(n4089), .DIN1(CRC_OUT_4_3), .DIN2(n4090) );
  xor2s1 U5839 ( .Q(n4090), .DIN1(WX7356), .DIN2(CRC_OUT_4_31) );
  nor2s1 U5840 ( .Q(WX7735), .DIN1(n3389), .DIN2(n4091) );
  xor2s1 U5841 ( .Q(n4091), .DIN1(WX7358), .DIN2(CRC_OUT_4_2) );
  nor2s1 U5842 ( .Q(WX7733), .DIN1(n3389), .DIN2(n4092) );
  xor2s1 U5843 ( .Q(n4092), .DIN1(WX7360), .DIN2(CRC_OUT_4_1) );
  nor2s1 U5844 ( .Q(WX7731), .DIN1(n3389), .DIN2(n4093) );
  xor2s1 U5845 ( .Q(n4093), .DIN1(WX7362), .DIN2(CRC_OUT_4_0) );
  nor2s1 U5846 ( .Q(WX7729), .DIN1(n3389), .DIN2(n4094) );
  xor2s1 U5847 ( .Q(n4094), .DIN1(WX7364), .DIN2(CRC_OUT_4_31) );
  and2s1 U5848 ( .Q(WX772), .DIN1(RESET), .DIN2(WX709) );
  and2s1 U5849 ( .Q(WX770), .DIN1(RESET), .DIN2(WX707) );
  and2s1 U5850 ( .Q(WX768), .DIN1(RESET), .DIN2(WX705) );
  and2s1 U5851 ( .Q(WX766), .DIN1(RESET), .DIN2(WX703) );
  and2s1 U5852 ( .Q(WX764), .DIN1(RESET), .DIN2(WX701) );
  and2s1 U5853 ( .Q(WX762), .DIN1(RESET), .DIN2(WX699) );
  and2s1 U5854 ( .Q(WX760), .DIN1(RESET), .DIN2(WX697) );
  and2s1 U5855 ( .Q(WX758), .DIN1(RESET), .DIN2(WX695) );
  and2s1 U5856 ( .Q(WX756), .DIN1(RESET), .DIN2(WX693) );
  and2s1 U5857 ( .Q(WX754), .DIN1(RESET), .DIN2(WX691) );
  and2s1 U5858 ( .Q(WX752), .DIN1(RESET), .DIN2(WX689) );
  and2s1 U5859 ( .Q(WX750), .DIN1(RESET), .DIN2(WX687) );
  and2s1 U5860 ( .Q(WX748), .DIN1(RESET), .DIN2(WX685) );
  and2s1 U5861 ( .Q(WX746), .DIN1(RESET), .DIN2(WX683) );
  and2s1 U5862 ( .Q(WX744), .DIN1(RESET), .DIN2(WX681) );
  and2s1 U5863 ( .Q(WX742), .DIN1(RESET), .DIN2(WX679) );
  and2s1 U5864 ( .Q(WX740), .DIN1(RESET), .DIN2(WX677) );
  and2s1 U5865 ( .Q(WX738), .DIN1(RESET), .DIN2(WX675) );
  and2s1 U5866 ( .Q(WX7363), .DIN1(RESET), .DIN2(WX7300) );
  and2s1 U5867 ( .Q(WX7361), .DIN1(RESET), .DIN2(WX7298) );
  and2s1 U5868 ( .Q(WX736), .DIN1(RESET), .DIN2(WX673) );
  and2s1 U5869 ( .Q(WX7359), .DIN1(RESET), .DIN2(WX7296) );
  and2s1 U5870 ( .Q(WX7357), .DIN1(RESET), .DIN2(WX7294) );
  and2s1 U5871 ( .Q(WX7355), .DIN1(RESET), .DIN2(WX7292) );
  and2s1 U5872 ( .Q(WX7353), .DIN1(RESET), .DIN2(WX7290) );
  and2s1 U5873 ( .Q(WX7351), .DIN1(RESET), .DIN2(WX7288) );
  and2s1 U5874 ( .Q(WX7349), .DIN1(RESET), .DIN2(WX7286) );
  and2s1 U5875 ( .Q(WX7347), .DIN1(RESET), .DIN2(WX7284) );
  and2s1 U5876 ( .Q(WX7345), .DIN1(RESET), .DIN2(WX7282) );
  and2s1 U5877 ( .Q(WX7343), .DIN1(RESET), .DIN2(WX7280) );
  and2s1 U5878 ( .Q(WX7341), .DIN1(RESET), .DIN2(WX7278) );
  and2s1 U5879 ( .Q(WX734), .DIN1(RESET), .DIN2(WX671) );
  and2s1 U5880 ( .Q(WX7339), .DIN1(RESET), .DIN2(WX7276) );
  and2s1 U5881 ( .Q(WX7337), .DIN1(RESET), .DIN2(WX7274) );
  and2s1 U5882 ( .Q(WX7335), .DIN1(RESET), .DIN2(WX7272) );
  and2s1 U5883 ( .Q(WX7333), .DIN1(RESET), .DIN2(WX7270) );
  and2s1 U5884 ( .Q(WX7331), .DIN1(RESET), .DIN2(WX7268) );
  and2s1 U5885 ( .Q(WX7329), .DIN1(RESET), .DIN2(WX7266) );
  and2s1 U5886 ( .Q(WX7327), .DIN1(RESET), .DIN2(WX7264) );
  and2s1 U5887 ( .Q(WX7325), .DIN1(RESET), .DIN2(WX7262) );
  and2s1 U5888 ( .Q(WX7323), .DIN1(RESET), .DIN2(WX7260) );
  and2s1 U5889 ( .Q(WX7321), .DIN1(RESET), .DIN2(WX7258) );
  and2s1 U5890 ( .Q(WX732), .DIN1(RESET), .DIN2(WX669) );
  and2s1 U5891 ( .Q(WX7319), .DIN1(RESET), .DIN2(WX7256) );
  and2s1 U5892 ( .Q(WX7317), .DIN1(RESET), .DIN2(WX7254) );
  and2s1 U5893 ( .Q(WX7315), .DIN1(RESET), .DIN2(WX7252) );
  and2s1 U5894 ( .Q(WX7313), .DIN1(RESET), .DIN2(WX7250) );
  and2s1 U5895 ( .Q(WX7311), .DIN1(RESET), .DIN2(WX7248) );
  and2s1 U5896 ( .Q(WX7309), .DIN1(RESET), .DIN2(WX7246) );
  and2s1 U5897 ( .Q(WX7307), .DIN1(RESET), .DIN2(WX7244) );
  and2s1 U5898 ( .Q(WX7305), .DIN1(RESET), .DIN2(WX7242) );
  and2s1 U5899 ( .Q(WX7303), .DIN1(RESET), .DIN2(WX7240) );
  and2s1 U5900 ( .Q(WX7301), .DIN1(RESET), .DIN2(WX7238) );
  and2s1 U5901 ( .Q(WX730), .DIN1(RESET), .DIN2(WX667) );
  and2s1 U5902 ( .Q(WX7299), .DIN1(RESET), .DIN2(WX7236) );
  and2s1 U5903 ( .Q(WX7297), .DIN1(RESET), .DIN2(WX7234) );
  and2s1 U5904 ( .Q(WX7295), .DIN1(RESET), .DIN2(WX7232) );
  and2s1 U5905 ( .Q(WX7293), .DIN1(RESET), .DIN2(WX7230) );
  and2s1 U5906 ( .Q(WX7291), .DIN1(RESET), .DIN2(WX7228) );
  and2s1 U5907 ( .Q(WX7289), .DIN1(RESET), .DIN2(WX7226) );
  and2s1 U5908 ( .Q(WX7287), .DIN1(RESET), .DIN2(WX7224) );
  and2s1 U5909 ( .Q(WX7285), .DIN1(RESET), .DIN2(WX7222) );
  and2s1 U5910 ( .Q(WX7283), .DIN1(RESET), .DIN2(WX7220) );
  and2s1 U5911 ( .Q(WX7281), .DIN1(RESET), .DIN2(WX7218) );
  and2s1 U5912 ( .Q(WX728), .DIN1(RESET), .DIN2(WX665) );
  and2s1 U5913 ( .Q(WX7279), .DIN1(RESET), .DIN2(WX7216) );
  and2s1 U5914 ( .Q(WX7277), .DIN1(RESET), .DIN2(WX7214) );
  and2s1 U5915 ( .Q(WX7275), .DIN1(RESET), .DIN2(WX7212) );
  and2s1 U5916 ( .Q(WX7273), .DIN1(RESET), .DIN2(WX7210) );
  and2s1 U5917 ( .Q(WX7271), .DIN1(RESET), .DIN2(WX7208) );
  and2s1 U5918 ( .Q(WX7269), .DIN1(RESET), .DIN2(WX7206) );
  nor2s1 U5919 ( .Q(WX7267), .DIN1(n3389), .DIN2(n2981) );
  nor2s1 U5920 ( .Q(WX7265), .DIN1(n3390), .DIN2(n2982) );
  nor2s1 U5921 ( .Q(WX7263), .DIN1(n3390), .DIN2(n2983) );
  nor2s1 U5922 ( .Q(WX7261), .DIN1(n3390), .DIN2(n2984) );
  and2s1 U5923 ( .Q(WX726), .DIN1(RESET), .DIN2(WX663) );
  nor2s1 U5924 ( .Q(WX7259), .DIN1(n3390), .DIN2(n2985) );
  nor2s1 U5925 ( .Q(WX7257), .DIN1(n3390), .DIN2(n2986) );
  nor2s1 U5926 ( .Q(WX7255), .DIN1(n3390), .DIN2(n2987) );
  nor2s1 U5927 ( .Q(WX7253), .DIN1(n3390), .DIN2(n2988) );
  nor2s1 U5928 ( .Q(WX7251), .DIN1(n3390), .DIN2(n2989) );
  nor2s1 U5929 ( .Q(WX7249), .DIN1(n3370), .DIN2(n2990) );
  nor2s1 U5930 ( .Q(WX7247), .DIN1(n3363), .DIN2(n2991) );
  nor2s1 U5931 ( .Q(WX7245), .DIN1(n3364), .DIN2(n2992) );
  nor2s1 U5932 ( .Q(WX7243), .DIN1(n3364), .DIN2(n2993) );
  nor2s1 U5933 ( .Q(WX7241), .DIN1(n3364), .DIN2(n2994) );
  and2s1 U5934 ( .Q(WX724), .DIN1(RESET), .DIN2(WX661) );
  nor2s1 U5935 ( .Q(WX7239), .DIN1(n3364), .DIN2(n2995) );
  nor2s1 U5936 ( .Q(WX7237), .DIN1(n3365), .DIN2(n2996) );
  nor2s1 U5937 ( .Q(WX7235), .DIN1(n3364), .DIN2(n3141) );
  nor2s1 U5938 ( .Q(WX7233), .DIN1(n3364), .DIN2(n3142) );
  nor2s1 U5939 ( .Q(WX7231), .DIN1(n3364), .DIN2(n3143) );
  nor2s1 U5940 ( .Q(WX7229), .DIN1(n3364), .DIN2(n3144) );
  nor2s1 U5941 ( .Q(WX7227), .DIN1(n3366), .DIN2(n3145) );
  nor2s1 U5942 ( .Q(WX7225), .DIN1(n3364), .DIN2(n3146) );
  nor2s1 U5943 ( .Q(WX7223), .DIN1(n3365), .DIN2(n3147) );
  nor2s1 U5944 ( .Q(WX7221), .DIN1(n3364), .DIN2(n3148) );
  and2s1 U5945 ( .Q(WX722), .DIN1(RESET), .DIN2(WX659) );
  nor2s1 U5946 ( .Q(WX7219), .DIN1(n3365), .DIN2(n3149) );
  nor2s1 U5947 ( .Q(WX7217), .DIN1(n3365), .DIN2(n3150) );
  nor2s1 U5948 ( .Q(WX7215), .DIN1(n3365), .DIN2(n3151) );
  nor2s1 U5949 ( .Q(WX7213), .DIN1(n3365), .DIN2(n3152) );
  nor2s1 U5950 ( .Q(WX7211), .DIN1(n3365), .DIN2(n3153) );
  nor2s1 U5951 ( .Q(WX7209), .DIN1(n3365), .DIN2(n3154) );
  nor2s1 U5952 ( .Q(WX7207), .DIN1(n3365), .DIN2(n3155) );
  nor2s1 U5953 ( .Q(WX7205), .DIN1(n3366), .DIN2(n3156) );
  and2s1 U5954 ( .Q(WX7203), .DIN1(RESET), .DIN2(WX7140) );
  and2s1 U5955 ( .Q(WX7201), .DIN1(RESET), .DIN2(WX7138) );
  and2s1 U5956 ( .Q(WX720), .DIN1(RESET), .DIN2(WX657) );
  and2s1 U5957 ( .Q(WX7199), .DIN1(RESET), .DIN2(WX7136) );
  and2s1 U5958 ( .Q(WX7197), .DIN1(RESET), .DIN2(WX7134) );
  and2s1 U5959 ( .Q(WX7195), .DIN1(RESET), .DIN2(WX7132) );
  and2s1 U5960 ( .Q(WX7193), .DIN1(RESET), .DIN2(WX7130) );
  and2s1 U5961 ( .Q(WX7191), .DIN1(RESET), .DIN2(WX7128) );
  and2s1 U5962 ( .Q(WX7189), .DIN1(RESET), .DIN2(WX7126) );
  and2s1 U5963 ( .Q(WX7187), .DIN1(RESET), .DIN2(WX7124) );
  and2s1 U5964 ( .Q(WX7185), .DIN1(RESET), .DIN2(WX7122) );
  and2s1 U5965 ( .Q(WX7183), .DIN1(RESET), .DIN2(WX7120) );
  and2s1 U5966 ( .Q(WX7181), .DIN1(RESET), .DIN2(WX7118) );
  and2s1 U5967 ( .Q(WX718), .DIN1(RESET), .DIN2(WX655) );
  and2s1 U5968 ( .Q(WX7179), .DIN1(RESET), .DIN2(WX7116) );
  and2s1 U5969 ( .Q(WX7177), .DIN1(RESET), .DIN2(WX7114) );
  and2s1 U5970 ( .Q(WX7175), .DIN1(RESET), .DIN2(WX7112) );
  and2s1 U5971 ( .Q(WX7173), .DIN1(RESET), .DIN2(WX7110) );
  nnd4s1 U5972 ( .Q(WX7171), .DIN1(n4095), .DIN2(n4096), .DIN3(n4097), .DIN4(
        n4098) );
  nnd2s1 U5973 ( .Q(n4098), .DIN1(n3468), .DIN2(n3825) );
  xor2s1 U5974 ( .Q(n3825), .DIN1(n4099), .DIN2(n4100) );
  xor2s1 U5975 ( .Q(n4100), .DIN1(WX8529), .DIN2(n3125) );
  xor2s1 U5976 ( .Q(n4099), .DIN1(n3221), .DIN2(WX8593) );
  nnd2s1 U5977 ( .Q(n4097), .DIN1(n3450), .DIN2(n4101) );
  nnd2s1 U5978 ( .Q(n4096), .DIN1(WX7012), .DIN2(n3513) );
  nnd2s1 U5979 ( .Q(n4095), .DIN1(CRC_OUT_4_0), .DIN2(n3545) );
  nnd4s1 U5980 ( .Q(WX7169), .DIN1(n4102), .DIN2(n4103), .DIN3(n4104), .DIN4(
        n4105) );
  nnd2s1 U5981 ( .Q(n4105), .DIN1(n3469), .DIN2(n3832) );
  xor2s1 U5982 ( .Q(n3832), .DIN1(n4106), .DIN2(n4107) );
  xor2s1 U5983 ( .Q(n4107), .DIN1(WX8527), .DIN2(n3126) );
  xor2s1 U5984 ( .Q(n4106), .DIN1(n3222), .DIN2(WX8591) );
  nnd2s1 U5985 ( .Q(n4104), .DIN1(n3450), .DIN2(n4108) );
  nnd2s1 U5986 ( .Q(n4103), .DIN1(WX7010), .DIN2(n3513) );
  nnd2s1 U5987 ( .Q(n4102), .DIN1(CRC_OUT_4_1), .DIN2(n3545) );
  nnd4s1 U5988 ( .Q(WX7167), .DIN1(n4109), .DIN2(n4110), .DIN3(n4111), .DIN4(
        n4112) );
  nnd2s1 U5989 ( .Q(n4112), .DIN1(n3469), .DIN2(n3839) );
  xor2s1 U5990 ( .Q(n3839), .DIN1(n4113), .DIN2(n4114) );
  xor2s1 U5991 ( .Q(n4114), .DIN1(WX8525), .DIN2(n3127) );
  xor2s1 U5992 ( .Q(n4113), .DIN1(n3223), .DIN2(WX8589) );
  nnd2s1 U5993 ( .Q(n4111), .DIN1(n3450), .DIN2(n4115) );
  nnd2s1 U5994 ( .Q(n4110), .DIN1(WX7008), .DIN2(n3513) );
  nnd2s1 U5995 ( .Q(n4109), .DIN1(CRC_OUT_4_2), .DIN2(n3545) );
  nnd4s1 U5996 ( .Q(WX7165), .DIN1(n4116), .DIN2(n4117), .DIN3(n4118), .DIN4(
        n4119) );
  nnd2s1 U5997 ( .Q(n4119), .DIN1(n3469), .DIN2(n3846) );
  xor2s1 U5998 ( .Q(n3846), .DIN1(n4120), .DIN2(n4121) );
  xor2s1 U5999 ( .Q(n4121), .DIN1(WX8523), .DIN2(n3128) );
  xor2s1 U6000 ( .Q(n4120), .DIN1(n3224), .DIN2(WX8587) );
  nnd2s1 U6001 ( .Q(n4118), .DIN1(n3449), .DIN2(n4122) );
  nnd2s1 U6002 ( .Q(n4117), .DIN1(WX7006), .DIN2(n3513) );
  nnd2s1 U6003 ( .Q(n4116), .DIN1(CRC_OUT_4_3), .DIN2(n3545) );
  nnd4s1 U6004 ( .Q(WX7163), .DIN1(n4123), .DIN2(n4124), .DIN3(n4125), .DIN4(
        n4126) );
  nnd2s1 U6005 ( .Q(n4126), .DIN1(n3469), .DIN2(n3853) );
  xor2s1 U6006 ( .Q(n3853), .DIN1(n4127), .DIN2(n4128) );
  xor2s1 U6007 ( .Q(n4128), .DIN1(WX8521), .DIN2(n3129) );
  xor2s1 U6008 ( .Q(n4127), .DIN1(n3225), .DIN2(WX8585) );
  nnd2s1 U6009 ( .Q(n4125), .DIN1(n3449), .DIN2(n4129) );
  nnd2s1 U6010 ( .Q(n4124), .DIN1(WX7004), .DIN2(n3513) );
  nnd2s1 U6011 ( .Q(n4123), .DIN1(CRC_OUT_4_4), .DIN2(n3545) );
  nnd4s1 U6012 ( .Q(WX7161), .DIN1(n4130), .DIN2(n4131), .DIN3(n4132), .DIN4(
        n4133) );
  nnd2s1 U6013 ( .Q(n4133), .DIN1(n3469), .DIN2(n3860) );
  xor2s1 U6014 ( .Q(n3860), .DIN1(n4134), .DIN2(n4135) );
  xor2s1 U6015 ( .Q(n4135), .DIN1(WX8519), .DIN2(n3130) );
  xor2s1 U6016 ( .Q(n4134), .DIN1(n3226), .DIN2(WX8583) );
  nnd2s1 U6017 ( .Q(n4132), .DIN1(n3449), .DIN2(n4136) );
  nnd2s1 U6018 ( .Q(n4131), .DIN1(WX7002), .DIN2(n3513) );
  nnd2s1 U6019 ( .Q(n4130), .DIN1(CRC_OUT_4_5), .DIN2(n3545) );
  and2s1 U6020 ( .Q(WX716), .DIN1(RESET), .DIN2(WX653) );
  nnd4s1 U6021 ( .Q(WX7159), .DIN1(n4137), .DIN2(n4138), .DIN3(n4139), .DIN4(
        n4140) );
  nnd2s1 U6022 ( .Q(n4140), .DIN1(n3469), .DIN2(n3867) );
  xor2s1 U6023 ( .Q(n3867), .DIN1(n4141), .DIN2(n4142) );
  xor2s1 U6024 ( .Q(n4142), .DIN1(WX8517), .DIN2(n3131) );
  xor2s1 U6025 ( .Q(n4141), .DIN1(n3227), .DIN2(WX8581) );
  nnd2s1 U6026 ( .Q(n4139), .DIN1(n3449), .DIN2(n4143) );
  nnd2s1 U6027 ( .Q(n4138), .DIN1(WX7000), .DIN2(n3513) );
  nnd2s1 U6028 ( .Q(n4137), .DIN1(CRC_OUT_4_6), .DIN2(n3545) );
  nnd4s1 U6029 ( .Q(WX7157), .DIN1(n4144), .DIN2(n4145), .DIN3(n4146), .DIN4(
        n4147) );
  nnd2s1 U6030 ( .Q(n4147), .DIN1(n3469), .DIN2(n3874) );
  xor2s1 U6031 ( .Q(n3874), .DIN1(n4148), .DIN2(n4149) );
  xor2s1 U6032 ( .Q(n4149), .DIN1(WX8515), .DIN2(n3132) );
  xor2s1 U6033 ( .Q(n4148), .DIN1(n3228), .DIN2(WX8579) );
  nnd2s1 U6034 ( .Q(n4146), .DIN1(n3449), .DIN2(n4150) );
  nnd2s1 U6035 ( .Q(n4145), .DIN1(WX6998), .DIN2(n3513) );
  nnd2s1 U6036 ( .Q(n4144), .DIN1(CRC_OUT_4_7), .DIN2(n3545) );
  nnd4s1 U6037 ( .Q(WX7155), .DIN1(n4151), .DIN2(n4152), .DIN3(n4153), .DIN4(
        n4154) );
  nnd2s1 U6038 ( .Q(n4154), .DIN1(n3469), .DIN2(n3881) );
  xor2s1 U6039 ( .Q(n3881), .DIN1(n4155), .DIN2(n4156) );
  xor2s1 U6040 ( .Q(n4156), .DIN1(WX8513), .DIN2(n3133) );
  xor2s1 U6041 ( .Q(n4155), .DIN1(n3229), .DIN2(WX8577) );
  nnd2s1 U6042 ( .Q(n4153), .DIN1(n3449), .DIN2(n4157) );
  nnd2s1 U6043 ( .Q(n4152), .DIN1(WX6996), .DIN2(n3512) );
  nnd2s1 U6044 ( .Q(n4151), .DIN1(CRC_OUT_4_8), .DIN2(n3544) );
  nnd4s1 U6045 ( .Q(WX7153), .DIN1(n4158), .DIN2(n4159), .DIN3(n4160), .DIN4(
        n4161) );
  nnd2s1 U6046 ( .Q(n4161), .DIN1(n3469), .DIN2(n3888) );
  xor2s1 U6047 ( .Q(n3888), .DIN1(n4162), .DIN2(n4163) );
  xor2s1 U6048 ( .Q(n4163), .DIN1(WX8511), .DIN2(n3134) );
  xor2s1 U6049 ( .Q(n4162), .DIN1(n3230), .DIN2(WX8575) );
  nnd2s1 U6050 ( .Q(n4160), .DIN1(n3449), .DIN2(n4164) );
  nnd2s1 U6051 ( .Q(n4159), .DIN1(WX6994), .DIN2(n3512) );
  nnd2s1 U6052 ( .Q(n4158), .DIN1(CRC_OUT_4_9), .DIN2(n3544) );
  nnd4s1 U6053 ( .Q(WX7151), .DIN1(n4165), .DIN2(n4166), .DIN3(n4167), .DIN4(
        n4168) );
  nnd2s1 U6054 ( .Q(n4168), .DIN1(n3469), .DIN2(n3895) );
  xor2s1 U6055 ( .Q(n3895), .DIN1(n4169), .DIN2(n4170) );
  xor2s1 U6056 ( .Q(n4170), .DIN1(WX8509), .DIN2(n3135) );
  xor2s1 U6057 ( .Q(n4169), .DIN1(n3231), .DIN2(WX8573) );
  nnd2s1 U6058 ( .Q(n4167), .DIN1(n3449), .DIN2(n4171) );
  nnd2s1 U6059 ( .Q(n4166), .DIN1(WX6992), .DIN2(n3512) );
  nnd2s1 U6060 ( .Q(n4165), .DIN1(CRC_OUT_4_10), .DIN2(n3544) );
  nnd4s1 U6061 ( .Q(WX7149), .DIN1(n4172), .DIN2(n4173), .DIN3(n4174), .DIN4(
        n4175) );
  nnd2s1 U6062 ( .Q(n4175), .DIN1(n3469), .DIN2(n3902) );
  xor2s1 U6063 ( .Q(n3902), .DIN1(n4176), .DIN2(n4177) );
  xor2s1 U6064 ( .Q(n4177), .DIN1(WX8507), .DIN2(n3136) );
  xor2s1 U6065 ( .Q(n4176), .DIN1(n3232), .DIN2(WX8571) );
  nnd2s1 U6066 ( .Q(n4174), .DIN1(n3449), .DIN2(n4178) );
  nnd2s1 U6067 ( .Q(n4173), .DIN1(WX6990), .DIN2(n3512) );
  nnd2s1 U6068 ( .Q(n4172), .DIN1(CRC_OUT_4_11), .DIN2(n3544) );
  nnd4s1 U6069 ( .Q(WX7147), .DIN1(n4179), .DIN2(n4180), .DIN3(n4181), .DIN4(
        n4182) );
  nnd2s1 U6070 ( .Q(n4182), .DIN1(n3469), .DIN2(n3909) );
  xor2s1 U6071 ( .Q(n3909), .DIN1(n4183), .DIN2(n4184) );
  xor2s1 U6072 ( .Q(n4184), .DIN1(WX8505), .DIN2(n3137) );
  xor2s1 U6073 ( .Q(n4183), .DIN1(n3233), .DIN2(WX8569) );
  nnd2s1 U6074 ( .Q(n4181), .DIN1(n3449), .DIN2(n4185) );
  nnd2s1 U6075 ( .Q(n4180), .DIN1(WX6988), .DIN2(n3512) );
  nnd2s1 U6076 ( .Q(n4179), .DIN1(CRC_OUT_4_12), .DIN2(n3544) );
  nnd4s1 U6077 ( .Q(WX7145), .DIN1(n4186), .DIN2(n4187), .DIN3(n4188), .DIN4(
        n4189) );
  nnd2s1 U6078 ( .Q(n4189), .DIN1(n3469), .DIN2(n3916) );
  xor2s1 U6079 ( .Q(n3916), .DIN1(n4190), .DIN2(n4191) );
  xor2s1 U6080 ( .Q(n4191), .DIN1(WX8503), .DIN2(n3138) );
  xor2s1 U6081 ( .Q(n4190), .DIN1(n3234), .DIN2(WX8567) );
  nnd2s1 U6082 ( .Q(n4188), .DIN1(n3449), .DIN2(n4192) );
  nnd2s1 U6083 ( .Q(n4187), .DIN1(WX6986), .DIN2(n3512) );
  nnd2s1 U6084 ( .Q(n4186), .DIN1(CRC_OUT_4_13), .DIN2(n3544) );
  nnd4s1 U6085 ( .Q(WX7143), .DIN1(n4193), .DIN2(n4194), .DIN3(n4195), .DIN4(
        n4196) );
  nnd2s1 U6086 ( .Q(n4196), .DIN1(n3470), .DIN2(n3923) );
  xor2s1 U6087 ( .Q(n3923), .DIN1(n4197), .DIN2(n4198) );
  xor2s1 U6088 ( .Q(n4198), .DIN1(WX8501), .DIN2(n3139) );
  xor2s1 U6089 ( .Q(n4197), .DIN1(n3235), .DIN2(WX8565) );
  nnd2s1 U6090 ( .Q(n4195), .DIN1(n3449), .DIN2(n4199) );
  nnd2s1 U6091 ( .Q(n4194), .DIN1(WX6984), .DIN2(n3512) );
  nnd2s1 U6092 ( .Q(n4193), .DIN1(CRC_OUT_4_14), .DIN2(n3544) );
  nnd4s1 U6093 ( .Q(WX7141), .DIN1(n4200), .DIN2(n4201), .DIN3(n4202), .DIN4(
        n4203) );
  nnd2s1 U6094 ( .Q(n4203), .DIN1(n3470), .DIN2(n3930) );
  xor2s1 U6095 ( .Q(n3930), .DIN1(n4204), .DIN2(n4205) );
  xor2s1 U6096 ( .Q(n4205), .DIN1(WX8499), .DIN2(n3140) );
  xor2s1 U6097 ( .Q(n4204), .DIN1(n3236), .DIN2(WX8563) );
  nnd2s1 U6098 ( .Q(n4202), .DIN1(n3449), .DIN2(n4206) );
  nnd2s1 U6099 ( .Q(n4201), .DIN1(WX6982), .DIN2(n3512) );
  nnd2s1 U6100 ( .Q(n4200), .DIN1(CRC_OUT_4_15), .DIN2(n3544) );
  and2s1 U6101 ( .Q(WX714), .DIN1(RESET), .DIN2(WX651) );
  nnd4s1 U6102 ( .Q(WX7139), .DIN1(n4207), .DIN2(n4208), .DIN3(n4209), .DIN4(
        n4210) );
  nnd2s1 U6103 ( .Q(n4210), .DIN1(n3470), .DIN2(n3939) );
  xor2s1 U6104 ( .Q(n3939), .DIN1(n4211), .DIN2(n4212) );
  xor2s1 U6105 ( .Q(n4212), .DIN1(n3561), .DIN2(WX8433) );
  xor2s1 U6106 ( .Q(n4211), .DIN1(n2965), .DIN2(n4213) );
  xor2s1 U6107 ( .Q(n4213), .DIN1(WX8625), .DIN2(WX8561) );
  nnd2s1 U6108 ( .Q(n4209), .DIN1(n3448), .DIN2(n4214) );
  nnd2s1 U6109 ( .Q(n4208), .DIN1(WX6980), .DIN2(n3512) );
  nnd2s1 U6110 ( .Q(n4207), .DIN1(CRC_OUT_4_16), .DIN2(n3544) );
  nnd4s1 U6111 ( .Q(WX7137), .DIN1(n4215), .DIN2(n4216), .DIN3(n4217), .DIN4(
        n4218) );
  nnd2s1 U6112 ( .Q(n4218), .DIN1(n3470), .DIN2(n3947) );
  xor2s1 U6113 ( .Q(n3947), .DIN1(n4219), .DIN2(n4220) );
  xor2s1 U6114 ( .Q(n4220), .DIN1(n3561), .DIN2(WX8431) );
  xor2s1 U6115 ( .Q(n4219), .DIN1(n2966), .DIN2(n4221) );
  xor2s1 U6116 ( .Q(n4221), .DIN1(WX8623), .DIN2(WX8559) );
  nnd2s1 U6117 ( .Q(n4217), .DIN1(n3448), .DIN2(n4222) );
  nnd2s1 U6118 ( .Q(n4216), .DIN1(WX6978), .DIN2(n3512) );
  nnd2s1 U6119 ( .Q(n4215), .DIN1(CRC_OUT_4_17), .DIN2(n3544) );
  nnd4s1 U6120 ( .Q(WX7135), .DIN1(n4223), .DIN2(n4224), .DIN3(n4225), .DIN4(
        n4226) );
  nnd2s1 U6121 ( .Q(n4226), .DIN1(n3470), .DIN2(n3955) );
  xor2s1 U6122 ( .Q(n3955), .DIN1(n4227), .DIN2(n4228) );
  xor2s1 U6123 ( .Q(n4228), .DIN1(n3561), .DIN2(WX8429) );
  xor2s1 U6124 ( .Q(n4227), .DIN1(n2967), .DIN2(n4229) );
  xor2s1 U6125 ( .Q(n4229), .DIN1(WX8621), .DIN2(WX8557) );
  nnd2s1 U6126 ( .Q(n4225), .DIN1(n3448), .DIN2(n4230) );
  nnd2s1 U6127 ( .Q(n4224), .DIN1(WX6976), .DIN2(n3512) );
  nnd2s1 U6128 ( .Q(n4223), .DIN1(CRC_OUT_4_18), .DIN2(n3544) );
  nnd4s1 U6129 ( .Q(WX7133), .DIN1(n4231), .DIN2(n4232), .DIN3(n4233), .DIN4(
        n4234) );
  nnd2s1 U6130 ( .Q(n4234), .DIN1(n3470), .DIN2(n3963) );
  xor2s1 U6131 ( .Q(n3963), .DIN1(n4235), .DIN2(n4236) );
  xor2s1 U6132 ( .Q(n4236), .DIN1(n3561), .DIN2(WX8427) );
  xor2s1 U6133 ( .Q(n4235), .DIN1(n2968), .DIN2(n4237) );
  xor2s1 U6134 ( .Q(n4237), .DIN1(WX8619), .DIN2(WX8555) );
  nnd2s1 U6135 ( .Q(n4233), .DIN1(n3448), .DIN2(n4238) );
  nnd2s1 U6136 ( .Q(n4232), .DIN1(WX6974), .DIN2(n3512) );
  nnd2s1 U6137 ( .Q(n4231), .DIN1(CRC_OUT_4_19), .DIN2(n3544) );
  nnd4s1 U6138 ( .Q(WX7131), .DIN1(n4239), .DIN2(n4240), .DIN3(n4241), .DIN4(
        n4242) );
  nnd2s1 U6139 ( .Q(n4242), .DIN1(n3470), .DIN2(n3971) );
  xor2s1 U6140 ( .Q(n3971), .DIN1(n4243), .DIN2(n4244) );
  xor2s1 U6141 ( .Q(n4244), .DIN1(n3561), .DIN2(WX8425) );
  xor2s1 U6142 ( .Q(n4243), .DIN1(n2969), .DIN2(n4245) );
  xor2s1 U6143 ( .Q(n4245), .DIN1(WX8617), .DIN2(WX8553) );
  nnd2s1 U6144 ( .Q(n4241), .DIN1(n3448), .DIN2(n4246) );
  nnd2s1 U6145 ( .Q(n4240), .DIN1(WX6972), .DIN2(n3511) );
  nnd2s1 U6146 ( .Q(n4239), .DIN1(CRC_OUT_4_20), .DIN2(n3543) );
  nnd4s1 U6147 ( .Q(WX7129), .DIN1(n4247), .DIN2(n4248), .DIN3(n4249), .DIN4(
        n4250) );
  nnd2s1 U6148 ( .Q(n4250), .DIN1(n3470), .DIN2(n3979) );
  xor2s1 U6149 ( .Q(n3979), .DIN1(n4251), .DIN2(n4252) );
  xor2s1 U6150 ( .Q(n4252), .DIN1(n3562), .DIN2(WX8423) );
  xor2s1 U6151 ( .Q(n4251), .DIN1(n2970), .DIN2(n4253) );
  xor2s1 U6152 ( .Q(n4253), .DIN1(WX8615), .DIN2(WX8551) );
  nnd2s1 U6153 ( .Q(n4249), .DIN1(n3448), .DIN2(n4254) );
  nnd2s1 U6154 ( .Q(n4248), .DIN1(WX6970), .DIN2(n3511) );
  nnd2s1 U6155 ( .Q(n4247), .DIN1(CRC_OUT_4_21), .DIN2(n3543) );
  nnd4s1 U6156 ( .Q(WX7127), .DIN1(n4255), .DIN2(n4256), .DIN3(n4257), .DIN4(
        n4258) );
  nnd2s1 U6157 ( .Q(n4258), .DIN1(n3470), .DIN2(n3987) );
  xor2s1 U6158 ( .Q(n3987), .DIN1(n4259), .DIN2(n4260) );
  xor2s1 U6159 ( .Q(n4260), .DIN1(n3562), .DIN2(WX8421) );
  xor2s1 U6160 ( .Q(n4259), .DIN1(n2971), .DIN2(n4261) );
  xor2s1 U6161 ( .Q(n4261), .DIN1(WX8613), .DIN2(WX8549) );
  nnd2s1 U6162 ( .Q(n4257), .DIN1(n3448), .DIN2(n4262) );
  nnd2s1 U6163 ( .Q(n4256), .DIN1(WX6968), .DIN2(n3511) );
  nnd2s1 U6164 ( .Q(n4255), .DIN1(CRC_OUT_4_22), .DIN2(n3543) );
  nnd4s1 U6165 ( .Q(WX7125), .DIN1(n4263), .DIN2(n4264), .DIN3(n4265), .DIN4(
        n4266) );
  nnd2s1 U6166 ( .Q(n4266), .DIN1(n3470), .DIN2(n3995) );
  xor2s1 U6167 ( .Q(n3995), .DIN1(n4267), .DIN2(n4268) );
  xor2s1 U6168 ( .Q(n4268), .DIN1(n3562), .DIN2(WX8419) );
  xor2s1 U6169 ( .Q(n4267), .DIN1(n2972), .DIN2(n4269) );
  xor2s1 U6170 ( .Q(n4269), .DIN1(WX8611), .DIN2(WX8547) );
  nnd2s1 U6171 ( .Q(n4265), .DIN1(n3448), .DIN2(n4270) );
  nnd2s1 U6172 ( .Q(n4264), .DIN1(WX6966), .DIN2(n3511) );
  nnd2s1 U6173 ( .Q(n4263), .DIN1(CRC_OUT_4_23), .DIN2(n3543) );
  nnd4s1 U6174 ( .Q(WX7123), .DIN1(n4271), .DIN2(n4272), .DIN3(n4273), .DIN4(
        n4274) );
  nnd2s1 U6175 ( .Q(n4274), .DIN1(n3470), .DIN2(n4003) );
  xor2s1 U6176 ( .Q(n4003), .DIN1(n4275), .DIN2(n4276) );
  xor2s1 U6177 ( .Q(n4276), .DIN1(n3562), .DIN2(WX8417) );
  xor2s1 U6178 ( .Q(n4275), .DIN1(n2973), .DIN2(n4277) );
  xor2s1 U6179 ( .Q(n4277), .DIN1(WX8609), .DIN2(WX8545) );
  nnd2s1 U6180 ( .Q(n4273), .DIN1(n3448), .DIN2(n4278) );
  nnd2s1 U6181 ( .Q(n4272), .DIN1(WX6964), .DIN2(n3511) );
  nnd2s1 U6182 ( .Q(n4271), .DIN1(CRC_OUT_4_24), .DIN2(n3543) );
  nnd4s1 U6183 ( .Q(WX7121), .DIN1(n4279), .DIN2(n4280), .DIN3(n4281), .DIN4(
        n4282) );
  nnd2s1 U6184 ( .Q(n4282), .DIN1(n3470), .DIN2(n4011) );
  xor2s1 U6185 ( .Q(n4011), .DIN1(n4283), .DIN2(n4284) );
  xor2s1 U6186 ( .Q(n4284), .DIN1(n3562), .DIN2(WX8415) );
  xor2s1 U6187 ( .Q(n4283), .DIN1(n2974), .DIN2(n4285) );
  xor2s1 U6188 ( .Q(n4285), .DIN1(WX8607), .DIN2(WX8543) );
  nnd2s1 U6189 ( .Q(n4281), .DIN1(n3448), .DIN2(n4286) );
  nnd2s1 U6190 ( .Q(n4280), .DIN1(WX6962), .DIN2(n3511) );
  nnd2s1 U6191 ( .Q(n4279), .DIN1(CRC_OUT_4_25), .DIN2(n3543) );
  and2s1 U6192 ( .Q(WX712), .DIN1(RESET), .DIN2(WX649) );
  nnd4s1 U6193 ( .Q(WX7119), .DIN1(n4287), .DIN2(n4288), .DIN3(n4289), .DIN4(
        n4290) );
  nnd2s1 U6194 ( .Q(n4290), .DIN1(n3470), .DIN2(n4019) );
  xor2s1 U6195 ( .Q(n4019), .DIN1(n4291), .DIN2(n4292) );
  xor2s1 U6196 ( .Q(n4292), .DIN1(n3562), .DIN2(WX8413) );
  xor2s1 U6197 ( .Q(n4291), .DIN1(n2975), .DIN2(n4293) );
  xor2s1 U6198 ( .Q(n4293), .DIN1(WX8605), .DIN2(WX8541) );
  nnd2s1 U6199 ( .Q(n4289), .DIN1(n3448), .DIN2(n4294) );
  nnd2s1 U6200 ( .Q(n4288), .DIN1(WX6960), .DIN2(n3511) );
  nnd2s1 U6201 ( .Q(n4287), .DIN1(CRC_OUT_4_26), .DIN2(n3543) );
  nnd4s1 U6202 ( .Q(WX7117), .DIN1(n4295), .DIN2(n4296), .DIN3(n4297), .DIN4(
        n4298) );
  nnd2s1 U6203 ( .Q(n4298), .DIN1(n3471), .DIN2(n4027) );
  xor2s1 U6204 ( .Q(n4027), .DIN1(n4299), .DIN2(n4300) );
  xor2s1 U6205 ( .Q(n4300), .DIN1(n3562), .DIN2(WX8411) );
  xor2s1 U6206 ( .Q(n4299), .DIN1(n2976), .DIN2(n4301) );
  xor2s1 U6207 ( .Q(n4301), .DIN1(WX8603), .DIN2(WX8539) );
  nnd2s1 U6208 ( .Q(n4297), .DIN1(n3448), .DIN2(n4302) );
  nnd2s1 U6209 ( .Q(n4296), .DIN1(WX6958), .DIN2(n3511) );
  nnd2s1 U6210 ( .Q(n4295), .DIN1(CRC_OUT_4_27), .DIN2(n3543) );
  nnd4s1 U6211 ( .Q(WX7115), .DIN1(n4303), .DIN2(n4304), .DIN3(n4305), .DIN4(
        n4306) );
  nnd2s1 U6212 ( .Q(n4306), .DIN1(n3471), .DIN2(n4035) );
  xor2s1 U6213 ( .Q(n4035), .DIN1(n4307), .DIN2(n4308) );
  xor2s1 U6214 ( .Q(n4308), .DIN1(n3563), .DIN2(WX8409) );
  xor2s1 U6215 ( .Q(n4307), .DIN1(n2977), .DIN2(n4309) );
  xor2s1 U6216 ( .Q(n4309), .DIN1(WX8601), .DIN2(WX8537) );
  nnd2s1 U6217 ( .Q(n4305), .DIN1(n3448), .DIN2(n4310) );
  nnd2s1 U6218 ( .Q(n4304), .DIN1(WX6956), .DIN2(n3511) );
  nnd2s1 U6219 ( .Q(n4303), .DIN1(CRC_OUT_4_28), .DIN2(n3543) );
  nnd4s1 U6220 ( .Q(WX7113), .DIN1(n4311), .DIN2(n4312), .DIN3(n4313), .DIN4(
        n4314) );
  nnd2s1 U6221 ( .Q(n4314), .DIN1(n3471), .DIN2(n4043) );
  xor2s1 U6222 ( .Q(n4043), .DIN1(n4315), .DIN2(n4316) );
  xor2s1 U6223 ( .Q(n4316), .DIN1(n3563), .DIN2(WX8407) );
  xor2s1 U6224 ( .Q(n4315), .DIN1(n2978), .DIN2(n4317) );
  xor2s1 U6225 ( .Q(n4317), .DIN1(WX8599), .DIN2(WX8535) );
  nnd2s1 U6226 ( .Q(n4313), .DIN1(n3447), .DIN2(n4318) );
  nnd2s1 U6227 ( .Q(n4312), .DIN1(WX6954), .DIN2(n3511) );
  nnd2s1 U6228 ( .Q(n4311), .DIN1(CRC_OUT_4_29), .DIN2(n3543) );
  nnd4s1 U6229 ( .Q(WX7111), .DIN1(n4319), .DIN2(n4320), .DIN3(n4321), .DIN4(
        n4322) );
  nnd2s1 U6230 ( .Q(n4322), .DIN1(n3471), .DIN2(n4051) );
  xor2s1 U6231 ( .Q(n4051), .DIN1(n4323), .DIN2(n4324) );
  xor2s1 U6232 ( .Q(n4324), .DIN1(n3563), .DIN2(WX8405) );
  xor2s1 U6233 ( .Q(n4323), .DIN1(n2979), .DIN2(n4325) );
  xor2s1 U6234 ( .Q(n4325), .DIN1(WX8597), .DIN2(WX8533) );
  nnd2s1 U6235 ( .Q(n4321), .DIN1(n3447), .DIN2(n4326) );
  nnd2s1 U6236 ( .Q(n4320), .DIN1(WX6952), .DIN2(n3511) );
  nnd2s1 U6237 ( .Q(n4319), .DIN1(CRC_OUT_4_30), .DIN2(n3543) );
  nnd4s1 U6238 ( .Q(WX7109), .DIN1(n4327), .DIN2(n4328), .DIN3(n4329), .DIN4(
        n4330) );
  nnd2s1 U6239 ( .Q(n4330), .DIN1(n3471), .DIN2(n4059) );
  xor2s1 U6240 ( .Q(n4059), .DIN1(n4331), .DIN2(n4332) );
  xor2s1 U6241 ( .Q(n4332), .DIN1(n3563), .DIN2(WX8403) );
  xor2s1 U6242 ( .Q(n4331), .DIN1(n2980), .DIN2(n4333) );
  xor2s1 U6243 ( .Q(n4333), .DIN1(WX8595), .DIN2(WX8531) );
  nnd2s1 U6244 ( .Q(n4329), .DIN1(n3447), .DIN2(n4334) );
  nnd2s1 U6245 ( .Q(n4328), .DIN1(WX6950), .DIN2(n3511) );
  nnd2s1 U6246 ( .Q(n4327), .DIN1(CRC_OUT_4_31), .DIN2(n3543) );
  and2s1 U6247 ( .Q(WX710), .DIN1(RESET), .DIN2(WX647) );
  and2s1 U6248 ( .Q(WX708), .DIN1(RESET), .DIN2(WX645) );
  nnd4s1 U6249 ( .Q(WX706), .DIN1(n4335), .DIN2(n4336), .DIN3(n4337), .DIN4(
        n4338) );
  nnd2s1 U6250 ( .Q(n4338), .DIN1(n3471), .DIN2(n4339) );
  nnd2s1 U6251 ( .Q(n4337), .DIN1(n3447), .DIN2(n4340) );
  hi1s1 U6252 ( .Q(n4340), .DIN(n4341) );
  nnd2s1 U6253 ( .Q(n4336), .DIN1(WX547), .DIN2(n3510) );
  nnd2s1 U6254 ( .Q(n4335), .DIN1(CRC_OUT_9_0), .DIN2(n3542) );
  nnd4s1 U6255 ( .Q(WX704), .DIN1(n4342), .DIN2(n4343), .DIN3(n4344), .DIN4(
        n4345) );
  nnd2s1 U6256 ( .Q(n4345), .DIN1(n3471), .DIN2(n4346) );
  nnd2s1 U6257 ( .Q(n4344), .DIN1(n3447), .DIN2(n4347) );
  hi1s1 U6258 ( .Q(n4347), .DIN(n4348) );
  nnd2s1 U6259 ( .Q(n4343), .DIN1(WX545), .DIN2(n3510) );
  nnd2s1 U6260 ( .Q(n4342), .DIN1(CRC_OUT_9_1), .DIN2(n3542) );
  nnd4s1 U6261 ( .Q(WX702), .DIN1(n4349), .DIN2(n4350), .DIN3(n4351), .DIN4(
        n4352) );
  nnd2s1 U6262 ( .Q(n4352), .DIN1(n3471), .DIN2(n4353) );
  nnd2s1 U6263 ( .Q(n4351), .DIN1(n3447), .DIN2(n4354) );
  hi1s1 U6264 ( .Q(n4354), .DIN(n4355) );
  nnd2s1 U6265 ( .Q(n4350), .DIN1(WX543), .DIN2(n3510) );
  nnd2s1 U6266 ( .Q(n4349), .DIN1(CRC_OUT_9_2), .DIN2(n3542) );
  nor2s1 U6267 ( .Q(WX7011), .DIN1(WX6950), .DIN2(n3363) );
  and2s1 U6268 ( .Q(WX7009), .DIN1(RESET), .DIN2(WX7012) );
  and2s1 U6269 ( .Q(WX7007), .DIN1(RESET), .DIN2(WX7010) );
  and2s1 U6270 ( .Q(WX7005), .DIN1(RESET), .DIN2(WX7008) );
  and2s1 U6271 ( .Q(WX7003), .DIN1(RESET), .DIN2(WX7006) );
  and2s1 U6272 ( .Q(WX7001), .DIN1(RESET), .DIN2(WX7004) );
  nnd4s1 U6273 ( .Q(WX700), .DIN1(n4356), .DIN2(n4357), .DIN3(n4358), .DIN4(
        n4359) );
  nnd2s1 U6274 ( .Q(n4359), .DIN1(n3471), .DIN2(n4360) );
  nnd2s1 U6275 ( .Q(n4358), .DIN1(n3447), .DIN2(n4361) );
  hi1s1 U6276 ( .Q(n4361), .DIN(n4362) );
  nnd2s1 U6277 ( .Q(n4357), .DIN1(WX541), .DIN2(n3510) );
  nnd2s1 U6278 ( .Q(n4356), .DIN1(CRC_OUT_9_3), .DIN2(n3542) );
  and2s1 U6279 ( .Q(WX6999), .DIN1(RESET), .DIN2(WX7002) );
  and2s1 U6280 ( .Q(WX6997), .DIN1(RESET), .DIN2(WX7000) );
  and2s1 U6281 ( .Q(WX6995), .DIN1(RESET), .DIN2(WX6998) );
  and2s1 U6282 ( .Q(WX6993), .DIN1(RESET), .DIN2(WX6996) );
  and2s1 U6283 ( .Q(WX6991), .DIN1(RESET), .DIN2(WX6994) );
  and2s1 U6284 ( .Q(WX6989), .DIN1(RESET), .DIN2(WX6992) );
  and2s1 U6285 ( .Q(WX6987), .DIN1(RESET), .DIN2(WX6990) );
  and2s1 U6286 ( .Q(WX6985), .DIN1(RESET), .DIN2(WX6988) );
  and2s1 U6287 ( .Q(WX6983), .DIN1(RESET), .DIN2(WX6986) );
  and2s1 U6288 ( .Q(WX6981), .DIN1(RESET), .DIN2(WX6984) );
  nnd4s1 U6289 ( .Q(WX698), .DIN1(n4363), .DIN2(n4364), .DIN3(n4365), .DIN4(
        n4366) );
  nnd2s1 U6290 ( .Q(n4366), .DIN1(n3471), .DIN2(n4367) );
  nnd2s1 U6291 ( .Q(n4365), .DIN1(n3447), .DIN2(n4368) );
  hi1s1 U6292 ( .Q(n4368), .DIN(n4369) );
  nnd2s1 U6293 ( .Q(n4364), .DIN1(WX539), .DIN2(n3510) );
  nnd2s1 U6294 ( .Q(n4363), .DIN1(CRC_OUT_9_4), .DIN2(n3542) );
  and2s1 U6295 ( .Q(WX6979), .DIN1(RESET), .DIN2(WX6982) );
  and2s1 U6296 ( .Q(WX6977), .DIN1(RESET), .DIN2(WX6980) );
  and2s1 U6297 ( .Q(WX6975), .DIN1(RESET), .DIN2(WX6978) );
  and2s1 U6298 ( .Q(WX6973), .DIN1(RESET), .DIN2(WX6976) );
  and2s1 U6299 ( .Q(WX6971), .DIN1(RESET), .DIN2(WX6974) );
  and2s1 U6300 ( .Q(WX6969), .DIN1(RESET), .DIN2(WX6972) );
  and2s1 U6301 ( .Q(WX6967), .DIN1(RESET), .DIN2(WX6970) );
  and2s1 U6302 ( .Q(WX6965), .DIN1(RESET), .DIN2(WX6968) );
  and2s1 U6303 ( .Q(WX6963), .DIN1(RESET), .DIN2(WX6966) );
  and2s1 U6304 ( .Q(WX6961), .DIN1(RESET), .DIN2(WX6964) );
  nnd4s1 U6305 ( .Q(WX696), .DIN1(n4370), .DIN2(n4371), .DIN3(n4372), .DIN4(
        n4373) );
  nnd2s1 U6306 ( .Q(n4373), .DIN1(n3471), .DIN2(n4374) );
  nnd2s1 U6307 ( .Q(n4372), .DIN1(n3447), .DIN2(n4375) );
  hi1s1 U6308 ( .Q(n4375), .DIN(n4376) );
  nnd2s1 U6309 ( .Q(n4371), .DIN1(WX537), .DIN2(n3510) );
  nnd2s1 U6310 ( .Q(n4370), .DIN1(CRC_OUT_9_5), .DIN2(n3542) );
  and2s1 U6311 ( .Q(WX6959), .DIN1(RESET), .DIN2(WX6962) );
  and2s1 U6312 ( .Q(WX6957), .DIN1(RESET), .DIN2(WX6960) );
  and2s1 U6313 ( .Q(WX6955), .DIN1(RESET), .DIN2(WX6958) );
  and2s1 U6314 ( .Q(WX6953), .DIN1(RESET), .DIN2(WX6956) );
  and2s1 U6315 ( .Q(WX6951), .DIN1(RESET), .DIN2(WX6954) );
  and2s1 U6316 ( .Q(WX6949), .DIN1(RESET), .DIN2(WX6952) );
  nnd4s1 U6317 ( .Q(WX694), .DIN1(n4377), .DIN2(n4378), .DIN3(n4379), .DIN4(
        n4380) );
  nnd2s1 U6318 ( .Q(n4380), .DIN1(n3471), .DIN2(n4381) );
  nnd2s1 U6319 ( .Q(n4379), .DIN1(n3447), .DIN2(n4382) );
  hi1s1 U6320 ( .Q(n4382), .DIN(n4383) );
  nnd2s1 U6321 ( .Q(n4378), .DIN1(WX535), .DIN2(n3510) );
  nnd2s1 U6322 ( .Q(n4377), .DIN1(CRC_OUT_9_6), .DIN2(n3542) );
  nnd4s1 U6323 ( .Q(WX692), .DIN1(n4384), .DIN2(n4385), .DIN3(n4386), .DIN4(
        n4387) );
  nnd2s1 U6324 ( .Q(n4387), .DIN1(n3471), .DIN2(n4388) );
  nnd2s1 U6325 ( .Q(n4386), .DIN1(n3447), .DIN2(n4389) );
  hi1s1 U6326 ( .Q(n4389), .DIN(n4390) );
  nnd2s1 U6327 ( .Q(n4385), .DIN1(WX533), .DIN2(n3510) );
  nnd2s1 U6328 ( .Q(n4384), .DIN1(CRC_OUT_9_7), .DIN2(n3542) );
  nnd4s1 U6329 ( .Q(WX690), .DIN1(n4391), .DIN2(n4392), .DIN3(n4393), .DIN4(
        n4394) );
  nnd2s1 U6330 ( .Q(n4394), .DIN1(n3472), .DIN2(n4395) );
  nnd2s1 U6331 ( .Q(n4393), .DIN1(n3447), .DIN2(n4396) );
  hi1s1 U6332 ( .Q(n4396), .DIN(n4397) );
  nnd2s1 U6333 ( .Q(n4392), .DIN1(WX531), .DIN2(n3510) );
  nnd2s1 U6334 ( .Q(n4391), .DIN1(CRC_OUT_9_8), .DIN2(n3542) );
  nnd4s1 U6335 ( .Q(WX688), .DIN1(n4398), .DIN2(n4399), .DIN3(n4400), .DIN4(
        n4401) );
  nnd2s1 U6336 ( .Q(n4401), .DIN1(n3472), .DIN2(n4402) );
  nnd2s1 U6337 ( .Q(n4400), .DIN1(n3447), .DIN2(n4403) );
  hi1s1 U6338 ( .Q(n4403), .DIN(n4404) );
  nnd2s1 U6339 ( .Q(n4399), .DIN1(WX529), .DIN2(n3510) );
  nnd2s1 U6340 ( .Q(n4398), .DIN1(CRC_OUT_9_9), .DIN2(n3542) );
  nnd4s1 U6341 ( .Q(WX686), .DIN1(n4405), .DIN2(n4406), .DIN3(n4407), .DIN4(
        n4408) );
  nnd2s1 U6342 ( .Q(n4408), .DIN1(n3472), .DIN2(n4409) );
  nnd2s1 U6343 ( .Q(n4407), .DIN1(n3446), .DIN2(n4410) );
  hi1s1 U6344 ( .Q(n4410), .DIN(n4411) );
  nnd2s1 U6345 ( .Q(n4406), .DIN1(WX527), .DIN2(n3510) );
  nnd2s1 U6346 ( .Q(n4405), .DIN1(CRC_OUT_9_10), .DIN2(n3542) );
  nnd4s1 U6347 ( .Q(WX684), .DIN1(n4412), .DIN2(n4413), .DIN3(n4414), .DIN4(
        n4415) );
  nnd2s1 U6348 ( .Q(n4415), .DIN1(n3472), .DIN2(n4416) );
  nnd2s1 U6349 ( .Q(n4414), .DIN1(n3446), .DIN2(n4417) );
  hi1s1 U6350 ( .Q(n4417), .DIN(n4418) );
  nnd2s1 U6351 ( .Q(n4413), .DIN1(WX525), .DIN2(n3510) );
  nnd2s1 U6352 ( .Q(n4412), .DIN1(CRC_OUT_9_11), .DIN2(n3542) );
  nnd4s1 U6353 ( .Q(WX682), .DIN1(n4419), .DIN2(n4420), .DIN3(n4421), .DIN4(
        n4422) );
  nnd2s1 U6354 ( .Q(n4422), .DIN1(n3472), .DIN2(n4423) );
  nnd2s1 U6355 ( .Q(n4421), .DIN1(n3446), .DIN2(n4424) );
  hi1s1 U6356 ( .Q(n4424), .DIN(n4425) );
  nnd2s1 U6357 ( .Q(n4420), .DIN1(WX523), .DIN2(n3509) );
  nnd2s1 U6358 ( .Q(n4419), .DIN1(CRC_OUT_9_12), .DIN2(n3541) );
  nnd4s1 U6359 ( .Q(WX680), .DIN1(n4426), .DIN2(n4427), .DIN3(n4428), .DIN4(
        n4429) );
  nnd2s1 U6360 ( .Q(n4429), .DIN1(n3472), .DIN2(n4430) );
  nnd2s1 U6361 ( .Q(n4428), .DIN1(n3446), .DIN2(n4431) );
  hi1s1 U6362 ( .Q(n4431), .DIN(n4432) );
  nnd2s1 U6363 ( .Q(n4427), .DIN1(WX521), .DIN2(n3509) );
  nnd2s1 U6364 ( .Q(n4426), .DIN1(CRC_OUT_9_13), .DIN2(n3541) );
  nnd4s1 U6365 ( .Q(WX678), .DIN1(n4433), .DIN2(n4434), .DIN3(n4435), .DIN4(
        n4436) );
  nnd2s1 U6366 ( .Q(n4436), .DIN1(n3472), .DIN2(n4437) );
  nnd2s1 U6367 ( .Q(n4435), .DIN1(n3446), .DIN2(n4438) );
  hi1s1 U6368 ( .Q(n4438), .DIN(n4439) );
  nnd2s1 U6369 ( .Q(n4434), .DIN1(WX519), .DIN2(n3509) );
  nnd2s1 U6370 ( .Q(n4433), .DIN1(CRC_OUT_9_14), .DIN2(n3541) );
  nnd4s1 U6371 ( .Q(WX676), .DIN1(n4440), .DIN2(n4441), .DIN3(n4442), .DIN4(
        n4443) );
  nnd2s1 U6372 ( .Q(n4443), .DIN1(n3472), .DIN2(n4444) );
  nnd2s1 U6373 ( .Q(n4442), .DIN1(n3446), .DIN2(n4445) );
  hi1s1 U6374 ( .Q(n4445), .DIN(n4446) );
  nnd2s1 U6375 ( .Q(n4441), .DIN1(WX517), .DIN2(n3509) );
  nnd2s1 U6376 ( .Q(n4440), .DIN1(CRC_OUT_9_15), .DIN2(n3541) );
  nnd4s1 U6377 ( .Q(WX674), .DIN1(n4447), .DIN2(n4448), .DIN3(n4449), .DIN4(
        n4450) );
  nnd2s1 U6378 ( .Q(n4450), .DIN1(n3472), .DIN2(n4451) );
  nnd2s1 U6379 ( .Q(n4449), .DIN1(n3446), .DIN2(n4452) );
  hi1s1 U6380 ( .Q(n4452), .DIN(n4453) );
  nnd2s1 U6381 ( .Q(n4448), .DIN1(WX515), .DIN2(n3509) );
  nnd2s1 U6382 ( .Q(n4447), .DIN1(CRC_OUT_9_16), .DIN2(n3541) );
  nnd4s1 U6383 ( .Q(WX672), .DIN1(n4454), .DIN2(n4455), .DIN3(n4456), .DIN4(
        n4457) );
  nnd2s1 U6384 ( .Q(n4457), .DIN1(n3472), .DIN2(n4458) );
  nnd2s1 U6385 ( .Q(n4456), .DIN1(n3446), .DIN2(n4459) );
  hi1s1 U6386 ( .Q(n4459), .DIN(n4460) );
  nnd2s1 U6387 ( .Q(n4455), .DIN1(WX513), .DIN2(n3509) );
  nnd2s1 U6388 ( .Q(n4454), .DIN1(CRC_OUT_9_17), .DIN2(n3541) );
  nnd4s1 U6389 ( .Q(WX670), .DIN1(n4461), .DIN2(n4462), .DIN3(n4463), .DIN4(
        n4464) );
  nnd2s1 U6390 ( .Q(n4464), .DIN1(n3472), .DIN2(n4465) );
  nnd2s1 U6391 ( .Q(n4463), .DIN1(n3446), .DIN2(n4466) );
  hi1s1 U6392 ( .Q(n4466), .DIN(n4467) );
  nnd2s1 U6393 ( .Q(n4462), .DIN1(WX511), .DIN2(n3509) );
  nnd2s1 U6394 ( .Q(n4461), .DIN1(CRC_OUT_9_18), .DIN2(n3541) );
  nnd4s1 U6395 ( .Q(WX668), .DIN1(n4468), .DIN2(n4469), .DIN3(n4470), .DIN4(
        n4471) );
  nnd2s1 U6396 ( .Q(n4471), .DIN1(n3472), .DIN2(n4472) );
  nnd2s1 U6397 ( .Q(n4470), .DIN1(WX509), .DIN2(n3509) );
  nnd2s1 U6398 ( .Q(n4469), .DIN1(CRC_OUT_9_19), .DIN2(n3541) );
  nnd2s1 U6399 ( .Q(n4468), .DIN1(n3446), .DIN2(n4473) );
  hi1s1 U6400 ( .Q(n4473), .DIN(n4474) );
  nnd4s1 U6401 ( .Q(WX666), .DIN1(n4475), .DIN2(n4476), .DIN3(n4477), .DIN4(
        n4478) );
  nnd2s1 U6402 ( .Q(n4478), .DIN1(n3472), .DIN2(n4479) );
  nnd2s1 U6403 ( .Q(n4477), .DIN1(WX507), .DIN2(n3509) );
  nnd2s1 U6404 ( .Q(n4476), .DIN1(CRC_OUT_9_20), .DIN2(n3541) );
  nnd2s1 U6405 ( .Q(n4475), .DIN1(n3446), .DIN2(n4480) );
  hi1s1 U6406 ( .Q(n4480), .DIN(n4481) );
  nnd4s1 U6407 ( .Q(WX664), .DIN1(n4482), .DIN2(n4483), .DIN3(n4484), .DIN4(
        n4485) );
  nnd2s1 U6408 ( .Q(n4485), .DIN1(n3473), .DIN2(n4486) );
  nnd2s1 U6409 ( .Q(n4484), .DIN1(WX505), .DIN2(n3509) );
  nnd2s1 U6410 ( .Q(n4483), .DIN1(CRC_OUT_9_21), .DIN2(n3541) );
  nnd2s1 U6411 ( .Q(n4482), .DIN1(n3446), .DIN2(n4487) );
  hi1s1 U6412 ( .Q(n4487), .DIN(n4488) );
  nnd4s1 U6413 ( .Q(WX662), .DIN1(n4489), .DIN2(n4490), .DIN3(n4491), .DIN4(
        n4492) );
  nnd2s1 U6414 ( .Q(n4492), .DIN1(n3473), .DIN2(n4493) );
  nnd2s1 U6415 ( .Q(n4491), .DIN1(WX503), .DIN2(n3509) );
  nnd2s1 U6416 ( .Q(n4490), .DIN1(CRC_OUT_9_22), .DIN2(n3541) );
  nnd2s1 U6417 ( .Q(n4489), .DIN1(n3446), .DIN2(n4494) );
  hi1s1 U6418 ( .Q(n4494), .DIN(n4495) );
  nnd4s1 U6419 ( .Q(WX660), .DIN1(n4496), .DIN2(n4497), .DIN3(n4498), .DIN4(
        n4499) );
  nnd2s1 U6420 ( .Q(n4499), .DIN1(n3473), .DIN2(n4500) );
  nnd2s1 U6421 ( .Q(n4498), .DIN1(WX501), .DIN2(n3509) );
  nnd2s1 U6422 ( .Q(n4497), .DIN1(CRC_OUT_9_23), .DIN2(n3541) );
  nnd2s1 U6423 ( .Q(n4496), .DIN1(n3445), .DIN2(n4501) );
  hi1s1 U6424 ( .Q(n4501), .DIN(n4502) );
  nnd4s1 U6425 ( .Q(WX658), .DIN1(n4503), .DIN2(n4504), .DIN3(n4505), .DIN4(
        n4506) );
  nnd2s1 U6426 ( .Q(n4506), .DIN1(n3473), .DIN2(n4507) );
  nnd2s1 U6427 ( .Q(n4505), .DIN1(WX499), .DIN2(n3508) );
  nnd2s1 U6428 ( .Q(n4504), .DIN1(CRC_OUT_9_24), .DIN2(n3540) );
  nnd2s1 U6429 ( .Q(n4503), .DIN1(n3445), .DIN2(n4508) );
  hi1s1 U6430 ( .Q(n4508), .DIN(n4509) );
  nnd4s1 U6431 ( .Q(WX656), .DIN1(n4510), .DIN2(n4511), .DIN3(n4512), .DIN4(
        n4513) );
  nnd2s1 U6432 ( .Q(n4513), .DIN1(n3473), .DIN2(n4514) );
  nnd2s1 U6433 ( .Q(n4512), .DIN1(WX497), .DIN2(n3508) );
  nnd2s1 U6434 ( .Q(n4511), .DIN1(CRC_OUT_9_25), .DIN2(n3540) );
  nnd2s1 U6435 ( .Q(n4510), .DIN1(n3445), .DIN2(n4515) );
  hi1s1 U6436 ( .Q(n4515), .DIN(n4516) );
  nnd4s1 U6437 ( .Q(WX654), .DIN1(n4517), .DIN2(n4518), .DIN3(n4519), .DIN4(
        n4520) );
  nnd2s1 U6438 ( .Q(n4520), .DIN1(n3473), .DIN2(n4521) );
  nnd2s1 U6439 ( .Q(n4519), .DIN1(WX495), .DIN2(n3508) );
  nnd2s1 U6440 ( .Q(n4518), .DIN1(CRC_OUT_9_26), .DIN2(n3540) );
  nnd2s1 U6441 ( .Q(n4517), .DIN1(n3445), .DIN2(n4522) );
  hi1s1 U6442 ( .Q(n4522), .DIN(n4523) );
  nnd4s1 U6443 ( .Q(WX652), .DIN1(n4524), .DIN2(n4525), .DIN3(n4526), .DIN4(
        n4527) );
  nnd2s1 U6444 ( .Q(n4527), .DIN1(n3473), .DIN2(n4528) );
  nnd2s1 U6445 ( .Q(n4526), .DIN1(WX493), .DIN2(n3508) );
  nnd2s1 U6446 ( .Q(n4525), .DIN1(CRC_OUT_9_27), .DIN2(n3540) );
  nnd2s1 U6447 ( .Q(n4524), .DIN1(n3445), .DIN2(n4529) );
  hi1s1 U6448 ( .Q(n4529), .DIN(n4530) );
  nnd4s1 U6449 ( .Q(WX650), .DIN1(n4531), .DIN2(n4532), .DIN3(n4533), .DIN4(
        n4534) );
  nnd2s1 U6450 ( .Q(n4534), .DIN1(n3473), .DIN2(n4535) );
  nnd2s1 U6451 ( .Q(n4533), .DIN1(WX491), .DIN2(n3508) );
  nnd2s1 U6452 ( .Q(n4532), .DIN1(CRC_OUT_9_28), .DIN2(n3540) );
  nnd2s1 U6453 ( .Q(n4531), .DIN1(n3445), .DIN2(n4536) );
  hi1s1 U6454 ( .Q(n4536), .DIN(n4537) );
  nor2s1 U6455 ( .Q(WX6498), .DIN1(n3366), .DIN2(n4538) );
  xor2s1 U6456 ( .Q(n4538), .DIN1(WX6009), .DIN2(CRC_OUT_5_30) );
  nor2s1 U6457 ( .Q(WX6496), .DIN1(n3366), .DIN2(n4539) );
  xor2s1 U6458 ( .Q(n4539), .DIN1(WX6011), .DIN2(CRC_OUT_5_29) );
  nor2s1 U6459 ( .Q(WX6494), .DIN1(n3366), .DIN2(n4540) );
  xor2s1 U6460 ( .Q(n4540), .DIN1(WX6013), .DIN2(CRC_OUT_5_28) );
  nor2s1 U6461 ( .Q(WX6492), .DIN1(n3366), .DIN2(n4541) );
  xor2s1 U6462 ( .Q(n4541), .DIN1(WX6015), .DIN2(CRC_OUT_5_27) );
  nor2s1 U6463 ( .Q(WX6490), .DIN1(n3367), .DIN2(n4542) );
  xor2s1 U6464 ( .Q(n4542), .DIN1(WX6017), .DIN2(CRC_OUT_5_26) );
  nor2s1 U6465 ( .Q(WX6488), .DIN1(n3366), .DIN2(n4543) );
  xor2s1 U6466 ( .Q(n4543), .DIN1(WX6019), .DIN2(CRC_OUT_5_25) );
  nor2s1 U6467 ( .Q(WX6486), .DIN1(n3366), .DIN2(n4544) );
  xor2s1 U6468 ( .Q(n4544), .DIN1(WX6021), .DIN2(CRC_OUT_5_24) );
  nor2s1 U6469 ( .Q(WX6484), .DIN1(n3366), .DIN2(n4545) );
  xor2s1 U6470 ( .Q(n4545), .DIN1(WX6023), .DIN2(CRC_OUT_5_23) );
  nor2s1 U6471 ( .Q(WX6482), .DIN1(n3367), .DIN2(n4546) );
  xor2s1 U6472 ( .Q(n4546), .DIN1(WX6025), .DIN2(CRC_OUT_5_22) );
  nor2s1 U6473 ( .Q(WX6480), .DIN1(n3366), .DIN2(n4547) );
  xor2s1 U6474 ( .Q(n4547), .DIN1(WX6027), .DIN2(CRC_OUT_5_21) );
  nnd4s1 U6475 ( .Q(WX648), .DIN1(n4548), .DIN2(n4549), .DIN3(n4550), .DIN4(
        n4551) );
  nnd2s1 U6476 ( .Q(n4551), .DIN1(n3473), .DIN2(n4552) );
  nnd2s1 U6477 ( .Q(n4550), .DIN1(WX489), .DIN2(n3508) );
  nnd2s1 U6478 ( .Q(n4549), .DIN1(CRC_OUT_9_29), .DIN2(n3540) );
  nnd2s1 U6479 ( .Q(n4548), .DIN1(n3445), .DIN2(n4553) );
  hi1s1 U6480 ( .Q(n4553), .DIN(n4554) );
  nor2s1 U6481 ( .Q(WX6478), .DIN1(n3367), .DIN2(n4555) );
  xor2s1 U6482 ( .Q(n4555), .DIN1(WX6029), .DIN2(CRC_OUT_5_20) );
  nor2s1 U6483 ( .Q(WX6476), .DIN1(n3367), .DIN2(n4556) );
  xor2s1 U6484 ( .Q(n4556), .DIN1(WX6031), .DIN2(CRC_OUT_5_19) );
  nor2s1 U6485 ( .Q(WX6474), .DIN1(n3367), .DIN2(n4557) );
  xor2s1 U6486 ( .Q(n4557), .DIN1(WX6033), .DIN2(CRC_OUT_5_18) );
  nor2s1 U6487 ( .Q(WX6472), .DIN1(n3367), .DIN2(n4558) );
  xor2s1 U6488 ( .Q(n4558), .DIN1(WX6035), .DIN2(CRC_OUT_5_17) );
  nor2s1 U6489 ( .Q(WX6470), .DIN1(n3368), .DIN2(n4559) );
  xor2s1 U6490 ( .Q(n4559), .DIN1(WX6037), .DIN2(CRC_OUT_5_16) );
  nor2s1 U6491 ( .Q(WX6468), .DIN1(n3367), .DIN2(n4560) );
  xor2s1 U6492 ( .Q(n4560), .DIN1(CRC_OUT_5_15), .DIN2(n4561) );
  xor2s1 U6493 ( .Q(n4561), .DIN1(WX6039), .DIN2(CRC_OUT_5_31) );
  nor2s1 U6494 ( .Q(WX6466), .DIN1(n3367), .DIN2(n4562) );
  xor2s1 U6495 ( .Q(n4562), .DIN1(WX6041), .DIN2(CRC_OUT_5_14) );
  nor2s1 U6496 ( .Q(WX6464), .DIN1(n3367), .DIN2(n4563) );
  xor2s1 U6497 ( .Q(n4563), .DIN1(WX6043), .DIN2(CRC_OUT_5_13) );
  nor2s1 U6498 ( .Q(WX6462), .DIN1(n3367), .DIN2(n4564) );
  xor2s1 U6499 ( .Q(n4564), .DIN1(WX6045), .DIN2(CRC_OUT_5_12) );
  nor2s1 U6500 ( .Q(WX6460), .DIN1(n3368), .DIN2(n4565) );
  xor2s1 U6501 ( .Q(n4565), .DIN1(WX6047), .DIN2(CRC_OUT_5_11) );
  nnd4s1 U6502 ( .Q(WX646), .DIN1(n4566), .DIN2(n4567), .DIN3(n4568), .DIN4(
        n4569) );
  nnd2s1 U6503 ( .Q(n4569), .DIN1(n3473), .DIN2(n4570) );
  nnd2s1 U6504 ( .Q(n4568), .DIN1(WX487), .DIN2(n3508) );
  nnd2s1 U6505 ( .Q(n4567), .DIN1(CRC_OUT_9_30), .DIN2(n3540) );
  nnd2s1 U6506 ( .Q(n4566), .DIN1(n3445), .DIN2(n4571) );
  hi1s1 U6507 ( .Q(n4571), .DIN(n4572) );
  nor2s1 U6508 ( .Q(WX6458), .DIN1(n3368), .DIN2(n4573) );
  xor2s1 U6509 ( .Q(n4573), .DIN1(CRC_OUT_5_10), .DIN2(n4574) );
  xor2s1 U6510 ( .Q(n4574), .DIN1(WX6049), .DIN2(CRC_OUT_5_31) );
  nor2s1 U6511 ( .Q(WX6456), .DIN1(n3368), .DIN2(n4575) );
  xor2s1 U6512 ( .Q(n4575), .DIN1(WX6051), .DIN2(CRC_OUT_5_9) );
  nor2s1 U6513 ( .Q(WX6454), .DIN1(n3368), .DIN2(n4576) );
  xor2s1 U6514 ( .Q(n4576), .DIN1(WX6053), .DIN2(CRC_OUT_5_8) );
  nor2s1 U6515 ( .Q(WX6452), .DIN1(n3369), .DIN2(n4577) );
  xor2s1 U6516 ( .Q(n4577), .DIN1(WX6055), .DIN2(CRC_OUT_5_7) );
  nor2s1 U6517 ( .Q(WX6450), .DIN1(n3368), .DIN2(n4578) );
  xor2s1 U6518 ( .Q(n4578), .DIN1(WX6057), .DIN2(CRC_OUT_5_6) );
  nor2s1 U6519 ( .Q(WX6448), .DIN1(n3368), .DIN2(n4579) );
  xor2s1 U6520 ( .Q(n4579), .DIN1(WX6059), .DIN2(CRC_OUT_5_5) );
  nor2s1 U6521 ( .Q(WX6446), .DIN1(n3368), .DIN2(n4580) );
  xor2s1 U6522 ( .Q(n4580), .DIN1(WX6061), .DIN2(CRC_OUT_5_4) );
  nor2s1 U6523 ( .Q(WX6444), .DIN1(n3368), .DIN2(n4581) );
  xor2s1 U6524 ( .Q(n4581), .DIN1(CRC_OUT_5_3), .DIN2(n4582) );
  xor2s1 U6525 ( .Q(n4582), .DIN1(WX6063), .DIN2(CRC_OUT_5_31) );
  nor2s1 U6526 ( .Q(WX6442), .DIN1(n3368), .DIN2(n4583) );
  xor2s1 U6527 ( .Q(n4583), .DIN1(WX6065), .DIN2(CRC_OUT_5_2) );
  nor2s1 U6528 ( .Q(WX6440), .DIN1(n3369), .DIN2(n4584) );
  xor2s1 U6529 ( .Q(n4584), .DIN1(WX6067), .DIN2(CRC_OUT_5_1) );
  nnd4s1 U6530 ( .Q(WX644), .DIN1(n4585), .DIN2(n4586), .DIN3(n4587), .DIN4(
        n4588) );
  nnd2s1 U6531 ( .Q(n4588), .DIN1(n3473), .DIN2(n4589) );
  nnd2s1 U6532 ( .Q(n4587), .DIN1(WX485), .DIN2(n3508) );
  nnd2s1 U6533 ( .Q(n4586), .DIN1(CRC_OUT_9_31), .DIN2(n3540) );
  nnd2s1 U6534 ( .Q(n4585), .DIN1(n3445), .DIN2(n4590) );
  hi1s1 U6535 ( .Q(n4590), .DIN(n4591) );
  nor2s1 U6536 ( .Q(WX6438), .DIN1(n3369), .DIN2(n4592) );
  xor2s1 U6537 ( .Q(n4592), .DIN1(WX6069), .DIN2(CRC_OUT_5_0) );
  nor2s1 U6538 ( .Q(WX6436), .DIN1(n3369), .DIN2(n4593) );
  xor2s1 U6539 ( .Q(n4593), .DIN1(WX6071), .DIN2(CRC_OUT_5_31) );
  and2s1 U6540 ( .Q(WX6070), .DIN1(RESET), .DIN2(WX6007) );
  and2s1 U6541 ( .Q(WX6068), .DIN1(RESET), .DIN2(WX6005) );
  and2s1 U6542 ( .Q(WX6066), .DIN1(RESET), .DIN2(WX6003) );
  and2s1 U6543 ( .Q(WX6064), .DIN1(RESET), .DIN2(WX6001) );
  and2s1 U6544 ( .Q(WX6062), .DIN1(RESET), .DIN2(WX5999) );
  and2s1 U6545 ( .Q(WX6060), .DIN1(RESET), .DIN2(WX5997) );
  and2s1 U6546 ( .Q(WX6058), .DIN1(RESET), .DIN2(WX5995) );
  and2s1 U6547 ( .Q(WX6056), .DIN1(RESET), .DIN2(WX5993) );
  and2s1 U6548 ( .Q(WX6054), .DIN1(RESET), .DIN2(WX5991) );
  and2s1 U6549 ( .Q(WX6052), .DIN1(RESET), .DIN2(WX5989) );
  and2s1 U6550 ( .Q(WX6050), .DIN1(RESET), .DIN2(WX5987) );
  and2s1 U6551 ( .Q(WX6048), .DIN1(RESET), .DIN2(WX5985) );
  and2s1 U6552 ( .Q(WX6046), .DIN1(RESET), .DIN2(WX5983) );
  and2s1 U6553 ( .Q(WX6044), .DIN1(RESET), .DIN2(WX5981) );
  and2s1 U6554 ( .Q(WX6042), .DIN1(RESET), .DIN2(WX5979) );
  and2s1 U6555 ( .Q(WX6040), .DIN1(RESET), .DIN2(WX5977) );
  and2s1 U6556 ( .Q(WX6038), .DIN1(RESET), .DIN2(WX5975) );
  and2s1 U6557 ( .Q(WX6036), .DIN1(RESET), .DIN2(WX5973) );
  and2s1 U6558 ( .Q(WX6034), .DIN1(RESET), .DIN2(WX5971) );
  and2s1 U6559 ( .Q(WX6032), .DIN1(RESET), .DIN2(WX5969) );
  and2s1 U6560 ( .Q(WX6030), .DIN1(RESET), .DIN2(WX5967) );
  and2s1 U6561 ( .Q(WX6028), .DIN1(RESET), .DIN2(WX5965) );
  and2s1 U6562 ( .Q(WX6026), .DIN1(RESET), .DIN2(WX5963) );
  and2s1 U6563 ( .Q(WX6024), .DIN1(RESET), .DIN2(WX5961) );
  and2s1 U6564 ( .Q(WX6022), .DIN1(RESET), .DIN2(WX5959) );
  and2s1 U6565 ( .Q(WX6020), .DIN1(RESET), .DIN2(WX5957) );
  and2s1 U6566 ( .Q(WX6018), .DIN1(RESET), .DIN2(WX5955) );
  and2s1 U6567 ( .Q(WX6016), .DIN1(RESET), .DIN2(WX5953) );
  and2s1 U6568 ( .Q(WX6014), .DIN1(RESET), .DIN2(WX5951) );
  and2s1 U6569 ( .Q(WX6012), .DIN1(RESET), .DIN2(WX5949) );
  and2s1 U6570 ( .Q(WX6010), .DIN1(RESET), .DIN2(WX5947) );
  and2s1 U6571 ( .Q(WX6008), .DIN1(RESET), .DIN2(WX5945) );
  and2s1 U6572 ( .Q(WX6006), .DIN1(RESET), .DIN2(WX5943) );
  and2s1 U6573 ( .Q(WX6004), .DIN1(RESET), .DIN2(WX5941) );
  and2s1 U6574 ( .Q(WX6002), .DIN1(RESET), .DIN2(WX5939) );
  and2s1 U6575 ( .Q(WX6000), .DIN1(RESET), .DIN2(WX5937) );
  and2s1 U6576 ( .Q(WX5998), .DIN1(RESET), .DIN2(WX5935) );
  and2s1 U6577 ( .Q(WX5996), .DIN1(RESET), .DIN2(WX5933) );
  and2s1 U6578 ( .Q(WX5994), .DIN1(RESET), .DIN2(WX5931) );
  and2s1 U6579 ( .Q(WX5992), .DIN1(RESET), .DIN2(WX5929) );
  and2s1 U6580 ( .Q(WX5990), .DIN1(RESET), .DIN2(WX5927) );
  and2s1 U6581 ( .Q(WX5988), .DIN1(RESET), .DIN2(WX5925) );
  and2s1 U6582 ( .Q(WX5986), .DIN1(RESET), .DIN2(WX5923) );
  and2s1 U6583 ( .Q(WX5984), .DIN1(RESET), .DIN2(WX5921) );
  and2s1 U6584 ( .Q(WX5982), .DIN1(RESET), .DIN2(WX5919) );
  and2s1 U6585 ( .Q(WX5980), .DIN1(RESET), .DIN2(WX5917) );
  and2s1 U6586 ( .Q(WX5978), .DIN1(RESET), .DIN2(WX5915) );
  and2s1 U6587 ( .Q(WX5976), .DIN1(RESET), .DIN2(WX5913) );
  nor2s1 U6588 ( .Q(WX5974), .DIN1(n3369), .DIN2(n2997) );
  nor2s1 U6589 ( .Q(WX5972), .DIN1(n3369), .DIN2(n2998) );
  nor2s1 U6590 ( .Q(WX5970), .DIN1(n3369), .DIN2(n2999) );
  nor2s1 U6591 ( .Q(WX5968), .DIN1(n3369), .DIN2(n3000) );
  nor2s1 U6592 ( .Q(WX5966), .DIN1(n3369), .DIN2(n3001) );
  nor2s1 U6593 ( .Q(WX5964), .DIN1(n3369), .DIN2(n3002) );
  nor2s1 U6594 ( .Q(WX5962), .DIN1(n3370), .DIN2(n3003) );
  nor2s1 U6595 ( .Q(WX5960), .DIN1(n3370), .DIN2(n3004) );
  nor2s1 U6596 ( .Q(WX5958), .DIN1(n3370), .DIN2(n3005) );
  nor2s1 U6597 ( .Q(WX5956), .DIN1(n3370), .DIN2(n3006) );
  nor2s1 U6598 ( .Q(WX5954), .DIN1(n3370), .DIN2(n3007) );
  nor2s1 U6599 ( .Q(WX5952), .DIN1(n3370), .DIN2(n3008) );
  nor2s1 U6600 ( .Q(WX5950), .DIN1(n3370), .DIN2(n3009) );
  nor2s1 U6601 ( .Q(WX5948), .DIN1(n3370), .DIN2(n3010) );
  nor2s1 U6602 ( .Q(WX5946), .DIN1(n3370), .DIN2(n3011) );
  nor2s1 U6603 ( .Q(WX5944), .DIN1(n3371), .DIN2(n3012) );
  nor2s1 U6604 ( .Q(WX5942), .DIN1(n3371), .DIN2(n3157) );
  nor2s1 U6605 ( .Q(WX5940), .DIN1(n3371), .DIN2(n3158) );
  nor2s1 U6606 ( .Q(WX5938), .DIN1(n3371), .DIN2(n3159) );
  nor2s1 U6607 ( .Q(WX5936), .DIN1(n3371), .DIN2(n3160) );
  nor2s1 U6608 ( .Q(WX5934), .DIN1(n3371), .DIN2(n3161) );
  nor2s1 U6609 ( .Q(WX5932), .DIN1(n3371), .DIN2(n3162) );
  nor2s1 U6610 ( .Q(WX5930), .DIN1(n3371), .DIN2(n3163) );
  nor2s1 U6611 ( .Q(WX5928), .DIN1(n3371), .DIN2(n3164) );
  nor2s1 U6612 ( .Q(WX5926), .DIN1(n3371), .DIN2(n3165) );
  nor2s1 U6613 ( .Q(WX5924), .DIN1(n3372), .DIN2(n3166) );
  nor2s1 U6614 ( .Q(WX5922), .DIN1(n3372), .DIN2(n3167) );
  nor2s1 U6615 ( .Q(WX5920), .DIN1(n3372), .DIN2(n3168) );
  nor2s1 U6616 ( .Q(WX5918), .DIN1(n3372), .DIN2(n3169) );
  nor2s1 U6617 ( .Q(WX5916), .DIN1(n3372), .DIN2(n3170) );
  nor2s1 U6618 ( .Q(WX5914), .DIN1(n3372), .DIN2(n3171) );
  nor2s1 U6619 ( .Q(WX5912), .DIN1(n3372), .DIN2(n3172) );
  and2s1 U6620 ( .Q(WX5910), .DIN1(RESET), .DIN2(WX5847) );
  and2s1 U6621 ( .Q(WX5908), .DIN1(RESET), .DIN2(WX5845) );
  and2s1 U6622 ( .Q(WX5906), .DIN1(RESET), .DIN2(WX5843) );
  and2s1 U6623 ( .Q(WX5904), .DIN1(RESET), .DIN2(WX5841) );
  and2s1 U6624 ( .Q(WX5902), .DIN1(RESET), .DIN2(WX5839) );
  and2s1 U6625 ( .Q(WX5900), .DIN1(RESET), .DIN2(WX5837) );
  and2s1 U6626 ( .Q(WX5898), .DIN1(RESET), .DIN2(WX5835) );
  and2s1 U6627 ( .Q(WX5896), .DIN1(RESET), .DIN2(WX5833) );
  and2s1 U6628 ( .Q(WX5894), .DIN1(RESET), .DIN2(WX5831) );
  and2s1 U6629 ( .Q(WX5892), .DIN1(RESET), .DIN2(WX5829) );
  and2s1 U6630 ( .Q(WX5890), .DIN1(RESET), .DIN2(WX5827) );
  and2s1 U6631 ( .Q(WX5888), .DIN1(RESET), .DIN2(WX5825) );
  and2s1 U6632 ( .Q(WX5886), .DIN1(RESET), .DIN2(WX5823) );
  and2s1 U6633 ( .Q(WX5884), .DIN1(RESET), .DIN2(WX5821) );
  and2s1 U6634 ( .Q(WX5882), .DIN1(RESET), .DIN2(WX5819) );
  and2s1 U6635 ( .Q(WX5880), .DIN1(RESET), .DIN2(WX5817) );
  nnd4s1 U6636 ( .Q(WX5878), .DIN1(n4594), .DIN2(n4595), .DIN3(n4596), .DIN4(
        n4597) );
  nnd2s1 U6637 ( .Q(n4597), .DIN1(n3473), .DIN2(n4101) );
  xor2s1 U6638 ( .Q(n4101), .DIN1(n4598), .DIN2(n4599) );
  xor2s1 U6639 ( .Q(n4599), .DIN1(WX7236), .DIN2(n3141) );
  xor2s1 U6640 ( .Q(n4598), .DIN1(n3237), .DIN2(WX7300) );
  nnd2s1 U6641 ( .Q(n4596), .DIN1(n3445), .DIN2(n4600) );
  nnd2s1 U6642 ( .Q(n4595), .DIN1(WX5719), .DIN2(n3508) );
  nnd2s1 U6643 ( .Q(n4594), .DIN1(CRC_OUT_5_0), .DIN2(n3540) );
  nnd4s1 U6644 ( .Q(WX5876), .DIN1(n4601), .DIN2(n4602), .DIN3(n4603), .DIN4(
        n4604) );
  nnd2s1 U6645 ( .Q(n4604), .DIN1(n3473), .DIN2(n4108) );
  xor2s1 U6646 ( .Q(n4108), .DIN1(n4605), .DIN2(n4606) );
  xor2s1 U6647 ( .Q(n4606), .DIN1(WX7234), .DIN2(n3142) );
  xor2s1 U6648 ( .Q(n4605), .DIN1(n3238), .DIN2(WX7298) );
  nnd2s1 U6649 ( .Q(n4603), .DIN1(n3445), .DIN2(n4607) );
  nnd2s1 U6650 ( .Q(n4602), .DIN1(WX5717), .DIN2(n3508) );
  nnd2s1 U6651 ( .Q(n4601), .DIN1(CRC_OUT_5_1), .DIN2(n3540) );
  nnd4s1 U6652 ( .Q(WX5874), .DIN1(n4608), .DIN2(n4609), .DIN3(n4610), .DIN4(
        n4611) );
  nnd2s1 U6653 ( .Q(n4611), .DIN1(n3474), .DIN2(n4115) );
  xor2s1 U6654 ( .Q(n4115), .DIN1(n4612), .DIN2(n4613) );
  xor2s1 U6655 ( .Q(n4613), .DIN1(WX7232), .DIN2(n3143) );
  xor2s1 U6656 ( .Q(n4612), .DIN1(n3239), .DIN2(WX7296) );
  nnd2s1 U6657 ( .Q(n4610), .DIN1(n3445), .DIN2(n4614) );
  nnd2s1 U6658 ( .Q(n4609), .DIN1(WX5715), .DIN2(n3508) );
  nnd2s1 U6659 ( .Q(n4608), .DIN1(CRC_OUT_5_2), .DIN2(n3540) );
  nnd4s1 U6660 ( .Q(WX5872), .DIN1(n4615), .DIN2(n4616), .DIN3(n4617), .DIN4(
        n4618) );
  nnd2s1 U6661 ( .Q(n4618), .DIN1(n3474), .DIN2(n4122) );
  xor2s1 U6662 ( .Q(n4122), .DIN1(n4619), .DIN2(n4620) );
  xor2s1 U6663 ( .Q(n4620), .DIN1(WX7230), .DIN2(n3144) );
  xor2s1 U6664 ( .Q(n4619), .DIN1(n3240), .DIN2(WX7294) );
  nnd2s1 U6665 ( .Q(n4617), .DIN1(n3445), .DIN2(n4621) );
  nnd2s1 U6666 ( .Q(n4616), .DIN1(WX5713), .DIN2(n3508) );
  nnd2s1 U6667 ( .Q(n4615), .DIN1(CRC_OUT_5_3), .DIN2(n3540) );
  nnd4s1 U6668 ( .Q(WX5870), .DIN1(n4622), .DIN2(n4623), .DIN3(n4624), .DIN4(
        n4625) );
  nnd2s1 U6669 ( .Q(n4625), .DIN1(n3474), .DIN2(n4129) );
  xor2s1 U6670 ( .Q(n4129), .DIN1(n4626), .DIN2(n4627) );
  xor2s1 U6671 ( .Q(n4627), .DIN1(WX7228), .DIN2(n3145) );
  xor2s1 U6672 ( .Q(n4626), .DIN1(n3241), .DIN2(WX7292) );
  nnd2s1 U6673 ( .Q(n4624), .DIN1(n3444), .DIN2(n4628) );
  nnd2s1 U6674 ( .Q(n4623), .DIN1(WX5711), .DIN2(n3507) );
  nnd2s1 U6675 ( .Q(n4622), .DIN1(CRC_OUT_5_4), .DIN2(n3539) );
  nnd4s1 U6676 ( .Q(WX5868), .DIN1(n4629), .DIN2(n4630), .DIN3(n4631), .DIN4(
        n4632) );
  nnd2s1 U6677 ( .Q(n4632), .DIN1(n3474), .DIN2(n4136) );
  xor2s1 U6678 ( .Q(n4136), .DIN1(n4633), .DIN2(n4634) );
  xor2s1 U6679 ( .Q(n4634), .DIN1(WX7226), .DIN2(n3146) );
  xor2s1 U6680 ( .Q(n4633), .DIN1(n3242), .DIN2(WX7290) );
  nnd2s1 U6681 ( .Q(n4631), .DIN1(n3444), .DIN2(n4635) );
  nnd2s1 U6682 ( .Q(n4630), .DIN1(WX5709), .DIN2(n3507) );
  nnd2s1 U6683 ( .Q(n4629), .DIN1(CRC_OUT_5_5), .DIN2(n3539) );
  nnd4s1 U6684 ( .Q(WX5866), .DIN1(n4636), .DIN2(n4637), .DIN3(n4638), .DIN4(
        n4639) );
  nnd2s1 U6685 ( .Q(n4639), .DIN1(n3474), .DIN2(n4143) );
  xor2s1 U6686 ( .Q(n4143), .DIN1(n4640), .DIN2(n4641) );
  xor2s1 U6687 ( .Q(n4641), .DIN1(WX7224), .DIN2(n3147) );
  xor2s1 U6688 ( .Q(n4640), .DIN1(n3243), .DIN2(WX7288) );
  nnd2s1 U6689 ( .Q(n4638), .DIN1(n3444), .DIN2(n4642) );
  nnd2s1 U6690 ( .Q(n4637), .DIN1(WX5707), .DIN2(n3507) );
  nnd2s1 U6691 ( .Q(n4636), .DIN1(CRC_OUT_5_6), .DIN2(n3539) );
  nnd4s1 U6692 ( .Q(WX5864), .DIN1(n4643), .DIN2(n4644), .DIN3(n4645), .DIN4(
        n4646) );
  nnd2s1 U6693 ( .Q(n4646), .DIN1(n3474), .DIN2(n4150) );
  xor2s1 U6694 ( .Q(n4150), .DIN1(n4647), .DIN2(n4648) );
  xor2s1 U6695 ( .Q(n4648), .DIN1(WX7222), .DIN2(n3148) );
  xor2s1 U6696 ( .Q(n4647), .DIN1(n3244), .DIN2(WX7286) );
  nnd2s1 U6697 ( .Q(n4645), .DIN1(n3444), .DIN2(n4649) );
  nnd2s1 U6698 ( .Q(n4644), .DIN1(WX5705), .DIN2(n3507) );
  nnd2s1 U6699 ( .Q(n4643), .DIN1(CRC_OUT_5_7), .DIN2(n3539) );
  nnd4s1 U6700 ( .Q(WX5862), .DIN1(n4650), .DIN2(n4651), .DIN3(n4652), .DIN4(
        n4653) );
  nnd2s1 U6701 ( .Q(n4653), .DIN1(n3474), .DIN2(n4157) );
  xor2s1 U6702 ( .Q(n4157), .DIN1(n4654), .DIN2(n4655) );
  xor2s1 U6703 ( .Q(n4655), .DIN1(WX7220), .DIN2(n3149) );
  xor2s1 U6704 ( .Q(n4654), .DIN1(n3245), .DIN2(WX7284) );
  nnd2s1 U6705 ( .Q(n4652), .DIN1(n3444), .DIN2(n4656) );
  nnd2s1 U6706 ( .Q(n4651), .DIN1(WX5703), .DIN2(n3507) );
  nnd2s1 U6707 ( .Q(n4650), .DIN1(CRC_OUT_5_8), .DIN2(n3539) );
  nnd4s1 U6708 ( .Q(WX5860), .DIN1(n4657), .DIN2(n4658), .DIN3(n4659), .DIN4(
        n4660) );
  nnd2s1 U6709 ( .Q(n4660), .DIN1(n3474), .DIN2(n4164) );
  xor2s1 U6710 ( .Q(n4164), .DIN1(n4661), .DIN2(n4662) );
  xor2s1 U6711 ( .Q(n4662), .DIN1(WX7218), .DIN2(n3150) );
  xor2s1 U6712 ( .Q(n4661), .DIN1(n3246), .DIN2(WX7282) );
  nnd2s1 U6713 ( .Q(n4659), .DIN1(n3444), .DIN2(n4663) );
  nnd2s1 U6714 ( .Q(n4658), .DIN1(WX5701), .DIN2(n3507) );
  nnd2s1 U6715 ( .Q(n4657), .DIN1(CRC_OUT_5_9), .DIN2(n3539) );
  nnd4s1 U6716 ( .Q(WX5858), .DIN1(n4664), .DIN2(n4665), .DIN3(n4666), .DIN4(
        n4667) );
  nnd2s1 U6717 ( .Q(n4667), .DIN1(n3474), .DIN2(n4171) );
  xor2s1 U6718 ( .Q(n4171), .DIN1(n4668), .DIN2(n4669) );
  xor2s1 U6719 ( .Q(n4669), .DIN1(WX7216), .DIN2(n3151) );
  xor2s1 U6720 ( .Q(n4668), .DIN1(n3247), .DIN2(WX7280) );
  nnd2s1 U6721 ( .Q(n4666), .DIN1(n3444), .DIN2(n4670) );
  nnd2s1 U6722 ( .Q(n4665), .DIN1(WX5699), .DIN2(n3507) );
  nnd2s1 U6723 ( .Q(n4664), .DIN1(CRC_OUT_5_10), .DIN2(n3539) );
  nnd4s1 U6724 ( .Q(WX5856), .DIN1(n4671), .DIN2(n4672), .DIN3(n4673), .DIN4(
        n4674) );
  nnd2s1 U6725 ( .Q(n4674), .DIN1(n3474), .DIN2(n4178) );
  xor2s1 U6726 ( .Q(n4178), .DIN1(n4675), .DIN2(n4676) );
  xor2s1 U6727 ( .Q(n4676), .DIN1(WX7214), .DIN2(n3152) );
  xor2s1 U6728 ( .Q(n4675), .DIN1(n3248), .DIN2(WX7278) );
  nnd2s1 U6729 ( .Q(n4673), .DIN1(n3444), .DIN2(n4677) );
  nnd2s1 U6730 ( .Q(n4672), .DIN1(WX5697), .DIN2(n3507) );
  nnd2s1 U6731 ( .Q(n4671), .DIN1(CRC_OUT_5_11), .DIN2(n3539) );
  nnd4s1 U6732 ( .Q(WX5854), .DIN1(n4678), .DIN2(n4679), .DIN3(n4680), .DIN4(
        n4681) );
  nnd2s1 U6733 ( .Q(n4681), .DIN1(n3474), .DIN2(n4185) );
  xor2s1 U6734 ( .Q(n4185), .DIN1(n4682), .DIN2(n4683) );
  xor2s1 U6735 ( .Q(n4683), .DIN1(WX7212), .DIN2(n3153) );
  xor2s1 U6736 ( .Q(n4682), .DIN1(n3249), .DIN2(WX7276) );
  nnd2s1 U6737 ( .Q(n4680), .DIN1(n3444), .DIN2(n4684) );
  nnd2s1 U6738 ( .Q(n4679), .DIN1(WX5695), .DIN2(n3507) );
  nnd2s1 U6739 ( .Q(n4678), .DIN1(CRC_OUT_5_12), .DIN2(n3539) );
  nnd4s1 U6740 ( .Q(WX5852), .DIN1(n4685), .DIN2(n4686), .DIN3(n4687), .DIN4(
        n4688) );
  nnd2s1 U6741 ( .Q(n4688), .DIN1(n3474), .DIN2(n4192) );
  xor2s1 U6742 ( .Q(n4192), .DIN1(n4689), .DIN2(n4690) );
  xor2s1 U6743 ( .Q(n4690), .DIN1(WX7210), .DIN2(n3154) );
  xor2s1 U6744 ( .Q(n4689), .DIN1(n3250), .DIN2(WX7274) );
  nnd2s1 U6745 ( .Q(n4687), .DIN1(n3444), .DIN2(n4691) );
  nnd2s1 U6746 ( .Q(n4686), .DIN1(WX5693), .DIN2(n3507) );
  nnd2s1 U6747 ( .Q(n4685), .DIN1(CRC_OUT_5_13), .DIN2(n3539) );
  nnd4s1 U6748 ( .Q(WX5850), .DIN1(n4692), .DIN2(n4693), .DIN3(n4694), .DIN4(
        n4695) );
  nnd2s1 U6749 ( .Q(n4695), .DIN1(n3474), .DIN2(n4199) );
  xor2s1 U6750 ( .Q(n4199), .DIN1(n4696), .DIN2(n4697) );
  xor2s1 U6751 ( .Q(n4697), .DIN1(WX7208), .DIN2(n3155) );
  xor2s1 U6752 ( .Q(n4696), .DIN1(n3251), .DIN2(WX7272) );
  nnd2s1 U6753 ( .Q(n4694), .DIN1(n3444), .DIN2(n4698) );
  nnd2s1 U6754 ( .Q(n4693), .DIN1(WX5691), .DIN2(n3507) );
  nnd2s1 U6755 ( .Q(n4692), .DIN1(CRC_OUT_5_14), .DIN2(n3539) );
  nnd4s1 U6756 ( .Q(WX5848), .DIN1(n4699), .DIN2(n4700), .DIN3(n4701), .DIN4(
        n4702) );
  nnd2s1 U6757 ( .Q(n4702), .DIN1(n3475), .DIN2(n4206) );
  xor2s1 U6758 ( .Q(n4206), .DIN1(n4703), .DIN2(n4704) );
  xor2s1 U6759 ( .Q(n4704), .DIN1(WX7206), .DIN2(n3156) );
  xor2s1 U6760 ( .Q(n4703), .DIN1(n3252), .DIN2(WX7270) );
  nnd2s1 U6761 ( .Q(n4701), .DIN1(n3444), .DIN2(n4705) );
  nnd2s1 U6762 ( .Q(n4700), .DIN1(WX5689), .DIN2(n3507) );
  nnd2s1 U6763 ( .Q(n4699), .DIN1(CRC_OUT_5_15), .DIN2(n3539) );
  nnd4s1 U6764 ( .Q(WX5846), .DIN1(n4706), .DIN2(n4707), .DIN3(n4708), .DIN4(
        n4709) );
  nnd2s1 U6765 ( .Q(n4709), .DIN1(n3475), .DIN2(n4214) );
  xor2s1 U6766 ( .Q(n4214), .DIN1(n4710), .DIN2(n4711) );
  xor2s1 U6767 ( .Q(n4711), .DIN1(n3563), .DIN2(WX7140) );
  xor2s1 U6768 ( .Q(n4710), .DIN1(n2981), .DIN2(n4712) );
  xor2s1 U6769 ( .Q(n4712), .DIN1(WX7332), .DIN2(WX7268) );
  nnd2s1 U6770 ( .Q(n4708), .DIN1(n3444), .DIN2(n4713) );
  nnd2s1 U6771 ( .Q(n4707), .DIN1(WX5687), .DIN2(n3506) );
  nnd2s1 U6772 ( .Q(n4706), .DIN1(CRC_OUT_5_16), .DIN2(n3538) );
  nnd4s1 U6773 ( .Q(WX5844), .DIN1(n4714), .DIN2(n4715), .DIN3(n4716), .DIN4(
        n4717) );
  nnd2s1 U6774 ( .Q(n4717), .DIN1(n3475), .DIN2(n4222) );
  xor2s1 U6775 ( .Q(n4222), .DIN1(n4718), .DIN2(n4719) );
  xor2s1 U6776 ( .Q(n4719), .DIN1(n3563), .DIN2(WX7138) );
  xor2s1 U6777 ( .Q(n4718), .DIN1(n2982), .DIN2(n4720) );
  xor2s1 U6778 ( .Q(n4720), .DIN1(WX7330), .DIN2(WX7266) );
  nnd2s1 U6779 ( .Q(n4716), .DIN1(n3443), .DIN2(n4721) );
  nnd2s1 U6780 ( .Q(n4715), .DIN1(WX5685), .DIN2(n3506) );
  nnd2s1 U6781 ( .Q(n4714), .DIN1(CRC_OUT_5_17), .DIN2(n3538) );
  nnd4s1 U6782 ( .Q(WX5842), .DIN1(n4722), .DIN2(n4723), .DIN3(n4724), .DIN4(
        n4725) );
  nnd2s1 U6783 ( .Q(n4725), .DIN1(n3475), .DIN2(n4230) );
  xor2s1 U6784 ( .Q(n4230), .DIN1(n4726), .DIN2(n4727) );
  xor2s1 U6785 ( .Q(n4727), .DIN1(n3563), .DIN2(WX7136) );
  xor2s1 U6786 ( .Q(n4726), .DIN1(n2983), .DIN2(n4728) );
  xor2s1 U6787 ( .Q(n4728), .DIN1(WX7328), .DIN2(WX7264) );
  nnd2s1 U6788 ( .Q(n4724), .DIN1(n3443), .DIN2(n4729) );
  nnd2s1 U6789 ( .Q(n4723), .DIN1(WX5683), .DIN2(n3506) );
  nnd2s1 U6790 ( .Q(n4722), .DIN1(CRC_OUT_5_18), .DIN2(n3538) );
  nnd4s1 U6791 ( .Q(WX5840), .DIN1(n4730), .DIN2(n4731), .DIN3(n4732), .DIN4(
        n4733) );
  nnd2s1 U6792 ( .Q(n4733), .DIN1(n3475), .DIN2(n4238) );
  xor2s1 U6793 ( .Q(n4238), .DIN1(n4734), .DIN2(n4735) );
  xor2s1 U6794 ( .Q(n4735), .DIN1(n3564), .DIN2(WX7134) );
  xor2s1 U6795 ( .Q(n4734), .DIN1(n2984), .DIN2(n4736) );
  xor2s1 U6796 ( .Q(n4736), .DIN1(WX7326), .DIN2(WX7262) );
  nnd2s1 U6797 ( .Q(n4732), .DIN1(n3443), .DIN2(n4737) );
  nnd2s1 U6798 ( .Q(n4731), .DIN1(WX5681), .DIN2(n3506) );
  nnd2s1 U6799 ( .Q(n4730), .DIN1(CRC_OUT_5_19), .DIN2(n3538) );
  nnd4s1 U6800 ( .Q(WX5838), .DIN1(n4738), .DIN2(n4739), .DIN3(n4740), .DIN4(
        n4741) );
  nnd2s1 U6801 ( .Q(n4741), .DIN1(n3475), .DIN2(n4246) );
  xor2s1 U6802 ( .Q(n4246), .DIN1(n4742), .DIN2(n4743) );
  xor2s1 U6803 ( .Q(n4743), .DIN1(n3564), .DIN2(WX7132) );
  xor2s1 U6804 ( .Q(n4742), .DIN1(n2985), .DIN2(n4744) );
  xor2s1 U6805 ( .Q(n4744), .DIN1(WX7324), .DIN2(WX7260) );
  nnd2s1 U6806 ( .Q(n4740), .DIN1(n3443), .DIN2(n4745) );
  nnd2s1 U6807 ( .Q(n4739), .DIN1(WX5679), .DIN2(n3506) );
  nnd2s1 U6808 ( .Q(n4738), .DIN1(CRC_OUT_5_20), .DIN2(n3538) );
  nnd4s1 U6809 ( .Q(WX5836), .DIN1(n4746), .DIN2(n4747), .DIN3(n4748), .DIN4(
        n4749) );
  nnd2s1 U6810 ( .Q(n4749), .DIN1(n3475), .DIN2(n4254) );
  xor2s1 U6811 ( .Q(n4254), .DIN1(n4750), .DIN2(n4751) );
  xor2s1 U6812 ( .Q(n4751), .DIN1(n3564), .DIN2(WX7130) );
  xor2s1 U6813 ( .Q(n4750), .DIN1(n2986), .DIN2(n4752) );
  xor2s1 U6814 ( .Q(n4752), .DIN1(WX7322), .DIN2(WX7258) );
  nnd2s1 U6815 ( .Q(n4748), .DIN1(n3443), .DIN2(n4753) );
  nnd2s1 U6816 ( .Q(n4747), .DIN1(WX5677), .DIN2(n3506) );
  nnd2s1 U6817 ( .Q(n4746), .DIN1(CRC_OUT_5_21), .DIN2(n3538) );
  nnd4s1 U6818 ( .Q(WX5834), .DIN1(n4754), .DIN2(n4755), .DIN3(n4756), .DIN4(
        n4757) );
  nnd2s1 U6819 ( .Q(n4757), .DIN1(n3475), .DIN2(n4262) );
  xor2s1 U6820 ( .Q(n4262), .DIN1(n4758), .DIN2(n4759) );
  xor2s1 U6821 ( .Q(n4759), .DIN1(n3564), .DIN2(WX7128) );
  xor2s1 U6822 ( .Q(n4758), .DIN1(n2987), .DIN2(n4760) );
  xor2s1 U6823 ( .Q(n4760), .DIN1(WX7320), .DIN2(WX7256) );
  nnd2s1 U6824 ( .Q(n4756), .DIN1(n3443), .DIN2(n4761) );
  nnd2s1 U6825 ( .Q(n4755), .DIN1(WX5675), .DIN2(n3506) );
  nnd2s1 U6826 ( .Q(n4754), .DIN1(CRC_OUT_5_22), .DIN2(n3538) );
  nnd4s1 U6827 ( .Q(WX5832), .DIN1(n4762), .DIN2(n4763), .DIN3(n4764), .DIN4(
        n4765) );
  nnd2s1 U6828 ( .Q(n4765), .DIN1(n3475), .DIN2(n4270) );
  xor2s1 U6829 ( .Q(n4270), .DIN1(n4766), .DIN2(n4767) );
  xor2s1 U6830 ( .Q(n4767), .DIN1(n3564), .DIN2(WX7126) );
  xor2s1 U6831 ( .Q(n4766), .DIN1(n2988), .DIN2(n4768) );
  xor2s1 U6832 ( .Q(n4768), .DIN1(WX7318), .DIN2(WX7254) );
  nnd2s1 U6833 ( .Q(n4764), .DIN1(n3443), .DIN2(n4769) );
  nnd2s1 U6834 ( .Q(n4763), .DIN1(WX5673), .DIN2(n3506) );
  nnd2s1 U6835 ( .Q(n4762), .DIN1(CRC_OUT_5_23), .DIN2(n3538) );
  nnd4s1 U6836 ( .Q(WX5830), .DIN1(n4770), .DIN2(n4771), .DIN3(n4772), .DIN4(
        n4773) );
  nnd2s1 U6837 ( .Q(n4773), .DIN1(n3475), .DIN2(n4278) );
  xor2s1 U6838 ( .Q(n4278), .DIN1(n4774), .DIN2(n4775) );
  xor2s1 U6839 ( .Q(n4775), .DIN1(n3564), .DIN2(WX7124) );
  xor2s1 U6840 ( .Q(n4774), .DIN1(n2989), .DIN2(n4776) );
  xor2s1 U6841 ( .Q(n4776), .DIN1(WX7316), .DIN2(WX7252) );
  nnd2s1 U6842 ( .Q(n4772), .DIN1(n3443), .DIN2(n4777) );
  nnd2s1 U6843 ( .Q(n4771), .DIN1(WX5671), .DIN2(n3506) );
  nnd2s1 U6844 ( .Q(n4770), .DIN1(CRC_OUT_5_24), .DIN2(n3538) );
  nnd4s1 U6845 ( .Q(WX5828), .DIN1(n4778), .DIN2(n4779), .DIN3(n4780), .DIN4(
        n4781) );
  nnd2s1 U6846 ( .Q(n4781), .DIN1(n3475), .DIN2(n4286) );
  xor2s1 U6847 ( .Q(n4286), .DIN1(n4782), .DIN2(n4783) );
  xor2s1 U6848 ( .Q(n4783), .DIN1(n3564), .DIN2(WX7122) );
  xor2s1 U6849 ( .Q(n4782), .DIN1(n2990), .DIN2(n4784) );
  xor2s1 U6850 ( .Q(n4784), .DIN1(WX7314), .DIN2(WX7250) );
  nnd2s1 U6851 ( .Q(n4780), .DIN1(n3443), .DIN2(n4785) );
  nnd2s1 U6852 ( .Q(n4779), .DIN1(WX5669), .DIN2(n3506) );
  nnd2s1 U6853 ( .Q(n4778), .DIN1(CRC_OUT_5_25), .DIN2(n3538) );
  nnd4s1 U6854 ( .Q(WX5826), .DIN1(n4786), .DIN2(n4787), .DIN3(n4788), .DIN4(
        n4789) );
  nnd2s1 U6855 ( .Q(n4789), .DIN1(n3475), .DIN2(n4294) );
  xor2s1 U6856 ( .Q(n4294), .DIN1(n4790), .DIN2(n4791) );
  xor2s1 U6857 ( .Q(n4791), .DIN1(n3565), .DIN2(WX7120) );
  xor2s1 U6858 ( .Q(n4790), .DIN1(n2991), .DIN2(n4792) );
  xor2s1 U6859 ( .Q(n4792), .DIN1(WX7312), .DIN2(WX7248) );
  nnd2s1 U6860 ( .Q(n4788), .DIN1(n3443), .DIN2(n4793) );
  nnd2s1 U6861 ( .Q(n4787), .DIN1(WX5667), .DIN2(n3506) );
  nnd2s1 U6862 ( .Q(n4786), .DIN1(CRC_OUT_5_26), .DIN2(n3538) );
  nnd4s1 U6863 ( .Q(WX5824), .DIN1(n4794), .DIN2(n4795), .DIN3(n4796), .DIN4(
        n4797) );
  nnd2s1 U6864 ( .Q(n4797), .DIN1(n3475), .DIN2(n4302) );
  xor2s1 U6865 ( .Q(n4302), .DIN1(n4798), .DIN2(n4799) );
  xor2s1 U6866 ( .Q(n4799), .DIN1(n3565), .DIN2(WX7118) );
  xor2s1 U6867 ( .Q(n4798), .DIN1(n2992), .DIN2(n4800) );
  xor2s1 U6868 ( .Q(n4800), .DIN1(WX7310), .DIN2(WX7246) );
  nnd2s1 U6869 ( .Q(n4796), .DIN1(n3443), .DIN2(n4801) );
  nnd2s1 U6870 ( .Q(n4795), .DIN1(WX5665), .DIN2(n3506) );
  nnd2s1 U6871 ( .Q(n4794), .DIN1(CRC_OUT_5_27), .DIN2(n3538) );
  nnd4s1 U6872 ( .Q(WX5822), .DIN1(n4802), .DIN2(n4803), .DIN3(n4804), .DIN4(
        n4805) );
  nnd2s1 U6873 ( .Q(n4805), .DIN1(n3476), .DIN2(n4310) );
  xor2s1 U6874 ( .Q(n4310), .DIN1(n4806), .DIN2(n4807) );
  xor2s1 U6875 ( .Q(n4807), .DIN1(n3565), .DIN2(WX7116) );
  xor2s1 U6876 ( .Q(n4806), .DIN1(n2993), .DIN2(n4808) );
  xor2s1 U6877 ( .Q(n4808), .DIN1(WX7308), .DIN2(WX7244) );
  nnd2s1 U6878 ( .Q(n4804), .DIN1(n3443), .DIN2(n4809) );
  nnd2s1 U6879 ( .Q(n4803), .DIN1(WX5663), .DIN2(n3505) );
  nnd2s1 U6880 ( .Q(n4802), .DIN1(CRC_OUT_5_28), .DIN2(n3537) );
  nnd4s1 U6881 ( .Q(WX5820), .DIN1(n4810), .DIN2(n4811), .DIN3(n4812), .DIN4(
        n4813) );
  nnd2s1 U6882 ( .Q(n4813), .DIN1(n3476), .DIN2(n4318) );
  xor2s1 U6883 ( .Q(n4318), .DIN1(n4814), .DIN2(n4815) );
  xor2s1 U6884 ( .Q(n4815), .DIN1(n3565), .DIN2(WX7114) );
  xor2s1 U6885 ( .Q(n4814), .DIN1(n2994), .DIN2(n4816) );
  xor2s1 U6886 ( .Q(n4816), .DIN1(WX7306), .DIN2(WX7242) );
  nnd2s1 U6887 ( .Q(n4812), .DIN1(n3443), .DIN2(n4817) );
  nnd2s1 U6888 ( .Q(n4811), .DIN1(WX5661), .DIN2(n3505) );
  nnd2s1 U6889 ( .Q(n4810), .DIN1(CRC_OUT_5_29), .DIN2(n3537) );
  nnd4s1 U6890 ( .Q(WX5818), .DIN1(n4818), .DIN2(n4819), .DIN3(n4820), .DIN4(
        n4821) );
  nnd2s1 U6891 ( .Q(n4821), .DIN1(n3476), .DIN2(n4326) );
  xor2s1 U6892 ( .Q(n4326), .DIN1(n4822), .DIN2(n4823) );
  xor2s1 U6893 ( .Q(n4823), .DIN1(n3565), .DIN2(WX7112) );
  xor2s1 U6894 ( .Q(n4822), .DIN1(n2995), .DIN2(n4824) );
  xor2s1 U6895 ( .Q(n4824), .DIN1(WX7304), .DIN2(WX7240) );
  nnd2s1 U6896 ( .Q(n4820), .DIN1(n3442), .DIN2(n4825) );
  nnd2s1 U6897 ( .Q(n4819), .DIN1(WX5659), .DIN2(n3505) );
  nnd2s1 U6898 ( .Q(n4818), .DIN1(CRC_OUT_5_30), .DIN2(n3537) );
  nnd4s1 U6899 ( .Q(WX5816), .DIN1(n4826), .DIN2(n4827), .DIN3(n4828), .DIN4(
        n4829) );
  nnd2s1 U6900 ( .Q(n4829), .DIN1(n3476), .DIN2(n4334) );
  xor2s1 U6901 ( .Q(n4334), .DIN1(n4830), .DIN2(n4831) );
  xor2s1 U6902 ( .Q(n4831), .DIN1(n3565), .DIN2(WX7110) );
  xor2s1 U6903 ( .Q(n4830), .DIN1(n2996), .DIN2(n4832) );
  xor2s1 U6904 ( .Q(n4832), .DIN1(WX7302), .DIN2(WX7238) );
  nnd2s1 U6905 ( .Q(n4828), .DIN1(n3442), .DIN2(n4833) );
  nnd2s1 U6906 ( .Q(n4827), .DIN1(WX5657), .DIN2(n3505) );
  nnd2s1 U6907 ( .Q(n4826), .DIN1(CRC_OUT_5_31), .DIN2(n3537) );
  nor2s1 U6908 ( .Q(WX5718), .DIN1(WX5657), .DIN2(n3363) );
  and2s1 U6909 ( .Q(WX5716), .DIN1(RESET), .DIN2(WX5719) );
  and2s1 U6910 ( .Q(WX5714), .DIN1(RESET), .DIN2(WX5717) );
  and2s1 U6911 ( .Q(WX5712), .DIN1(RESET), .DIN2(WX5715) );
  and2s1 U6912 ( .Q(WX5710), .DIN1(RESET), .DIN2(WX5713) );
  and2s1 U6913 ( .Q(WX5708), .DIN1(RESET), .DIN2(WX5711) );
  and2s1 U6914 ( .Q(WX5706), .DIN1(RESET), .DIN2(WX5709) );
  and2s1 U6915 ( .Q(WX5704), .DIN1(RESET), .DIN2(WX5707) );
  and2s1 U6916 ( .Q(WX5702), .DIN1(RESET), .DIN2(WX5705) );
  and2s1 U6917 ( .Q(WX5700), .DIN1(RESET), .DIN2(WX5703) );
  and2s1 U6918 ( .Q(WX5698), .DIN1(RESET), .DIN2(WX5701) );
  and2s1 U6919 ( .Q(WX5696), .DIN1(RESET), .DIN2(WX5699) );
  and2s1 U6920 ( .Q(WX5694), .DIN1(RESET), .DIN2(WX5697) );
  and2s1 U6921 ( .Q(WX5692), .DIN1(RESET), .DIN2(WX5695) );
  and2s1 U6922 ( .Q(WX5690), .DIN1(RESET), .DIN2(WX5693) );
  and2s1 U6923 ( .Q(WX5688), .DIN1(RESET), .DIN2(WX5691) );
  and2s1 U6924 ( .Q(WX5686), .DIN1(RESET), .DIN2(WX5689) );
  and2s1 U6925 ( .Q(WX5684), .DIN1(RESET), .DIN2(WX5687) );
  and2s1 U6926 ( .Q(WX5682), .DIN1(RESET), .DIN2(WX5685) );
  and2s1 U6927 ( .Q(WX5680), .DIN1(RESET), .DIN2(WX5683) );
  and2s1 U6928 ( .Q(WX5678), .DIN1(RESET), .DIN2(WX5681) );
  and2s1 U6929 ( .Q(WX5676), .DIN1(RESET), .DIN2(WX5679) );
  and2s1 U6930 ( .Q(WX5674), .DIN1(RESET), .DIN2(WX5677) );
  and2s1 U6931 ( .Q(WX5672), .DIN1(RESET), .DIN2(WX5675) );
  and2s1 U6932 ( .Q(WX5670), .DIN1(RESET), .DIN2(WX5673) );
  and2s1 U6933 ( .Q(WX5668), .DIN1(RESET), .DIN2(WX5671) );
  and2s1 U6934 ( .Q(WX5666), .DIN1(RESET), .DIN2(WX5669) );
  and2s1 U6935 ( .Q(WX5664), .DIN1(RESET), .DIN2(WX5667) );
  and2s1 U6936 ( .Q(WX5662), .DIN1(RESET), .DIN2(WX5665) );
  and2s1 U6937 ( .Q(WX5660), .DIN1(RESET), .DIN2(WX5663) );
  and2s1 U6938 ( .Q(WX5658), .DIN1(RESET), .DIN2(WX5661) );
  and2s1 U6939 ( .Q(WX5656), .DIN1(RESET), .DIN2(WX5659) );
  nor2s1 U6940 ( .Q(WX546), .DIN1(WX485), .DIN2(n3363) );
  and2s1 U6941 ( .Q(WX544), .DIN1(RESET), .DIN2(WX547) );
  and2s1 U6942 ( .Q(WX542), .DIN1(RESET), .DIN2(WX545) );
  and2s1 U6943 ( .Q(WX540), .DIN1(RESET), .DIN2(WX543) );
  and2s1 U6944 ( .Q(WX538), .DIN1(RESET), .DIN2(WX541) );
  and2s1 U6945 ( .Q(WX536), .DIN1(RESET), .DIN2(WX539) );
  and2s1 U6946 ( .Q(WX534), .DIN1(RESET), .DIN2(WX537) );
  and2s1 U6947 ( .Q(WX532), .DIN1(RESET), .DIN2(WX535) );
  and2s1 U6948 ( .Q(WX530), .DIN1(RESET), .DIN2(WX533) );
  and2s1 U6949 ( .Q(WX528), .DIN1(RESET), .DIN2(WX531) );
  and2s1 U6950 ( .Q(WX526), .DIN1(RESET), .DIN2(WX529) );
  and2s1 U6951 ( .Q(WX524), .DIN1(RESET), .DIN2(WX527) );
  and2s1 U6952 ( .Q(WX522), .DIN1(RESET), .DIN2(WX525) );
  nor2s1 U6953 ( .Q(WX5205), .DIN1(n3372), .DIN2(n4834) );
  xor2s1 U6954 ( .Q(n4834), .DIN1(WX4716), .DIN2(CRC_OUT_6_30) );
  nor2s1 U6955 ( .Q(WX5203), .DIN1(n3372), .DIN2(n4835) );
  xor2s1 U6956 ( .Q(n4835), .DIN1(WX4718), .DIN2(CRC_OUT_6_29) );
  nor2s1 U6957 ( .Q(WX5201), .DIN1(n3372), .DIN2(n4836) );
  xor2s1 U6958 ( .Q(n4836), .DIN1(WX4720), .DIN2(CRC_OUT_6_28) );
  and2s1 U6959 ( .Q(WX520), .DIN1(RESET), .DIN2(WX523) );
  nor2s1 U6960 ( .Q(WX5199), .DIN1(n3373), .DIN2(n4837) );
  xor2s1 U6961 ( .Q(n4837), .DIN1(WX4722), .DIN2(CRC_OUT_6_27) );
  nor2s1 U6962 ( .Q(WX5197), .DIN1(n3373), .DIN2(n4838) );
  xor2s1 U6963 ( .Q(n4838), .DIN1(WX4724), .DIN2(CRC_OUT_6_26) );
  nor2s1 U6964 ( .Q(WX5195), .DIN1(n3373), .DIN2(n4839) );
  xor2s1 U6965 ( .Q(n4839), .DIN1(WX4726), .DIN2(CRC_OUT_6_25) );
  nor2s1 U6966 ( .Q(WX5193), .DIN1(n3373), .DIN2(n4840) );
  xor2s1 U6967 ( .Q(n4840), .DIN1(WX4728), .DIN2(CRC_OUT_6_24) );
  nor2s1 U6968 ( .Q(WX5191), .DIN1(n3373), .DIN2(n4841) );
  xor2s1 U6969 ( .Q(n4841), .DIN1(WX4730), .DIN2(CRC_OUT_6_23) );
  nor2s1 U6970 ( .Q(WX5189), .DIN1(n3373), .DIN2(n4842) );
  xor2s1 U6971 ( .Q(n4842), .DIN1(WX4732), .DIN2(CRC_OUT_6_22) );
  nor2s1 U6972 ( .Q(WX5187), .DIN1(n3373), .DIN2(n4843) );
  xor2s1 U6973 ( .Q(n4843), .DIN1(WX4734), .DIN2(CRC_OUT_6_21) );
  nor2s1 U6974 ( .Q(WX5185), .DIN1(n3373), .DIN2(n4844) );
  xor2s1 U6975 ( .Q(n4844), .DIN1(WX4736), .DIN2(CRC_OUT_6_20) );
  nor2s1 U6976 ( .Q(WX5183), .DIN1(n3373), .DIN2(n4845) );
  xor2s1 U6977 ( .Q(n4845), .DIN1(WX4738), .DIN2(CRC_OUT_6_19) );
  nor2s1 U6978 ( .Q(WX5181), .DIN1(n3373), .DIN2(n4846) );
  xor2s1 U6979 ( .Q(n4846), .DIN1(WX4740), .DIN2(CRC_OUT_6_18) );
  and2s1 U6980 ( .Q(WX518), .DIN1(RESET), .DIN2(WX521) );
  nor2s1 U6981 ( .Q(WX5179), .DIN1(n3374), .DIN2(n4847) );
  xor2s1 U6982 ( .Q(n4847), .DIN1(WX4742), .DIN2(CRC_OUT_6_17) );
  nor2s1 U6983 ( .Q(WX5177), .DIN1(n3374), .DIN2(n4848) );
  xor2s1 U6984 ( .Q(n4848), .DIN1(WX4744), .DIN2(CRC_OUT_6_16) );
  nor2s1 U6985 ( .Q(WX5175), .DIN1(n3374), .DIN2(n4849) );
  xor2s1 U6986 ( .Q(n4849), .DIN1(CRC_OUT_6_15), .DIN2(n4850) );
  xor2s1 U6987 ( .Q(n4850), .DIN1(WX4746), .DIN2(CRC_OUT_6_31) );
  nor2s1 U6988 ( .Q(WX5173), .DIN1(n3374), .DIN2(n4851) );
  xor2s1 U6989 ( .Q(n4851), .DIN1(WX4748), .DIN2(CRC_OUT_6_14) );
  nor2s1 U6990 ( .Q(WX5171), .DIN1(n3374), .DIN2(n4852) );
  xor2s1 U6991 ( .Q(n4852), .DIN1(WX4750), .DIN2(CRC_OUT_6_13) );
  nor2s1 U6992 ( .Q(WX5169), .DIN1(n3374), .DIN2(n4853) );
  xor2s1 U6993 ( .Q(n4853), .DIN1(WX4752), .DIN2(CRC_OUT_6_12) );
  nor2s1 U6994 ( .Q(WX5167), .DIN1(n3374), .DIN2(n4854) );
  xor2s1 U6995 ( .Q(n4854), .DIN1(WX4754), .DIN2(CRC_OUT_6_11) );
  nor2s1 U6996 ( .Q(WX5165), .DIN1(n3374), .DIN2(n4855) );
  xor2s1 U6997 ( .Q(n4855), .DIN1(CRC_OUT_6_10), .DIN2(n4856) );
  xor2s1 U6998 ( .Q(n4856), .DIN1(WX4756), .DIN2(CRC_OUT_6_31) );
  nor2s1 U6999 ( .Q(WX5163), .DIN1(n3374), .DIN2(n4857) );
  xor2s1 U7000 ( .Q(n4857), .DIN1(WX4758), .DIN2(CRC_OUT_6_9) );
  nor2s1 U7001 ( .Q(WX5161), .DIN1(n3374), .DIN2(n4858) );
  xor2s1 U7002 ( .Q(n4858), .DIN1(WX4760), .DIN2(CRC_OUT_6_8) );
  and2s1 U7003 ( .Q(WX516), .DIN1(RESET), .DIN2(WX519) );
  nor2s1 U7004 ( .Q(WX5159), .DIN1(n3375), .DIN2(n4859) );
  xor2s1 U7005 ( .Q(n4859), .DIN1(WX4762), .DIN2(CRC_OUT_6_7) );
  nor2s1 U7006 ( .Q(WX5157), .DIN1(n3375), .DIN2(n4860) );
  xor2s1 U7007 ( .Q(n4860), .DIN1(WX4764), .DIN2(CRC_OUT_6_6) );
  nor2s1 U7008 ( .Q(WX5155), .DIN1(n3375), .DIN2(n4861) );
  xor2s1 U7009 ( .Q(n4861), .DIN1(WX4766), .DIN2(CRC_OUT_6_5) );
  nor2s1 U7010 ( .Q(WX5153), .DIN1(n3375), .DIN2(n4862) );
  xor2s1 U7011 ( .Q(n4862), .DIN1(WX4768), .DIN2(CRC_OUT_6_4) );
  nor2s1 U7012 ( .Q(WX5151), .DIN1(n3375), .DIN2(n4863) );
  xor2s1 U7013 ( .Q(n4863), .DIN1(CRC_OUT_6_3), .DIN2(n4864) );
  xor2s1 U7014 ( .Q(n4864), .DIN1(WX4770), .DIN2(CRC_OUT_6_31) );
  nor2s1 U7015 ( .Q(WX5149), .DIN1(n3375), .DIN2(n4865) );
  xor2s1 U7016 ( .Q(n4865), .DIN1(WX4772), .DIN2(CRC_OUT_6_2) );
  nor2s1 U7017 ( .Q(WX5147), .DIN1(n3375), .DIN2(n4866) );
  xor2s1 U7018 ( .Q(n4866), .DIN1(WX4774), .DIN2(CRC_OUT_6_1) );
  nor2s1 U7019 ( .Q(WX5145), .DIN1(n3375), .DIN2(n4867) );
  xor2s1 U7020 ( .Q(n4867), .DIN1(WX4776), .DIN2(CRC_OUT_6_0) );
  nor2s1 U7021 ( .Q(WX5143), .DIN1(n3375), .DIN2(n4868) );
  xor2s1 U7022 ( .Q(n4868), .DIN1(WX4778), .DIN2(CRC_OUT_6_31) );
  and2s1 U7023 ( .Q(WX514), .DIN1(RESET), .DIN2(WX517) );
  and2s1 U7024 ( .Q(WX512), .DIN1(RESET), .DIN2(WX515) );
  and2s1 U7025 ( .Q(WX510), .DIN1(RESET), .DIN2(WX513) );
  and2s1 U7026 ( .Q(WX508), .DIN1(RESET), .DIN2(WX511) );
  and2s1 U7027 ( .Q(WX506), .DIN1(RESET), .DIN2(WX509) );
  and2s1 U7028 ( .Q(WX504), .DIN1(RESET), .DIN2(WX507) );
  and2s1 U7029 ( .Q(WX502), .DIN1(RESET), .DIN2(WX505) );
  and2s1 U7030 ( .Q(WX500), .DIN1(RESET), .DIN2(WX503) );
  and2s1 U7031 ( .Q(WX498), .DIN1(RESET), .DIN2(WX501) );
  and2s1 U7032 ( .Q(WX496), .DIN1(RESET), .DIN2(WX499) );
  and2s1 U7033 ( .Q(WX494), .DIN1(RESET), .DIN2(WX497) );
  and2s1 U7034 ( .Q(WX492), .DIN1(RESET), .DIN2(WX495) );
  and2s1 U7035 ( .Q(WX490), .DIN1(RESET), .DIN2(WX493) );
  and2s1 U7036 ( .Q(WX488), .DIN1(RESET), .DIN2(WX491) );
  and2s1 U7037 ( .Q(WX486), .DIN1(RESET), .DIN2(WX489) );
  and2s1 U7038 ( .Q(WX484), .DIN1(RESET), .DIN2(WX487) );
  and2s1 U7039 ( .Q(WX4777), .DIN1(RESET), .DIN2(WX4714) );
  and2s1 U7040 ( .Q(WX4775), .DIN1(RESET), .DIN2(WX4712) );
  and2s1 U7041 ( .Q(WX4773), .DIN1(RESET), .DIN2(WX4710) );
  and2s1 U7042 ( .Q(WX4771), .DIN1(RESET), .DIN2(WX4708) );
  and2s1 U7043 ( .Q(WX4769), .DIN1(RESET), .DIN2(WX4706) );
  and2s1 U7044 ( .Q(WX4767), .DIN1(RESET), .DIN2(WX4704) );
  and2s1 U7045 ( .Q(WX4765), .DIN1(RESET), .DIN2(WX4702) );
  and2s1 U7046 ( .Q(WX4763), .DIN1(RESET), .DIN2(WX4700) );
  and2s1 U7047 ( .Q(WX4761), .DIN1(RESET), .DIN2(WX4698) );
  and2s1 U7048 ( .Q(WX4759), .DIN1(RESET), .DIN2(WX4696) );
  and2s1 U7049 ( .Q(WX4757), .DIN1(RESET), .DIN2(WX4694) );
  and2s1 U7050 ( .Q(WX4755), .DIN1(RESET), .DIN2(WX4692) );
  and2s1 U7051 ( .Q(WX4753), .DIN1(RESET), .DIN2(WX4690) );
  and2s1 U7052 ( .Q(WX4751), .DIN1(RESET), .DIN2(WX4688) );
  and2s1 U7053 ( .Q(WX4749), .DIN1(RESET), .DIN2(WX4686) );
  and2s1 U7054 ( .Q(WX4747), .DIN1(RESET), .DIN2(WX4684) );
  and2s1 U7055 ( .Q(WX4745), .DIN1(RESET), .DIN2(WX4682) );
  and2s1 U7056 ( .Q(WX4743), .DIN1(RESET), .DIN2(WX4680) );
  and2s1 U7057 ( .Q(WX4741), .DIN1(RESET), .DIN2(WX4678) );
  and2s1 U7058 ( .Q(WX4739), .DIN1(RESET), .DIN2(WX4676) );
  and2s1 U7059 ( .Q(WX4737), .DIN1(RESET), .DIN2(WX4674) );
  and2s1 U7060 ( .Q(WX4735), .DIN1(RESET), .DIN2(WX4672) );
  and2s1 U7061 ( .Q(WX4733), .DIN1(RESET), .DIN2(WX4670) );
  and2s1 U7062 ( .Q(WX4731), .DIN1(RESET), .DIN2(WX4668) );
  and2s1 U7063 ( .Q(WX4729), .DIN1(RESET), .DIN2(WX4666) );
  and2s1 U7064 ( .Q(WX4727), .DIN1(RESET), .DIN2(WX4664) );
  and2s1 U7065 ( .Q(WX4725), .DIN1(RESET), .DIN2(WX4662) );
  and2s1 U7066 ( .Q(WX4723), .DIN1(RESET), .DIN2(WX4660) );
  and2s1 U7067 ( .Q(WX4721), .DIN1(RESET), .DIN2(WX4658) );
  and2s1 U7068 ( .Q(WX4719), .DIN1(RESET), .DIN2(WX4656) );
  and2s1 U7069 ( .Q(WX4717), .DIN1(RESET), .DIN2(WX4654) );
  and2s1 U7070 ( .Q(WX4715), .DIN1(RESET), .DIN2(WX4652) );
  and2s1 U7071 ( .Q(WX4713), .DIN1(RESET), .DIN2(WX4650) );
  and2s1 U7072 ( .Q(WX4711), .DIN1(RESET), .DIN2(WX4648) );
  and2s1 U7073 ( .Q(WX4709), .DIN1(RESET), .DIN2(WX4646) );
  and2s1 U7074 ( .Q(WX4707), .DIN1(RESET), .DIN2(WX4644) );
  and2s1 U7075 ( .Q(WX4705), .DIN1(RESET), .DIN2(WX4642) );
  and2s1 U7076 ( .Q(WX4703), .DIN1(RESET), .DIN2(WX4640) );
  and2s1 U7077 ( .Q(WX4701), .DIN1(RESET), .DIN2(WX4638) );
  and2s1 U7078 ( .Q(WX4699), .DIN1(RESET), .DIN2(WX4636) );
  and2s1 U7079 ( .Q(WX4697), .DIN1(RESET), .DIN2(WX4634) );
  and2s1 U7080 ( .Q(WX4695), .DIN1(RESET), .DIN2(WX4632) );
  and2s1 U7081 ( .Q(WX4693), .DIN1(RESET), .DIN2(WX4630) );
  and2s1 U7082 ( .Q(WX4691), .DIN1(RESET), .DIN2(WX4628) );
  and2s1 U7083 ( .Q(WX4689), .DIN1(RESET), .DIN2(WX4626) );
  and2s1 U7084 ( .Q(WX4687), .DIN1(RESET), .DIN2(WX4624) );
  and2s1 U7085 ( .Q(WX4685), .DIN1(RESET), .DIN2(WX4622) );
  and2s1 U7086 ( .Q(WX4683), .DIN1(RESET), .DIN2(WX4620) );
  nor2s1 U7087 ( .Q(WX4681), .DIN1(n3375), .DIN2(n3013) );
  nor2s1 U7088 ( .Q(WX4679), .DIN1(n3376), .DIN2(n3014) );
  nor2s1 U7089 ( .Q(WX4677), .DIN1(n3376), .DIN2(n3015) );
  nor2s1 U7090 ( .Q(WX4675), .DIN1(n3376), .DIN2(n3016) );
  nor2s1 U7091 ( .Q(WX4673), .DIN1(n3376), .DIN2(n3017) );
  nor2s1 U7092 ( .Q(WX4671), .DIN1(n3376), .DIN2(n3018) );
  nor2s1 U7093 ( .Q(WX4669), .DIN1(n3376), .DIN2(n3019) );
  nor2s1 U7094 ( .Q(WX4667), .DIN1(n3376), .DIN2(n3020) );
  nor2s1 U7095 ( .Q(WX4665), .DIN1(n3376), .DIN2(n3021) );
  nor2s1 U7096 ( .Q(WX4663), .DIN1(n3376), .DIN2(n3022) );
  nor2s1 U7097 ( .Q(WX4661), .DIN1(n3376), .DIN2(n3023) );
  nor2s1 U7098 ( .Q(WX4659), .DIN1(n3377), .DIN2(n3024) );
  nor2s1 U7099 ( .Q(WX4657), .DIN1(n3377), .DIN2(n3025) );
  nor2s1 U7100 ( .Q(WX4655), .DIN1(n3411), .DIN2(n3026) );
  nor2s1 U7101 ( .Q(WX4653), .DIN1(n3404), .DIN2(n3027) );
  nor2s1 U7102 ( .Q(WX4651), .DIN1(n3404), .DIN2(n3028) );
  nor2s1 U7103 ( .Q(WX4649), .DIN1(n3404), .DIN2(n3173) );
  nor2s1 U7104 ( .Q(WX4647), .DIN1(n3404), .DIN2(n3174) );
  nor2s1 U7105 ( .Q(WX4645), .DIN1(n3405), .DIN2(n3175) );
  nor2s1 U7106 ( .Q(WX4643), .DIN1(n3405), .DIN2(n3176) );
  nor2s1 U7107 ( .Q(WX4641), .DIN1(n3405), .DIN2(n3177) );
  nor2s1 U7108 ( .Q(WX4639), .DIN1(n3405), .DIN2(n3178) );
  nor2s1 U7109 ( .Q(WX4637), .DIN1(n3405), .DIN2(n3179) );
  nor2s1 U7110 ( .Q(WX4635), .DIN1(n3405), .DIN2(n3180) );
  nor2s1 U7111 ( .Q(WX4633), .DIN1(n3405), .DIN2(n3181) );
  nor2s1 U7112 ( .Q(WX4631), .DIN1(n3405), .DIN2(n3182) );
  nor2s1 U7113 ( .Q(WX4629), .DIN1(n3405), .DIN2(n3183) );
  nor2s1 U7114 ( .Q(WX4627), .DIN1(n3405), .DIN2(n3184) );
  nor2s1 U7115 ( .Q(WX4625), .DIN1(n3406), .DIN2(n3185) );
  nor2s1 U7116 ( .Q(WX4623), .DIN1(n3406), .DIN2(n3186) );
  nor2s1 U7117 ( .Q(WX4621), .DIN1(n3406), .DIN2(n3187) );
  nor2s1 U7118 ( .Q(WX4619), .DIN1(n3406), .DIN2(n3188) );
  and2s1 U7119 ( .Q(WX4617), .DIN1(RESET), .DIN2(WX4554) );
  and2s1 U7120 ( .Q(WX4615), .DIN1(RESET), .DIN2(WX4552) );
  and2s1 U7121 ( .Q(WX4613), .DIN1(RESET), .DIN2(WX4550) );
  and2s1 U7122 ( .Q(WX4611), .DIN1(RESET), .DIN2(WX4548) );
  and2s1 U7123 ( .Q(WX4609), .DIN1(RESET), .DIN2(WX4546) );
  and2s1 U7124 ( .Q(WX4607), .DIN1(RESET), .DIN2(WX4544) );
  and2s1 U7125 ( .Q(WX4605), .DIN1(RESET), .DIN2(WX4542) );
  and2s1 U7126 ( .Q(WX4603), .DIN1(RESET), .DIN2(WX4540) );
  and2s1 U7127 ( .Q(WX4601), .DIN1(RESET), .DIN2(WX4538) );
  and2s1 U7128 ( .Q(WX4599), .DIN1(RESET), .DIN2(WX4536) );
  and2s1 U7129 ( .Q(WX4597), .DIN1(RESET), .DIN2(WX4534) );
  and2s1 U7130 ( .Q(WX4595), .DIN1(RESET), .DIN2(WX4532) );
  and2s1 U7131 ( .Q(WX4593), .DIN1(RESET), .DIN2(WX4530) );
  and2s1 U7132 ( .Q(WX4591), .DIN1(RESET), .DIN2(WX4528) );
  and2s1 U7133 ( .Q(WX4589), .DIN1(RESET), .DIN2(WX4526) );
  and2s1 U7134 ( .Q(WX4587), .DIN1(RESET), .DIN2(WX4524) );
  nnd4s1 U7135 ( .Q(WX4585), .DIN1(n4869), .DIN2(n4870), .DIN3(n4871), .DIN4(
        n4872) );
  nnd2s1 U7136 ( .Q(n4872), .DIN1(n3476), .DIN2(n4600) );
  xor2s1 U7137 ( .Q(n4600), .DIN1(n4873), .DIN2(n4874) );
  xor2s1 U7138 ( .Q(n4874), .DIN1(WX5943), .DIN2(n3157) );
  xor2s1 U7139 ( .Q(n4873), .DIN1(n3253), .DIN2(WX6007) );
  nnd2s1 U7140 ( .Q(n4871), .DIN1(n3442), .DIN2(n4875) );
  nnd2s1 U7141 ( .Q(n4870), .DIN1(WX4426), .DIN2(n3505) );
  nnd2s1 U7142 ( .Q(n4869), .DIN1(CRC_OUT_6_0), .DIN2(n3537) );
  nnd4s1 U7143 ( .Q(WX4583), .DIN1(n4876), .DIN2(n4877), .DIN3(n4878), .DIN4(
        n4879) );
  nnd2s1 U7144 ( .Q(n4879), .DIN1(n3476), .DIN2(n4607) );
  xor2s1 U7145 ( .Q(n4607), .DIN1(n4880), .DIN2(n4881) );
  xor2s1 U7146 ( .Q(n4881), .DIN1(WX5941), .DIN2(n3158) );
  xor2s1 U7147 ( .Q(n4880), .DIN1(n3254), .DIN2(WX6005) );
  nnd2s1 U7148 ( .Q(n4878), .DIN1(n3442), .DIN2(n4882) );
  nnd2s1 U7149 ( .Q(n4877), .DIN1(WX4424), .DIN2(n3505) );
  nnd2s1 U7150 ( .Q(n4876), .DIN1(CRC_OUT_6_1), .DIN2(n3537) );
  nnd4s1 U7151 ( .Q(WX4581), .DIN1(n4883), .DIN2(n4884), .DIN3(n4885), .DIN4(
        n4886) );
  nnd2s1 U7152 ( .Q(n4886), .DIN1(n3476), .DIN2(n4614) );
  xor2s1 U7153 ( .Q(n4614), .DIN1(n4887), .DIN2(n4888) );
  xor2s1 U7154 ( .Q(n4888), .DIN1(WX5939), .DIN2(n3159) );
  xor2s1 U7155 ( .Q(n4887), .DIN1(n3255), .DIN2(WX6003) );
  nnd2s1 U7156 ( .Q(n4885), .DIN1(n3442), .DIN2(n4889) );
  nnd2s1 U7157 ( .Q(n4884), .DIN1(WX4422), .DIN2(n3505) );
  nnd2s1 U7158 ( .Q(n4883), .DIN1(CRC_OUT_6_2), .DIN2(n3537) );
  nnd4s1 U7159 ( .Q(WX4579), .DIN1(n4890), .DIN2(n4891), .DIN3(n4892), .DIN4(
        n4893) );
  nnd2s1 U7160 ( .Q(n4893), .DIN1(n3476), .DIN2(n4621) );
  xor2s1 U7161 ( .Q(n4621), .DIN1(n4894), .DIN2(n4895) );
  xor2s1 U7162 ( .Q(n4895), .DIN1(WX5937), .DIN2(n3160) );
  xor2s1 U7163 ( .Q(n4894), .DIN1(n3256), .DIN2(WX6001) );
  nnd2s1 U7164 ( .Q(n4892), .DIN1(n3442), .DIN2(n4896) );
  nnd2s1 U7165 ( .Q(n4891), .DIN1(WX4420), .DIN2(n3505) );
  nnd2s1 U7166 ( .Q(n4890), .DIN1(CRC_OUT_6_3), .DIN2(n3537) );
  nnd4s1 U7167 ( .Q(WX4577), .DIN1(n4897), .DIN2(n4898), .DIN3(n4899), .DIN4(
        n4900) );
  nnd2s1 U7168 ( .Q(n4900), .DIN1(n3476), .DIN2(n4628) );
  xor2s1 U7169 ( .Q(n4628), .DIN1(n4901), .DIN2(n4902) );
  xor2s1 U7170 ( .Q(n4902), .DIN1(WX5935), .DIN2(n3161) );
  xor2s1 U7171 ( .Q(n4901), .DIN1(n3257), .DIN2(WX5999) );
  nnd2s1 U7172 ( .Q(n4899), .DIN1(n3442), .DIN2(n4903) );
  nnd2s1 U7173 ( .Q(n4898), .DIN1(WX4418), .DIN2(n3505) );
  nnd2s1 U7174 ( .Q(n4897), .DIN1(CRC_OUT_6_4), .DIN2(n3537) );
  nnd4s1 U7175 ( .Q(WX4575), .DIN1(n4904), .DIN2(n4905), .DIN3(n4906), .DIN4(
        n4907) );
  nnd2s1 U7176 ( .Q(n4907), .DIN1(n3476), .DIN2(n4635) );
  xor2s1 U7177 ( .Q(n4635), .DIN1(n4908), .DIN2(n4909) );
  xor2s1 U7178 ( .Q(n4909), .DIN1(WX5933), .DIN2(n3162) );
  xor2s1 U7179 ( .Q(n4908), .DIN1(n3258), .DIN2(WX5997) );
  nnd2s1 U7180 ( .Q(n4906), .DIN1(n3442), .DIN2(n4910) );
  nnd2s1 U7181 ( .Q(n4905), .DIN1(WX4416), .DIN2(n3505) );
  nnd2s1 U7182 ( .Q(n4904), .DIN1(CRC_OUT_6_5), .DIN2(n3537) );
  nnd4s1 U7183 ( .Q(WX4573), .DIN1(n4911), .DIN2(n4912), .DIN3(n4913), .DIN4(
        n4914) );
  nnd2s1 U7184 ( .Q(n4914), .DIN1(n3476), .DIN2(n4642) );
  xor2s1 U7185 ( .Q(n4642), .DIN1(n4915), .DIN2(n4916) );
  xor2s1 U7186 ( .Q(n4916), .DIN1(WX5931), .DIN2(n3163) );
  xor2s1 U7187 ( .Q(n4915), .DIN1(n3259), .DIN2(WX5995) );
  nnd2s1 U7188 ( .Q(n4913), .DIN1(n3442), .DIN2(n4917) );
  nnd2s1 U7189 ( .Q(n4912), .DIN1(WX4414), .DIN2(n3505) );
  nnd2s1 U7190 ( .Q(n4911), .DIN1(CRC_OUT_6_6), .DIN2(n3537) );
  nnd4s1 U7191 ( .Q(WX4571), .DIN1(n4918), .DIN2(n4919), .DIN3(n4920), .DIN4(
        n4921) );
  nnd2s1 U7192 ( .Q(n4921), .DIN1(n3476), .DIN2(n4649) );
  xor2s1 U7193 ( .Q(n4649), .DIN1(n4922), .DIN2(n4923) );
  xor2s1 U7194 ( .Q(n4923), .DIN1(WX5929), .DIN2(n3164) );
  xor2s1 U7195 ( .Q(n4922), .DIN1(n3260), .DIN2(WX5993) );
  nnd2s1 U7196 ( .Q(n4920), .DIN1(n3442), .DIN2(n4924) );
  nnd2s1 U7197 ( .Q(n4919), .DIN1(WX4412), .DIN2(n3505) );
  nnd2s1 U7198 ( .Q(n4918), .DIN1(CRC_OUT_6_7), .DIN2(n3537) );
  nnd4s1 U7199 ( .Q(WX4569), .DIN1(n4925), .DIN2(n4926), .DIN3(n4927), .DIN4(
        n4928) );
  nnd2s1 U7200 ( .Q(n4928), .DIN1(n3476), .DIN2(n4656) );
  xor2s1 U7201 ( .Q(n4656), .DIN1(n4929), .DIN2(n4930) );
  xor2s1 U7202 ( .Q(n4930), .DIN1(WX5927), .DIN2(n3165) );
  xor2s1 U7203 ( .Q(n4929), .DIN1(n3261), .DIN2(WX5991) );
  nnd2s1 U7204 ( .Q(n4927), .DIN1(n3442), .DIN2(n4931) );
  nnd2s1 U7205 ( .Q(n4926), .DIN1(WX4410), .DIN2(n3504) );
  nnd2s1 U7206 ( .Q(n4925), .DIN1(CRC_OUT_6_8), .DIN2(n3536) );
  nnd4s1 U7207 ( .Q(WX4567), .DIN1(n4932), .DIN2(n4933), .DIN3(n4934), .DIN4(
        n4935) );
  nnd2s1 U7208 ( .Q(n4935), .DIN1(n3477), .DIN2(n4663) );
  xor2s1 U7209 ( .Q(n4663), .DIN1(n4936), .DIN2(n4937) );
  xor2s1 U7210 ( .Q(n4937), .DIN1(WX5925), .DIN2(n3166) );
  xor2s1 U7211 ( .Q(n4936), .DIN1(n3262), .DIN2(WX5989) );
  nnd2s1 U7212 ( .Q(n4934), .DIN1(n3442), .DIN2(n4938) );
  nnd2s1 U7213 ( .Q(n4933), .DIN1(WX4408), .DIN2(n3504) );
  nnd2s1 U7214 ( .Q(n4932), .DIN1(CRC_OUT_6_9), .DIN2(n3536) );
  nnd4s1 U7215 ( .Q(WX4565), .DIN1(n4939), .DIN2(n4940), .DIN3(n4941), .DIN4(
        n4942) );
  nnd2s1 U7216 ( .Q(n4942), .DIN1(n3477), .DIN2(n4670) );
  xor2s1 U7217 ( .Q(n4670), .DIN1(n4943), .DIN2(n4944) );
  xor2s1 U7218 ( .Q(n4944), .DIN1(WX5923), .DIN2(n3167) );
  xor2s1 U7219 ( .Q(n4943), .DIN1(n3263), .DIN2(WX5987) );
  nnd2s1 U7220 ( .Q(n4941), .DIN1(n3442), .DIN2(n4945) );
  nnd2s1 U7221 ( .Q(n4940), .DIN1(WX4406), .DIN2(n3504) );
  nnd2s1 U7222 ( .Q(n4939), .DIN1(CRC_OUT_6_10), .DIN2(n3536) );
  nnd4s1 U7223 ( .Q(WX4563), .DIN1(n4946), .DIN2(n4947), .DIN3(n4948), .DIN4(
        n4949) );
  nnd2s1 U7224 ( .Q(n4949), .DIN1(n3477), .DIN2(n4677) );
  xor2s1 U7225 ( .Q(n4677), .DIN1(n4950), .DIN2(n4951) );
  xor2s1 U7226 ( .Q(n4951), .DIN1(WX5921), .DIN2(n3168) );
  xor2s1 U7227 ( .Q(n4950), .DIN1(n3264), .DIN2(WX5985) );
  nnd2s1 U7228 ( .Q(n4948), .DIN1(n3441), .DIN2(n4952) );
  nnd2s1 U7229 ( .Q(n4947), .DIN1(WX4404), .DIN2(n3504) );
  nnd2s1 U7230 ( .Q(n4946), .DIN1(CRC_OUT_6_11), .DIN2(n3536) );
  nnd4s1 U7231 ( .Q(WX4561), .DIN1(n4953), .DIN2(n4954), .DIN3(n4955), .DIN4(
        n4956) );
  nnd2s1 U7232 ( .Q(n4956), .DIN1(n3477), .DIN2(n4684) );
  xor2s1 U7233 ( .Q(n4684), .DIN1(n4957), .DIN2(n4958) );
  xor2s1 U7234 ( .Q(n4958), .DIN1(WX5919), .DIN2(n3169) );
  xor2s1 U7235 ( .Q(n4957), .DIN1(n3265), .DIN2(WX5983) );
  nnd2s1 U7236 ( .Q(n4955), .DIN1(n3441), .DIN2(n4959) );
  nnd2s1 U7237 ( .Q(n4954), .DIN1(WX4402), .DIN2(n3504) );
  nnd2s1 U7238 ( .Q(n4953), .DIN1(CRC_OUT_6_12), .DIN2(n3536) );
  nnd4s1 U7239 ( .Q(WX4559), .DIN1(n4960), .DIN2(n4961), .DIN3(n4962), .DIN4(
        n4963) );
  nnd2s1 U7240 ( .Q(n4963), .DIN1(n3477), .DIN2(n4691) );
  xor2s1 U7241 ( .Q(n4691), .DIN1(n4964), .DIN2(n4965) );
  xor2s1 U7242 ( .Q(n4965), .DIN1(WX5917), .DIN2(n3170) );
  xor2s1 U7243 ( .Q(n4964), .DIN1(n3266), .DIN2(WX5981) );
  nnd2s1 U7244 ( .Q(n4962), .DIN1(n3441), .DIN2(n4966) );
  nnd2s1 U7245 ( .Q(n4961), .DIN1(WX4400), .DIN2(n3504) );
  nnd2s1 U7246 ( .Q(n4960), .DIN1(CRC_OUT_6_13), .DIN2(n3536) );
  nnd4s1 U7247 ( .Q(WX4557), .DIN1(n4967), .DIN2(n4968), .DIN3(n4969), .DIN4(
        n4970) );
  nnd2s1 U7248 ( .Q(n4970), .DIN1(n3477), .DIN2(n4698) );
  xor2s1 U7249 ( .Q(n4698), .DIN1(n4971), .DIN2(n4972) );
  xor2s1 U7250 ( .Q(n4972), .DIN1(WX5915), .DIN2(n3171) );
  xor2s1 U7251 ( .Q(n4971), .DIN1(n3267), .DIN2(WX5979) );
  nnd2s1 U7252 ( .Q(n4969), .DIN1(n3441), .DIN2(n4973) );
  nnd2s1 U7253 ( .Q(n4968), .DIN1(WX4398), .DIN2(n3504) );
  nnd2s1 U7254 ( .Q(n4967), .DIN1(CRC_OUT_6_14), .DIN2(n3536) );
  nnd4s1 U7255 ( .Q(WX4555), .DIN1(n4974), .DIN2(n4975), .DIN3(n4976), .DIN4(
        n4977) );
  nnd2s1 U7256 ( .Q(n4977), .DIN1(n3477), .DIN2(n4705) );
  xor2s1 U7257 ( .Q(n4705), .DIN1(n4978), .DIN2(n4979) );
  xor2s1 U7258 ( .Q(n4979), .DIN1(WX5913), .DIN2(n3172) );
  xor2s1 U7259 ( .Q(n4978), .DIN1(n3268), .DIN2(WX5977) );
  nnd2s1 U7260 ( .Q(n4976), .DIN1(n3441), .DIN2(n4980) );
  nnd2s1 U7261 ( .Q(n4975), .DIN1(WX4396), .DIN2(n3504) );
  nnd2s1 U7262 ( .Q(n4974), .DIN1(CRC_OUT_6_15), .DIN2(n3536) );
  nnd4s1 U7263 ( .Q(WX4553), .DIN1(n4981), .DIN2(n4982), .DIN3(n4983), .DIN4(
        n4984) );
  nnd2s1 U7264 ( .Q(n4984), .DIN1(n3477), .DIN2(n4713) );
  xor2s1 U7265 ( .Q(n4713), .DIN1(n4985), .DIN2(n4986) );
  xor2s1 U7266 ( .Q(n4986), .DIN1(n3565), .DIN2(WX5847) );
  xor2s1 U7267 ( .Q(n4985), .DIN1(n2997), .DIN2(n4987) );
  xor2s1 U7268 ( .Q(n4987), .DIN1(WX6039), .DIN2(WX5975) );
  nnd2s1 U7269 ( .Q(n4983), .DIN1(n3441), .DIN2(n4988) );
  nnd2s1 U7270 ( .Q(n4982), .DIN1(WX4394), .DIN2(n3504) );
  nnd2s1 U7271 ( .Q(n4981), .DIN1(CRC_OUT_6_16), .DIN2(n3536) );
  nnd4s1 U7272 ( .Q(WX4551), .DIN1(n4989), .DIN2(n4990), .DIN3(n4991), .DIN4(
        n4992) );
  nnd2s1 U7273 ( .Q(n4992), .DIN1(n3477), .DIN2(n4721) );
  xor2s1 U7274 ( .Q(n4721), .DIN1(n4993), .DIN2(n4994) );
  xor2s1 U7275 ( .Q(n4994), .DIN1(n3566), .DIN2(WX5845) );
  xor2s1 U7276 ( .Q(n4993), .DIN1(n2998), .DIN2(n4995) );
  xor2s1 U7277 ( .Q(n4995), .DIN1(WX6037), .DIN2(WX5973) );
  nnd2s1 U7278 ( .Q(n4991), .DIN1(n3441), .DIN2(n4996) );
  nnd2s1 U7279 ( .Q(n4990), .DIN1(WX4392), .DIN2(n3504) );
  nnd2s1 U7280 ( .Q(n4989), .DIN1(CRC_OUT_6_17), .DIN2(n3536) );
  nnd4s1 U7281 ( .Q(WX4549), .DIN1(n4997), .DIN2(n4998), .DIN3(n4999), .DIN4(
        n5000) );
  nnd2s1 U7282 ( .Q(n5000), .DIN1(n3477), .DIN2(n4729) );
  xor2s1 U7283 ( .Q(n4729), .DIN1(n5001), .DIN2(n5002) );
  xor2s1 U7284 ( .Q(n5002), .DIN1(n3566), .DIN2(WX5843) );
  xor2s1 U7285 ( .Q(n5001), .DIN1(n2999), .DIN2(n5003) );
  xor2s1 U7286 ( .Q(n5003), .DIN1(WX6035), .DIN2(WX5971) );
  nnd2s1 U7287 ( .Q(n4999), .DIN1(n3441), .DIN2(n5004) );
  nnd2s1 U7288 ( .Q(n4998), .DIN1(WX4390), .DIN2(n3504) );
  nnd2s1 U7289 ( .Q(n4997), .DIN1(CRC_OUT_6_18), .DIN2(n3536) );
  nnd4s1 U7290 ( .Q(WX4547), .DIN1(n5005), .DIN2(n5006), .DIN3(n5007), .DIN4(
        n5008) );
  nnd2s1 U7291 ( .Q(n5008), .DIN1(n3477), .DIN2(n4737) );
  xor2s1 U7292 ( .Q(n4737), .DIN1(n5009), .DIN2(n5010) );
  xor2s1 U7293 ( .Q(n5010), .DIN1(n3566), .DIN2(WX5841) );
  xor2s1 U7294 ( .Q(n5009), .DIN1(n3000), .DIN2(n5011) );
  xor2s1 U7295 ( .Q(n5011), .DIN1(WX6033), .DIN2(WX5969) );
  nnd2s1 U7296 ( .Q(n5007), .DIN1(n3441), .DIN2(n5012) );
  nnd2s1 U7297 ( .Q(n5006), .DIN1(WX4388), .DIN2(n3504) );
  nnd2s1 U7298 ( .Q(n5005), .DIN1(CRC_OUT_6_19), .DIN2(n3536) );
  nnd4s1 U7299 ( .Q(WX4545), .DIN1(n5013), .DIN2(n5014), .DIN3(n5015), .DIN4(
        n5016) );
  nnd2s1 U7300 ( .Q(n5016), .DIN1(n3477), .DIN2(n4745) );
  xor2s1 U7301 ( .Q(n4745), .DIN1(n5017), .DIN2(n5018) );
  xor2s1 U7302 ( .Q(n5018), .DIN1(n3566), .DIN2(WX5839) );
  xor2s1 U7303 ( .Q(n5017), .DIN1(n3001), .DIN2(n5019) );
  xor2s1 U7304 ( .Q(n5019), .DIN1(WX6031), .DIN2(WX5967) );
  nnd2s1 U7305 ( .Q(n5015), .DIN1(n3441), .DIN2(n5020) );
  nnd2s1 U7306 ( .Q(n5014), .DIN1(WX4386), .DIN2(n3503) );
  nnd2s1 U7307 ( .Q(n5013), .DIN1(CRC_OUT_6_20), .DIN2(n3535) );
  nnd4s1 U7308 ( .Q(WX4543), .DIN1(n5021), .DIN2(n5022), .DIN3(n5023), .DIN4(
        n5024) );
  nnd2s1 U7309 ( .Q(n5024), .DIN1(n3477), .DIN2(n4753) );
  xor2s1 U7310 ( .Q(n4753), .DIN1(n5025), .DIN2(n5026) );
  xor2s1 U7311 ( .Q(n5026), .DIN1(n3566), .DIN2(WX5837) );
  xor2s1 U7312 ( .Q(n5025), .DIN1(n3002), .DIN2(n5027) );
  xor2s1 U7313 ( .Q(n5027), .DIN1(WX6029), .DIN2(WX5965) );
  nnd2s1 U7314 ( .Q(n5023), .DIN1(n3441), .DIN2(n5028) );
  nnd2s1 U7315 ( .Q(n5022), .DIN1(WX4384), .DIN2(n3503) );
  nnd2s1 U7316 ( .Q(n5021), .DIN1(CRC_OUT_6_21), .DIN2(n3535) );
  nnd4s1 U7317 ( .Q(WX4541), .DIN1(n5029), .DIN2(n5030), .DIN3(n5031), .DIN4(
        n5032) );
  nnd2s1 U7318 ( .Q(n5032), .DIN1(n3478), .DIN2(n4761) );
  xor2s1 U7319 ( .Q(n4761), .DIN1(n5033), .DIN2(n5034) );
  xor2s1 U7320 ( .Q(n5034), .DIN1(n3566), .DIN2(WX5835) );
  xor2s1 U7321 ( .Q(n5033), .DIN1(n3003), .DIN2(n5035) );
  xor2s1 U7322 ( .Q(n5035), .DIN1(WX6027), .DIN2(WX5963) );
  nnd2s1 U7323 ( .Q(n5031), .DIN1(n3441), .DIN2(n5036) );
  nnd2s1 U7324 ( .Q(n5030), .DIN1(WX4382), .DIN2(n3503) );
  nnd2s1 U7325 ( .Q(n5029), .DIN1(CRC_OUT_6_22), .DIN2(n3535) );
  nnd4s1 U7326 ( .Q(WX4539), .DIN1(n5037), .DIN2(n5038), .DIN3(n5039), .DIN4(
        n5040) );
  nnd2s1 U7327 ( .Q(n5040), .DIN1(n3478), .DIN2(n4769) );
  xor2s1 U7328 ( .Q(n4769), .DIN1(n5041), .DIN2(n5042) );
  xor2s1 U7329 ( .Q(n5042), .DIN1(n3566), .DIN2(WX5833) );
  xor2s1 U7330 ( .Q(n5041), .DIN1(n3004), .DIN2(n5043) );
  xor2s1 U7331 ( .Q(n5043), .DIN1(WX6025), .DIN2(WX5961) );
  nnd2s1 U7332 ( .Q(n5039), .DIN1(n3441), .DIN2(n5044) );
  nnd2s1 U7333 ( .Q(n5038), .DIN1(WX4380), .DIN2(n3503) );
  nnd2s1 U7334 ( .Q(n5037), .DIN1(CRC_OUT_6_23), .DIN2(n3535) );
  nnd4s1 U7335 ( .Q(WX4537), .DIN1(n5045), .DIN2(n5046), .DIN3(n5047), .DIN4(
        n5048) );
  nnd2s1 U7336 ( .Q(n5048), .DIN1(n3478), .DIN2(n4777) );
  xor2s1 U7337 ( .Q(n4777), .DIN1(n5049), .DIN2(n5050) );
  xor2s1 U7338 ( .Q(n5050), .DIN1(n3567), .DIN2(WX5831) );
  xor2s1 U7339 ( .Q(n5049), .DIN1(n3005), .DIN2(n5051) );
  xor2s1 U7340 ( .Q(n5051), .DIN1(WX6023), .DIN2(WX5959) );
  nnd2s1 U7341 ( .Q(n5047), .DIN1(n3440), .DIN2(n5052) );
  nnd2s1 U7342 ( .Q(n5046), .DIN1(WX4378), .DIN2(n3503) );
  nnd2s1 U7343 ( .Q(n5045), .DIN1(CRC_OUT_6_24), .DIN2(n3535) );
  nnd4s1 U7344 ( .Q(WX4535), .DIN1(n5053), .DIN2(n5054), .DIN3(n5055), .DIN4(
        n5056) );
  nnd2s1 U7345 ( .Q(n5056), .DIN1(n3478), .DIN2(n4785) );
  xor2s1 U7346 ( .Q(n4785), .DIN1(n5057), .DIN2(n5058) );
  xor2s1 U7347 ( .Q(n5058), .DIN1(n3567), .DIN2(WX5829) );
  xor2s1 U7348 ( .Q(n5057), .DIN1(n3006), .DIN2(n5059) );
  xor2s1 U7349 ( .Q(n5059), .DIN1(WX6021), .DIN2(WX5957) );
  nnd2s1 U7350 ( .Q(n5055), .DIN1(n3440), .DIN2(n5060) );
  nnd2s1 U7351 ( .Q(n5054), .DIN1(WX4376), .DIN2(n3503) );
  nnd2s1 U7352 ( .Q(n5053), .DIN1(CRC_OUT_6_25), .DIN2(n3535) );
  nnd4s1 U7353 ( .Q(WX4533), .DIN1(n5061), .DIN2(n5062), .DIN3(n5063), .DIN4(
        n5064) );
  nnd2s1 U7354 ( .Q(n5064), .DIN1(n3478), .DIN2(n4793) );
  xor2s1 U7355 ( .Q(n4793), .DIN1(n5065), .DIN2(n5066) );
  xor2s1 U7356 ( .Q(n5066), .DIN1(n3567), .DIN2(WX5827) );
  xor2s1 U7357 ( .Q(n5065), .DIN1(n3007), .DIN2(n5067) );
  xor2s1 U7358 ( .Q(n5067), .DIN1(WX6019), .DIN2(WX5955) );
  nnd2s1 U7359 ( .Q(n5063), .DIN1(n3440), .DIN2(n5068) );
  nnd2s1 U7360 ( .Q(n5062), .DIN1(WX4374), .DIN2(n3503) );
  nnd2s1 U7361 ( .Q(n5061), .DIN1(CRC_OUT_6_26), .DIN2(n3535) );
  nnd4s1 U7362 ( .Q(WX4531), .DIN1(n5069), .DIN2(n5070), .DIN3(n5071), .DIN4(
        n5072) );
  nnd2s1 U7363 ( .Q(n5072), .DIN1(n3478), .DIN2(n4801) );
  xor2s1 U7364 ( .Q(n4801), .DIN1(n5073), .DIN2(n5074) );
  xor2s1 U7365 ( .Q(n5074), .DIN1(n3567), .DIN2(WX5825) );
  xor2s1 U7366 ( .Q(n5073), .DIN1(n3008), .DIN2(n5075) );
  xor2s1 U7367 ( .Q(n5075), .DIN1(WX6017), .DIN2(WX5953) );
  nnd2s1 U7368 ( .Q(n5071), .DIN1(n3440), .DIN2(n5076) );
  nnd2s1 U7369 ( .Q(n5070), .DIN1(WX4372), .DIN2(n3503) );
  nnd2s1 U7370 ( .Q(n5069), .DIN1(CRC_OUT_6_27), .DIN2(n3535) );
  nnd4s1 U7371 ( .Q(WX4529), .DIN1(n5077), .DIN2(n5078), .DIN3(n5079), .DIN4(
        n5080) );
  nnd2s1 U7372 ( .Q(n5080), .DIN1(n3478), .DIN2(n4809) );
  xor2s1 U7373 ( .Q(n4809), .DIN1(n5081), .DIN2(n5082) );
  xor2s1 U7374 ( .Q(n5082), .DIN1(n3567), .DIN2(WX5823) );
  xor2s1 U7375 ( .Q(n5081), .DIN1(n3009), .DIN2(n5083) );
  xor2s1 U7376 ( .Q(n5083), .DIN1(WX6015), .DIN2(WX5951) );
  nnd2s1 U7377 ( .Q(n5079), .DIN1(n3440), .DIN2(n5084) );
  nnd2s1 U7378 ( .Q(n5078), .DIN1(WX4370), .DIN2(n3503) );
  nnd2s1 U7379 ( .Q(n5077), .DIN1(CRC_OUT_6_28), .DIN2(n3535) );
  nnd4s1 U7380 ( .Q(WX4527), .DIN1(n5085), .DIN2(n5086), .DIN3(n5087), .DIN4(
        n5088) );
  nnd2s1 U7381 ( .Q(n5088), .DIN1(n3478), .DIN2(n4817) );
  xor2s1 U7382 ( .Q(n4817), .DIN1(n5089), .DIN2(n5090) );
  xor2s1 U7383 ( .Q(n5090), .DIN1(n3567), .DIN2(WX5821) );
  xor2s1 U7384 ( .Q(n5089), .DIN1(n3010), .DIN2(n5091) );
  xor2s1 U7385 ( .Q(n5091), .DIN1(WX6013), .DIN2(WX5949) );
  nnd2s1 U7386 ( .Q(n5087), .DIN1(n3440), .DIN2(n5092) );
  nnd2s1 U7387 ( .Q(n5086), .DIN1(WX4368), .DIN2(n3503) );
  nnd2s1 U7388 ( .Q(n5085), .DIN1(CRC_OUT_6_29), .DIN2(n3535) );
  nnd4s1 U7389 ( .Q(WX4525), .DIN1(n5093), .DIN2(n5094), .DIN3(n5095), .DIN4(
        n5096) );
  nnd2s1 U7390 ( .Q(n5096), .DIN1(n3478), .DIN2(n4825) );
  xor2s1 U7391 ( .Q(n4825), .DIN1(n5097), .DIN2(n5098) );
  xor2s1 U7392 ( .Q(n5098), .DIN1(n3567), .DIN2(WX5819) );
  xor2s1 U7393 ( .Q(n5097), .DIN1(n3011), .DIN2(n5099) );
  xor2s1 U7394 ( .Q(n5099), .DIN1(WX6011), .DIN2(WX5947) );
  nnd2s1 U7395 ( .Q(n5095), .DIN1(n3440), .DIN2(n5100) );
  nnd2s1 U7396 ( .Q(n5094), .DIN1(WX4366), .DIN2(n3503) );
  nnd2s1 U7397 ( .Q(n5093), .DIN1(CRC_OUT_6_30), .DIN2(n3535) );
  nnd4s1 U7398 ( .Q(WX4523), .DIN1(n5101), .DIN2(n5102), .DIN3(n5103), .DIN4(
        n5104) );
  nnd2s1 U7399 ( .Q(n5104), .DIN1(n3478), .DIN2(n4833) );
  xor2s1 U7400 ( .Q(n4833), .DIN1(n5105), .DIN2(n5106) );
  xor2s1 U7401 ( .Q(n5106), .DIN1(n3568), .DIN2(WX5817) );
  xor2s1 U7402 ( .Q(n5105), .DIN1(n3012), .DIN2(n5107) );
  xor2s1 U7403 ( .Q(n5107), .DIN1(WX6009), .DIN2(WX5945) );
  nnd2s1 U7404 ( .Q(n5103), .DIN1(n3440), .DIN2(n5108) );
  nnd2s1 U7405 ( .Q(n5102), .DIN1(WX4364), .DIN2(n3503) );
  nnd2s1 U7406 ( .Q(n5101), .DIN1(CRC_OUT_6_31), .DIN2(n3535) );
  nor2s1 U7407 ( .Q(WX4425), .DIN1(WX4364), .DIN2(n3363) );
  and2s1 U7408 ( .Q(WX4423), .DIN1(RESET), .DIN2(WX4426) );
  and2s1 U7409 ( .Q(WX4421), .DIN1(RESET), .DIN2(WX4424) );
  and2s1 U7410 ( .Q(WX4419), .DIN1(RESET), .DIN2(WX4422) );
  and2s1 U7411 ( .Q(WX4417), .DIN1(RESET), .DIN2(WX4420) );
  and2s1 U7412 ( .Q(WX4415), .DIN1(RESET), .DIN2(WX4418) );
  and2s1 U7413 ( .Q(WX4413), .DIN1(RESET), .DIN2(WX4416) );
  and2s1 U7414 ( .Q(WX4411), .DIN1(RESET), .DIN2(WX4414) );
  and2s1 U7415 ( .Q(WX4409), .DIN1(RESET), .DIN2(WX4412) );
  and2s1 U7416 ( .Q(WX4407), .DIN1(RESET), .DIN2(WX4410) );
  and2s1 U7417 ( .Q(WX4405), .DIN1(RESET), .DIN2(WX4408) );
  and2s1 U7418 ( .Q(WX4403), .DIN1(RESET), .DIN2(WX4406) );
  and2s1 U7419 ( .Q(WX4401), .DIN1(RESET), .DIN2(WX4404) );
  and2s1 U7420 ( .Q(WX4399), .DIN1(RESET), .DIN2(WX4402) );
  and2s1 U7421 ( .Q(WX4397), .DIN1(RESET), .DIN2(WX4400) );
  and2s1 U7422 ( .Q(WX4395), .DIN1(RESET), .DIN2(WX4398) );
  and2s1 U7423 ( .Q(WX4393), .DIN1(RESET), .DIN2(WX4396) );
  and2s1 U7424 ( .Q(WX4391), .DIN1(RESET), .DIN2(WX4394) );
  and2s1 U7425 ( .Q(WX4389), .DIN1(RESET), .DIN2(WX4392) );
  and2s1 U7426 ( .Q(WX4387), .DIN1(RESET), .DIN2(WX4390) );
  and2s1 U7427 ( .Q(WX4385), .DIN1(RESET), .DIN2(WX4388) );
  and2s1 U7428 ( .Q(WX4383), .DIN1(RESET), .DIN2(WX4386) );
  and2s1 U7429 ( .Q(WX4381), .DIN1(RESET), .DIN2(WX4384) );
  and2s1 U7430 ( .Q(WX4379), .DIN1(RESET), .DIN2(WX4382) );
  and2s1 U7431 ( .Q(WX4377), .DIN1(RESET), .DIN2(WX4380) );
  and2s1 U7432 ( .Q(WX4375), .DIN1(RESET), .DIN2(WX4378) );
  and2s1 U7433 ( .Q(WX4373), .DIN1(RESET), .DIN2(WX4376) );
  and2s1 U7434 ( .Q(WX4371), .DIN1(RESET), .DIN2(WX4374) );
  and2s1 U7435 ( .Q(WX4369), .DIN1(RESET), .DIN2(WX4372) );
  and2s1 U7436 ( .Q(WX4367), .DIN1(RESET), .DIN2(WX4370) );
  and2s1 U7437 ( .Q(WX4365), .DIN1(RESET), .DIN2(WX4368) );
  and2s1 U7438 ( .Q(WX4363), .DIN1(RESET), .DIN2(WX4366) );
  nor2s1 U7439 ( .Q(WX3912), .DIN1(n3406), .DIN2(n5109) );
  xor2s1 U7440 ( .Q(n5109), .DIN1(WX3423), .DIN2(CRC_OUT_7_30) );
  nor2s1 U7441 ( .Q(WX3910), .DIN1(n3406), .DIN2(n5110) );
  xor2s1 U7442 ( .Q(n5110), .DIN1(WX3425), .DIN2(CRC_OUT_7_29) );
  nor2s1 U7443 ( .Q(WX3908), .DIN1(n3406), .DIN2(n5111) );
  xor2s1 U7444 ( .Q(n5111), .DIN1(WX3427), .DIN2(CRC_OUT_7_28) );
  nor2s1 U7445 ( .Q(WX3906), .DIN1(n3406), .DIN2(n5112) );
  xor2s1 U7446 ( .Q(n5112), .DIN1(WX3429), .DIN2(CRC_OUT_7_27) );
  nor2s1 U7447 ( .Q(WX3904), .DIN1(n3406), .DIN2(n5113) );
  xor2s1 U7448 ( .Q(n5113), .DIN1(WX3431), .DIN2(CRC_OUT_7_26) );
  nor2s1 U7449 ( .Q(WX3902), .DIN1(n3406), .DIN2(n5114) );
  xor2s1 U7450 ( .Q(n5114), .DIN1(WX3433), .DIN2(CRC_OUT_7_25) );
  nor2s1 U7451 ( .Q(WX3900), .DIN1(n3407), .DIN2(n5115) );
  xor2s1 U7452 ( .Q(n5115), .DIN1(WX3435), .DIN2(CRC_OUT_7_24) );
  nor2s1 U7453 ( .Q(WX3898), .DIN1(n3407), .DIN2(n5116) );
  xor2s1 U7454 ( .Q(n5116), .DIN1(WX3437), .DIN2(CRC_OUT_7_23) );
  nor2s1 U7455 ( .Q(WX3896), .DIN1(n3407), .DIN2(n5117) );
  xor2s1 U7456 ( .Q(n5117), .DIN1(WX3439), .DIN2(CRC_OUT_7_22) );
  nor2s1 U7457 ( .Q(WX3894), .DIN1(n3407), .DIN2(n5118) );
  xor2s1 U7458 ( .Q(n5118), .DIN1(WX3441), .DIN2(CRC_OUT_7_21) );
  nor2s1 U7459 ( .Q(WX3892), .DIN1(n3407), .DIN2(n5119) );
  xor2s1 U7460 ( .Q(n5119), .DIN1(WX3443), .DIN2(CRC_OUT_7_20) );
  nor2s1 U7461 ( .Q(WX3890), .DIN1(n3407), .DIN2(n5120) );
  xor2s1 U7462 ( .Q(n5120), .DIN1(WX3445), .DIN2(CRC_OUT_7_19) );
  nor2s1 U7463 ( .Q(WX3888), .DIN1(n3407), .DIN2(n5121) );
  xor2s1 U7464 ( .Q(n5121), .DIN1(WX3447), .DIN2(CRC_OUT_7_18) );
  nor2s1 U7465 ( .Q(WX3886), .DIN1(n3407), .DIN2(n5122) );
  xor2s1 U7466 ( .Q(n5122), .DIN1(WX3449), .DIN2(CRC_OUT_7_17) );
  nor2s1 U7467 ( .Q(WX3884), .DIN1(n3407), .DIN2(n5123) );
  xor2s1 U7468 ( .Q(n5123), .DIN1(WX3451), .DIN2(CRC_OUT_7_16) );
  nor2s1 U7469 ( .Q(WX3882), .DIN1(n3407), .DIN2(n5124) );
  xor2s1 U7470 ( .Q(n5124), .DIN1(CRC_OUT_7_15), .DIN2(n5125) );
  xor2s1 U7471 ( .Q(n5125), .DIN1(WX3453), .DIN2(CRC_OUT_7_31) );
  nor2s1 U7472 ( .Q(WX3880), .DIN1(n3408), .DIN2(n5126) );
  xor2s1 U7473 ( .Q(n5126), .DIN1(WX3455), .DIN2(CRC_OUT_7_14) );
  nor2s1 U7474 ( .Q(WX3878), .DIN1(n3408), .DIN2(n5127) );
  xor2s1 U7475 ( .Q(n5127), .DIN1(WX3457), .DIN2(CRC_OUT_7_13) );
  nor2s1 U7476 ( .Q(WX3876), .DIN1(n3408), .DIN2(n5128) );
  xor2s1 U7477 ( .Q(n5128), .DIN1(WX3459), .DIN2(CRC_OUT_7_12) );
  nor2s1 U7478 ( .Q(WX3874), .DIN1(n3408), .DIN2(n5129) );
  xor2s1 U7479 ( .Q(n5129), .DIN1(WX3461), .DIN2(CRC_OUT_7_11) );
  nor2s1 U7480 ( .Q(WX3872), .DIN1(n3408), .DIN2(n5130) );
  xor2s1 U7481 ( .Q(n5130), .DIN1(CRC_OUT_7_10), .DIN2(n5131) );
  xor2s1 U7482 ( .Q(n5131), .DIN1(WX3463), .DIN2(CRC_OUT_7_31) );
  nor2s1 U7483 ( .Q(WX3870), .DIN1(n3408), .DIN2(n5132) );
  xor2s1 U7484 ( .Q(n5132), .DIN1(WX3465), .DIN2(CRC_OUT_7_9) );
  nor2s1 U7485 ( .Q(WX3868), .DIN1(n3408), .DIN2(n5133) );
  xor2s1 U7486 ( .Q(n5133), .DIN1(WX3467), .DIN2(CRC_OUT_7_8) );
  nor2s1 U7487 ( .Q(WX3866), .DIN1(n3408), .DIN2(n5134) );
  xor2s1 U7488 ( .Q(n5134), .DIN1(WX3469), .DIN2(CRC_OUT_7_7) );
  nor2s1 U7489 ( .Q(WX3864), .DIN1(n3408), .DIN2(n5135) );
  xor2s1 U7490 ( .Q(n5135), .DIN1(WX3471), .DIN2(CRC_OUT_7_6) );
  nor2s1 U7491 ( .Q(WX3862), .DIN1(n3408), .DIN2(n5136) );
  xor2s1 U7492 ( .Q(n5136), .DIN1(WX3473), .DIN2(CRC_OUT_7_5) );
  nor2s1 U7493 ( .Q(WX3860), .DIN1(n3409), .DIN2(n5137) );
  xor2s1 U7494 ( .Q(n5137), .DIN1(WX3475), .DIN2(CRC_OUT_7_4) );
  nor2s1 U7495 ( .Q(WX3858), .DIN1(n3409), .DIN2(n5138) );
  xor2s1 U7496 ( .Q(n5138), .DIN1(CRC_OUT_7_3), .DIN2(n5139) );
  xor2s1 U7497 ( .Q(n5139), .DIN1(WX3477), .DIN2(CRC_OUT_7_31) );
  nor2s1 U7498 ( .Q(WX3856), .DIN1(n3409), .DIN2(n5140) );
  xor2s1 U7499 ( .Q(n5140), .DIN1(WX3479), .DIN2(CRC_OUT_7_2) );
  nor2s1 U7500 ( .Q(WX3854), .DIN1(n3409), .DIN2(n5141) );
  xor2s1 U7501 ( .Q(n5141), .DIN1(WX3481), .DIN2(CRC_OUT_7_1) );
  nor2s1 U7502 ( .Q(WX3852), .DIN1(n3409), .DIN2(n5142) );
  xor2s1 U7503 ( .Q(n5142), .DIN1(WX3483), .DIN2(CRC_OUT_7_0) );
  nor2s1 U7504 ( .Q(WX3850), .DIN1(n3409), .DIN2(n5143) );
  xor2s1 U7505 ( .Q(n5143), .DIN1(WX3485), .DIN2(CRC_OUT_7_31) );
  and2s1 U7506 ( .Q(WX3484), .DIN1(RESET), .DIN2(WX3421) );
  and2s1 U7507 ( .Q(WX3482), .DIN1(RESET), .DIN2(WX3419) );
  and2s1 U7508 ( .Q(WX3480), .DIN1(RESET), .DIN2(WX3417) );
  and2s1 U7509 ( .Q(WX3478), .DIN1(RESET), .DIN2(WX3415) );
  and2s1 U7510 ( .Q(WX3476), .DIN1(RESET), .DIN2(WX3413) );
  and2s1 U7511 ( .Q(WX3474), .DIN1(RESET), .DIN2(WX3411) );
  and2s1 U7512 ( .Q(WX3472), .DIN1(RESET), .DIN2(WX3409) );
  and2s1 U7513 ( .Q(WX3470), .DIN1(RESET), .DIN2(WX3407) );
  and2s1 U7514 ( .Q(WX3468), .DIN1(RESET), .DIN2(WX3405) );
  and2s1 U7515 ( .Q(WX3466), .DIN1(RESET), .DIN2(WX3403) );
  and2s1 U7516 ( .Q(WX3464), .DIN1(RESET), .DIN2(WX3401) );
  and2s1 U7517 ( .Q(WX3462), .DIN1(RESET), .DIN2(WX3399) );
  and2s1 U7518 ( .Q(WX3460), .DIN1(RESET), .DIN2(WX3397) );
  and2s1 U7519 ( .Q(WX3458), .DIN1(RESET), .DIN2(WX3395) );
  and2s1 U7520 ( .Q(WX3456), .DIN1(RESET), .DIN2(WX3393) );
  and2s1 U7521 ( .Q(WX3454), .DIN1(RESET), .DIN2(WX3391) );
  and2s1 U7522 ( .Q(WX3452), .DIN1(RESET), .DIN2(WX3389) );
  and2s1 U7523 ( .Q(WX3450), .DIN1(RESET), .DIN2(WX3387) );
  and2s1 U7524 ( .Q(WX3448), .DIN1(RESET), .DIN2(WX3385) );
  and2s1 U7525 ( .Q(WX3446), .DIN1(RESET), .DIN2(WX3383) );
  and2s1 U7526 ( .Q(WX3444), .DIN1(RESET), .DIN2(WX3381) );
  and2s1 U7527 ( .Q(WX3442), .DIN1(RESET), .DIN2(WX3379) );
  and2s1 U7528 ( .Q(WX3440), .DIN1(RESET), .DIN2(WX3377) );
  and2s1 U7529 ( .Q(WX3438), .DIN1(RESET), .DIN2(WX3375) );
  and2s1 U7530 ( .Q(WX3436), .DIN1(RESET), .DIN2(WX3373) );
  and2s1 U7531 ( .Q(WX3434), .DIN1(RESET), .DIN2(WX3371) );
  and2s1 U7532 ( .Q(WX3432), .DIN1(RESET), .DIN2(WX3369) );
  and2s1 U7533 ( .Q(WX3430), .DIN1(RESET), .DIN2(WX3367) );
  and2s1 U7534 ( .Q(WX3428), .DIN1(RESET), .DIN2(WX3365) );
  and2s1 U7535 ( .Q(WX3426), .DIN1(RESET), .DIN2(WX3363) );
  and2s1 U7536 ( .Q(WX3424), .DIN1(RESET), .DIN2(WX3361) );
  and2s1 U7537 ( .Q(WX3422), .DIN1(RESET), .DIN2(WX3359) );
  and2s1 U7538 ( .Q(WX3420), .DIN1(RESET), .DIN2(WX3357) );
  and2s1 U7539 ( .Q(WX3418), .DIN1(RESET), .DIN2(WX3355) );
  and2s1 U7540 ( .Q(WX3416), .DIN1(RESET), .DIN2(WX3353) );
  and2s1 U7541 ( .Q(WX3414), .DIN1(RESET), .DIN2(WX3351) );
  and2s1 U7542 ( .Q(WX3412), .DIN1(RESET), .DIN2(WX3349) );
  and2s1 U7543 ( .Q(WX3410), .DIN1(RESET), .DIN2(WX3347) );
  and2s1 U7544 ( .Q(WX3408), .DIN1(RESET), .DIN2(WX3345) );
  and2s1 U7545 ( .Q(WX3406), .DIN1(RESET), .DIN2(WX3343) );
  and2s1 U7546 ( .Q(WX3404), .DIN1(RESET), .DIN2(WX3341) );
  and2s1 U7547 ( .Q(WX3402), .DIN1(RESET), .DIN2(WX3339) );
  and2s1 U7548 ( .Q(WX3400), .DIN1(RESET), .DIN2(WX3337) );
  and2s1 U7549 ( .Q(WX3398), .DIN1(RESET), .DIN2(WX3335) );
  and2s1 U7550 ( .Q(WX3396), .DIN1(RESET), .DIN2(WX3333) );
  and2s1 U7551 ( .Q(WX3394), .DIN1(RESET), .DIN2(WX3331) );
  and2s1 U7552 ( .Q(WX3392), .DIN1(RESET), .DIN2(WX3329) );
  and2s1 U7553 ( .Q(WX3390), .DIN1(RESET), .DIN2(WX3327) );
  nor2s1 U7554 ( .Q(WX3388), .DIN1(n3409), .DIN2(n3045) );
  nor2s1 U7555 ( .Q(WX3386), .DIN1(n3409), .DIN2(n3047) );
  nor2s1 U7556 ( .Q(WX3384), .DIN1(n3409), .DIN2(n3049) );
  nor2s1 U7557 ( .Q(WX3382), .DIN1(n3409), .DIN2(n3051) );
  nor2s1 U7558 ( .Q(WX3380), .DIN1(n3410), .DIN2(n3053) );
  nor2s1 U7559 ( .Q(WX3378), .DIN1(n3410), .DIN2(n3055) );
  nor2s1 U7560 ( .Q(WX3376), .DIN1(n3410), .DIN2(n3057) );
  nor2s1 U7561 ( .Q(WX3374), .DIN1(n3410), .DIN2(n3059) );
  nor2s1 U7562 ( .Q(WX3372), .DIN1(n3410), .DIN2(n3061) );
  nor2s1 U7563 ( .Q(WX3370), .DIN1(n3410), .DIN2(n3063) );
  nor2s1 U7564 ( .Q(WX3368), .DIN1(n3410), .DIN2(n3065) );
  nor2s1 U7565 ( .Q(WX3366), .DIN1(n3410), .DIN2(n3067) );
  nor2s1 U7566 ( .Q(WX3364), .DIN1(n3410), .DIN2(n3069) );
  nor2s1 U7567 ( .Q(WX3362), .DIN1(n3410), .DIN2(n3071) );
  nor2s1 U7568 ( .Q(WX3360), .DIN1(n3411), .DIN2(n3073) );
  nor2s1 U7569 ( .Q(WX3358), .DIN1(n3411), .DIN2(n3075) );
  nor2s1 U7570 ( .Q(WX3356), .DIN1(n3411), .DIN2(n3189) );
  nor2s1 U7571 ( .Q(WX3354), .DIN1(n3411), .DIN2(n3190) );
  nor2s1 U7572 ( .Q(WX3352), .DIN1(n3411), .DIN2(n3191) );
  nor2s1 U7573 ( .Q(WX3350), .DIN1(n3411), .DIN2(n3192) );
  nor2s1 U7574 ( .Q(WX3348), .DIN1(n3411), .DIN2(n3193) );
  nor2s1 U7575 ( .Q(WX3346), .DIN1(n3411), .DIN2(n3194) );
  nor2s1 U7576 ( .Q(WX3344), .DIN1(n3411), .DIN2(n3195) );
  nor2s1 U7577 ( .Q(WX3342), .DIN1(n3412), .DIN2(n3196) );
  nor2s1 U7578 ( .Q(WX3340), .DIN1(n3412), .DIN2(n3197) );
  nor2s1 U7579 ( .Q(WX3338), .DIN1(n3412), .DIN2(n3198) );
  nor2s1 U7580 ( .Q(WX3336), .DIN1(n3412), .DIN2(n3199) );
  nor2s1 U7581 ( .Q(WX3334), .DIN1(n3412), .DIN2(n3200) );
  nor2s1 U7582 ( .Q(WX3332), .DIN1(n3412), .DIN2(n3201) );
  nor2s1 U7583 ( .Q(WX3330), .DIN1(n3412), .DIN2(n3202) );
  nor2s1 U7584 ( .Q(WX3328), .DIN1(n3412), .DIN2(n3203) );
  nor2s1 U7585 ( .Q(WX3326), .DIN1(n3412), .DIN2(n3204) );
  and2s1 U7586 ( .Q(WX3324), .DIN1(RESET), .DIN2(WX3261) );
  and2s1 U7587 ( .Q(WX3322), .DIN1(RESET), .DIN2(WX3259) );
  and2s1 U7588 ( .Q(WX3320), .DIN1(RESET), .DIN2(WX3257) );
  and2s1 U7589 ( .Q(WX3318), .DIN1(RESET), .DIN2(WX3255) );
  and2s1 U7590 ( .Q(WX3316), .DIN1(RESET), .DIN2(WX3253) );
  and2s1 U7591 ( .Q(WX3314), .DIN1(RESET), .DIN2(WX3251) );
  and2s1 U7592 ( .Q(WX3312), .DIN1(RESET), .DIN2(WX3249) );
  and2s1 U7593 ( .Q(WX3310), .DIN1(RESET), .DIN2(WX3247) );
  and2s1 U7594 ( .Q(WX3308), .DIN1(RESET), .DIN2(WX3245) );
  and2s1 U7595 ( .Q(WX3306), .DIN1(RESET), .DIN2(WX3243) );
  and2s1 U7596 ( .Q(WX3304), .DIN1(RESET), .DIN2(WX3241) );
  and2s1 U7597 ( .Q(WX3302), .DIN1(RESET), .DIN2(WX3239) );
  and2s1 U7598 ( .Q(WX3300), .DIN1(RESET), .DIN2(WX3237) );
  and2s1 U7599 ( .Q(WX3298), .DIN1(RESET), .DIN2(WX3235) );
  and2s1 U7600 ( .Q(WX3296), .DIN1(RESET), .DIN2(WX3233) );
  and2s1 U7601 ( .Q(WX3294), .DIN1(RESET), .DIN2(WX3231) );
  nnd4s1 U7602 ( .Q(WX3292), .DIN1(n5144), .DIN2(n5145), .DIN3(n5146), .DIN4(
        n5147) );
  nnd2s1 U7603 ( .Q(n5147), .DIN1(n3478), .DIN2(n4875) );
  xor2s1 U7604 ( .Q(n4875), .DIN1(n5148), .DIN2(n5149) );
  xor2s1 U7605 ( .Q(n5149), .DIN1(WX4650), .DIN2(n3173) );
  xor2s1 U7606 ( .Q(n5148), .DIN1(n3269), .DIN2(WX4714) );
  nnd2s1 U7607 ( .Q(n5146), .DIN1(n3440), .DIN2(n5150) );
  nnd2s1 U7608 ( .Q(n5145), .DIN1(WX3133), .DIN2(n3502) );
  nnd2s1 U7609 ( .Q(n5144), .DIN1(CRC_OUT_7_0), .DIN2(n3534) );
  nnd4s1 U7610 ( .Q(WX3290), .DIN1(n5151), .DIN2(n5152), .DIN3(n5153), .DIN4(
        n5154) );
  nnd2s1 U7611 ( .Q(n5154), .DIN1(n3478), .DIN2(n4882) );
  xor2s1 U7612 ( .Q(n4882), .DIN1(n5155), .DIN2(n5156) );
  xor2s1 U7613 ( .Q(n5156), .DIN1(WX4648), .DIN2(n3174) );
  xor2s1 U7614 ( .Q(n5155), .DIN1(n3270), .DIN2(WX4712) );
  nnd2s1 U7615 ( .Q(n5153), .DIN1(n3440), .DIN2(n5157) );
  nnd2s1 U7616 ( .Q(n5152), .DIN1(WX3131), .DIN2(n3502) );
  nnd2s1 U7617 ( .Q(n5151), .DIN1(CRC_OUT_7_1), .DIN2(n3534) );
  nnd4s1 U7618 ( .Q(WX3288), .DIN1(n5158), .DIN2(n5159), .DIN3(n5160), .DIN4(
        n5161) );
  nnd2s1 U7619 ( .Q(n5161), .DIN1(n3478), .DIN2(n4889) );
  xor2s1 U7620 ( .Q(n4889), .DIN1(n5162), .DIN2(n5163) );
  xor2s1 U7621 ( .Q(n5163), .DIN1(WX4646), .DIN2(n3175) );
  xor2s1 U7622 ( .Q(n5162), .DIN1(n3271), .DIN2(WX4710) );
  nnd2s1 U7623 ( .Q(n5160), .DIN1(n3440), .DIN2(n5164) );
  nnd2s1 U7624 ( .Q(n5159), .DIN1(WX3129), .DIN2(n3502) );
  nnd2s1 U7625 ( .Q(n5158), .DIN1(CRC_OUT_7_2), .DIN2(n3534) );
  nnd4s1 U7626 ( .Q(WX3286), .DIN1(n5165), .DIN2(n5166), .DIN3(n5167), .DIN4(
        n5168) );
  nnd2s1 U7627 ( .Q(n5168), .DIN1(n3479), .DIN2(n4896) );
  xor2s1 U7628 ( .Q(n4896), .DIN1(n5169), .DIN2(n5170) );
  xor2s1 U7629 ( .Q(n5170), .DIN1(WX4644), .DIN2(n3176) );
  xor2s1 U7630 ( .Q(n5169), .DIN1(n3272), .DIN2(WX4708) );
  nnd2s1 U7631 ( .Q(n5167), .DIN1(n3440), .DIN2(n5171) );
  nnd2s1 U7632 ( .Q(n5166), .DIN1(WX3127), .DIN2(n3502) );
  nnd2s1 U7633 ( .Q(n5165), .DIN1(CRC_OUT_7_3), .DIN2(n3534) );
  nnd4s1 U7634 ( .Q(WX3284), .DIN1(n5172), .DIN2(n5173), .DIN3(n5174), .DIN4(
        n5175) );
  nnd2s1 U7635 ( .Q(n5175), .DIN1(n3479), .DIN2(n4903) );
  xor2s1 U7636 ( .Q(n4903), .DIN1(n5176), .DIN2(n5177) );
  xor2s1 U7637 ( .Q(n5177), .DIN1(WX4642), .DIN2(n3177) );
  xor2s1 U7638 ( .Q(n5176), .DIN1(n3273), .DIN2(WX4706) );
  nnd2s1 U7639 ( .Q(n5174), .DIN1(n3440), .DIN2(n5178) );
  nnd2s1 U7640 ( .Q(n5173), .DIN1(WX3125), .DIN2(n3502) );
  nnd2s1 U7641 ( .Q(n5172), .DIN1(CRC_OUT_7_4), .DIN2(n3534) );
  nnd4s1 U7642 ( .Q(WX3282), .DIN1(n5179), .DIN2(n5180), .DIN3(n5181), .DIN4(
        n5182) );
  nnd2s1 U7643 ( .Q(n5182), .DIN1(n3479), .DIN2(n4910) );
  xor2s1 U7644 ( .Q(n4910), .DIN1(n5183), .DIN2(n5184) );
  xor2s1 U7645 ( .Q(n5184), .DIN1(WX4640), .DIN2(n3178) );
  xor2s1 U7646 ( .Q(n5183), .DIN1(n3274), .DIN2(WX4704) );
  nnd2s1 U7647 ( .Q(n5181), .DIN1(n3439), .DIN2(n5185) );
  nnd2s1 U7648 ( .Q(n5180), .DIN1(WX3123), .DIN2(n3502) );
  nnd2s1 U7649 ( .Q(n5179), .DIN1(CRC_OUT_7_5), .DIN2(n3534) );
  nnd4s1 U7650 ( .Q(WX3280), .DIN1(n5186), .DIN2(n5187), .DIN3(n5188), .DIN4(
        n5189) );
  nnd2s1 U7651 ( .Q(n5189), .DIN1(n3479), .DIN2(n4917) );
  xor2s1 U7652 ( .Q(n4917), .DIN1(n5190), .DIN2(n5191) );
  xor2s1 U7653 ( .Q(n5191), .DIN1(WX4638), .DIN2(n3179) );
  xor2s1 U7654 ( .Q(n5190), .DIN1(n3275), .DIN2(WX4702) );
  nnd2s1 U7655 ( .Q(n5188), .DIN1(n3439), .DIN2(n5192) );
  nnd2s1 U7656 ( .Q(n5187), .DIN1(WX3121), .DIN2(n3502) );
  nnd2s1 U7657 ( .Q(n5186), .DIN1(CRC_OUT_7_6), .DIN2(n3534) );
  nnd4s1 U7658 ( .Q(WX3278), .DIN1(n5193), .DIN2(n5194), .DIN3(n5195), .DIN4(
        n5196) );
  nnd2s1 U7659 ( .Q(n5196), .DIN1(n3479), .DIN2(n4924) );
  xor2s1 U7660 ( .Q(n4924), .DIN1(n5197), .DIN2(n5198) );
  xor2s1 U7661 ( .Q(n5198), .DIN1(WX4636), .DIN2(n3180) );
  xor2s1 U7662 ( .Q(n5197), .DIN1(n3276), .DIN2(WX4700) );
  nnd2s1 U7663 ( .Q(n5195), .DIN1(n3439), .DIN2(n5199) );
  nnd2s1 U7664 ( .Q(n5194), .DIN1(WX3119), .DIN2(n3502) );
  nnd2s1 U7665 ( .Q(n5193), .DIN1(CRC_OUT_7_7), .DIN2(n3534) );
  nnd4s1 U7666 ( .Q(WX3276), .DIN1(n5200), .DIN2(n5201), .DIN3(n5202), .DIN4(
        n5203) );
  nnd2s1 U7667 ( .Q(n5203), .DIN1(n3479), .DIN2(n4931) );
  xor2s1 U7668 ( .Q(n4931), .DIN1(n5204), .DIN2(n5205) );
  xor2s1 U7669 ( .Q(n5205), .DIN1(WX4634), .DIN2(n3181) );
  xor2s1 U7670 ( .Q(n5204), .DIN1(n3277), .DIN2(WX4698) );
  nnd2s1 U7671 ( .Q(n5202), .DIN1(n3439), .DIN2(n5206) );
  nnd2s1 U7672 ( .Q(n5201), .DIN1(WX3117), .DIN2(n3502) );
  nnd2s1 U7673 ( .Q(n5200), .DIN1(CRC_OUT_7_8), .DIN2(n3534) );
  nnd4s1 U7674 ( .Q(WX3274), .DIN1(n5207), .DIN2(n5208), .DIN3(n5209), .DIN4(
        n5210) );
  nnd2s1 U7675 ( .Q(n5210), .DIN1(n3479), .DIN2(n4938) );
  xor2s1 U7676 ( .Q(n4938), .DIN1(n5211), .DIN2(n5212) );
  xor2s1 U7677 ( .Q(n5212), .DIN1(WX4632), .DIN2(n3182) );
  xor2s1 U7678 ( .Q(n5211), .DIN1(n3278), .DIN2(WX4696) );
  nnd2s1 U7679 ( .Q(n5209), .DIN1(n3439), .DIN2(n5213) );
  nnd2s1 U7680 ( .Q(n5208), .DIN1(WX3115), .DIN2(n3502) );
  nnd2s1 U7681 ( .Q(n5207), .DIN1(CRC_OUT_7_9), .DIN2(n3534) );
  nnd4s1 U7682 ( .Q(WX3272), .DIN1(n5214), .DIN2(n5215), .DIN3(n5216), .DIN4(
        n5217) );
  nnd2s1 U7683 ( .Q(n5217), .DIN1(n3479), .DIN2(n4945) );
  xor2s1 U7684 ( .Q(n4945), .DIN1(n5218), .DIN2(n5219) );
  xor2s1 U7685 ( .Q(n5219), .DIN1(WX4630), .DIN2(n3183) );
  xor2s1 U7686 ( .Q(n5218), .DIN1(n3279), .DIN2(WX4694) );
  nnd2s1 U7687 ( .Q(n5216), .DIN1(n3439), .DIN2(n5220) );
  nnd2s1 U7688 ( .Q(n5215), .DIN1(WX3113), .DIN2(n3502) );
  nnd2s1 U7689 ( .Q(n5214), .DIN1(CRC_OUT_7_10), .DIN2(n3534) );
  nnd4s1 U7690 ( .Q(WX3270), .DIN1(n5221), .DIN2(n5222), .DIN3(n5223), .DIN4(
        n5224) );
  nnd2s1 U7691 ( .Q(n5224), .DIN1(n3479), .DIN2(n4952) );
  xor2s1 U7692 ( .Q(n4952), .DIN1(n5225), .DIN2(n5226) );
  xor2s1 U7693 ( .Q(n5226), .DIN1(WX4628), .DIN2(n3184) );
  xor2s1 U7694 ( .Q(n5225), .DIN1(n3280), .DIN2(WX4692) );
  nnd2s1 U7695 ( .Q(n5223), .DIN1(n3439), .DIN2(n5227) );
  nnd2s1 U7696 ( .Q(n5222), .DIN1(WX3111), .DIN2(n3502) );
  nnd2s1 U7697 ( .Q(n5221), .DIN1(CRC_OUT_7_11), .DIN2(n3534) );
  nnd4s1 U7698 ( .Q(WX3268), .DIN1(n5228), .DIN2(n5229), .DIN3(n5230), .DIN4(
        n5231) );
  nnd2s1 U7699 ( .Q(n5231), .DIN1(n3479), .DIN2(n4959) );
  xor2s1 U7700 ( .Q(n4959), .DIN1(n5232), .DIN2(n5233) );
  xor2s1 U7701 ( .Q(n5233), .DIN1(WX4626), .DIN2(n3185) );
  xor2s1 U7702 ( .Q(n5232), .DIN1(n3281), .DIN2(WX4690) );
  nnd2s1 U7703 ( .Q(n5230), .DIN1(n3439), .DIN2(n5234) );
  nnd2s1 U7704 ( .Q(n5229), .DIN1(WX3109), .DIN2(n3501) );
  nnd2s1 U7705 ( .Q(n5228), .DIN1(CRC_OUT_7_12), .DIN2(n3533) );
  nnd4s1 U7706 ( .Q(WX3266), .DIN1(n5235), .DIN2(n5236), .DIN3(n5237), .DIN4(
        n5238) );
  nnd2s1 U7707 ( .Q(n5238), .DIN1(n3479), .DIN2(n4966) );
  xor2s1 U7708 ( .Q(n4966), .DIN1(n5239), .DIN2(n5240) );
  xor2s1 U7709 ( .Q(n5240), .DIN1(WX4624), .DIN2(n3186) );
  xor2s1 U7710 ( .Q(n5239), .DIN1(n3282), .DIN2(WX4688) );
  nnd2s1 U7711 ( .Q(n5237), .DIN1(n3439), .DIN2(n5241) );
  nnd2s1 U7712 ( .Q(n5236), .DIN1(WX3107), .DIN2(n3501) );
  nnd2s1 U7713 ( .Q(n5235), .DIN1(CRC_OUT_7_13), .DIN2(n3533) );
  nnd4s1 U7714 ( .Q(WX3264), .DIN1(n5242), .DIN2(n5243), .DIN3(n5244), .DIN4(
        n5245) );
  nnd2s1 U7715 ( .Q(n5245), .DIN1(n3479), .DIN2(n4973) );
  xor2s1 U7716 ( .Q(n4973), .DIN1(n5246), .DIN2(n5247) );
  xor2s1 U7717 ( .Q(n5247), .DIN1(WX4622), .DIN2(n3187) );
  xor2s1 U7718 ( .Q(n5246), .DIN1(n3283), .DIN2(WX4686) );
  nnd2s1 U7719 ( .Q(n5244), .DIN1(n3439), .DIN2(n5248) );
  nnd2s1 U7720 ( .Q(n5243), .DIN1(WX3105), .DIN2(n3501) );
  nnd2s1 U7721 ( .Q(n5242), .DIN1(CRC_OUT_7_14), .DIN2(n3533) );
  nnd4s1 U7722 ( .Q(WX3262), .DIN1(n5249), .DIN2(n5250), .DIN3(n5251), .DIN4(
        n5252) );
  nnd2s1 U7723 ( .Q(n5252), .DIN1(n3479), .DIN2(n4980) );
  xor2s1 U7724 ( .Q(n4980), .DIN1(n5253), .DIN2(n5254) );
  xor2s1 U7725 ( .Q(n5254), .DIN1(WX4620), .DIN2(n3188) );
  xor2s1 U7726 ( .Q(n5253), .DIN1(n3284), .DIN2(WX4684) );
  nnd2s1 U7727 ( .Q(n5251), .DIN1(n3439), .DIN2(n5255) );
  nnd2s1 U7728 ( .Q(n5250), .DIN1(WX3103), .DIN2(n3501) );
  nnd2s1 U7729 ( .Q(n5249), .DIN1(CRC_OUT_7_15), .DIN2(n3533) );
  nnd4s1 U7730 ( .Q(WX3260), .DIN1(n5256), .DIN2(n5257), .DIN3(n5258), .DIN4(
        n5259) );
  nnd2s1 U7731 ( .Q(n5259), .DIN1(n3480), .DIN2(n4988) );
  xor2s1 U7732 ( .Q(n4988), .DIN1(n5260), .DIN2(n5261) );
  xor2s1 U7733 ( .Q(n5261), .DIN1(n3568), .DIN2(WX4554) );
  xor2s1 U7734 ( .Q(n5260), .DIN1(n3013), .DIN2(n5262) );
  xor2s1 U7735 ( .Q(n5262), .DIN1(WX4746), .DIN2(WX4682) );
  nnd2s1 U7736 ( .Q(n5258), .DIN1(n3439), .DIN2(n5263) );
  nnd2s1 U7737 ( .Q(n5257), .DIN1(WX3101), .DIN2(n3501) );
  nnd2s1 U7738 ( .Q(n5256), .DIN1(CRC_OUT_7_16), .DIN2(n3533) );
  nnd4s1 U7739 ( .Q(WX3258), .DIN1(n5264), .DIN2(n5265), .DIN3(n5266), .DIN4(
        n5267) );
  nnd2s1 U7740 ( .Q(n5267), .DIN1(n3480), .DIN2(n4996) );
  xor2s1 U7741 ( .Q(n4996), .DIN1(n5268), .DIN2(n5269) );
  xor2s1 U7742 ( .Q(n5269), .DIN1(n3568), .DIN2(WX4552) );
  xor2s1 U7743 ( .Q(n5268), .DIN1(n3014), .DIN2(n5270) );
  xor2s1 U7744 ( .Q(n5270), .DIN1(WX4744), .DIN2(WX4680) );
  nnd2s1 U7745 ( .Q(n5266), .DIN1(n3439), .DIN2(n5271) );
  nnd2s1 U7746 ( .Q(n5265), .DIN1(WX3099), .DIN2(n3501) );
  nnd2s1 U7747 ( .Q(n5264), .DIN1(CRC_OUT_7_17), .DIN2(n3533) );
  nnd4s1 U7748 ( .Q(WX3256), .DIN1(n5272), .DIN2(n5273), .DIN3(n5274), .DIN4(
        n5275) );
  nnd2s1 U7749 ( .Q(n5275), .DIN1(n3480), .DIN2(n5004) );
  xor2s1 U7750 ( .Q(n5004), .DIN1(n5276), .DIN2(n5277) );
  xor2s1 U7751 ( .Q(n5277), .DIN1(n3568), .DIN2(WX4550) );
  xor2s1 U7752 ( .Q(n5276), .DIN1(n3015), .DIN2(n5278) );
  xor2s1 U7753 ( .Q(n5278), .DIN1(WX4742), .DIN2(WX4678) );
  nnd2s1 U7754 ( .Q(n5274), .DIN1(n3438), .DIN2(n5279) );
  nnd2s1 U7755 ( .Q(n5273), .DIN1(WX3097), .DIN2(n3501) );
  nnd2s1 U7756 ( .Q(n5272), .DIN1(CRC_OUT_7_18), .DIN2(n3533) );
  nnd4s1 U7757 ( .Q(WX3254), .DIN1(n5280), .DIN2(n5281), .DIN3(n5282), .DIN4(
        n5283) );
  nnd2s1 U7758 ( .Q(n5283), .DIN1(n3480), .DIN2(n5012) );
  xor2s1 U7759 ( .Q(n5012), .DIN1(n5284), .DIN2(n5285) );
  xor2s1 U7760 ( .Q(n5285), .DIN1(n3568), .DIN2(WX4548) );
  xor2s1 U7761 ( .Q(n5284), .DIN1(n3016), .DIN2(n5286) );
  xor2s1 U7762 ( .Q(n5286), .DIN1(WX4740), .DIN2(WX4676) );
  nnd2s1 U7763 ( .Q(n5282), .DIN1(n3438), .DIN2(n5287) );
  nnd2s1 U7764 ( .Q(n5281), .DIN1(WX3095), .DIN2(n3501) );
  nnd2s1 U7765 ( .Q(n5280), .DIN1(CRC_OUT_7_19), .DIN2(n3533) );
  nnd4s1 U7766 ( .Q(WX3252), .DIN1(n5288), .DIN2(n5289), .DIN3(n5290), .DIN4(
        n5291) );
  nnd2s1 U7767 ( .Q(n5291), .DIN1(n3480), .DIN2(n5020) );
  xor2s1 U7768 ( .Q(n5020), .DIN1(n5292), .DIN2(n5293) );
  xor2s1 U7769 ( .Q(n5293), .DIN1(n3568), .DIN2(WX4546) );
  xor2s1 U7770 ( .Q(n5292), .DIN1(n3017), .DIN2(n5294) );
  xor2s1 U7771 ( .Q(n5294), .DIN1(WX4738), .DIN2(WX4674) );
  nnd2s1 U7772 ( .Q(n5290), .DIN1(n3438), .DIN2(n5295) );
  nnd2s1 U7773 ( .Q(n5289), .DIN1(WX3093), .DIN2(n3501) );
  nnd2s1 U7774 ( .Q(n5288), .DIN1(CRC_OUT_7_20), .DIN2(n3533) );
  nnd4s1 U7775 ( .Q(WX3250), .DIN1(n5296), .DIN2(n5297), .DIN3(n5298), .DIN4(
        n5299) );
  nnd2s1 U7776 ( .Q(n5299), .DIN1(n3480), .DIN2(n5028) );
  xor2s1 U7777 ( .Q(n5028), .DIN1(n5300), .DIN2(n5301) );
  xor2s1 U7778 ( .Q(n5301), .DIN1(n3568), .DIN2(WX4544) );
  xor2s1 U7779 ( .Q(n5300), .DIN1(n3018), .DIN2(n5302) );
  xor2s1 U7780 ( .Q(n5302), .DIN1(WX4736), .DIN2(WX4672) );
  nnd2s1 U7781 ( .Q(n5298), .DIN1(n3438), .DIN2(n5303) );
  nnd2s1 U7782 ( .Q(n5297), .DIN1(WX3091), .DIN2(n3501) );
  nnd2s1 U7783 ( .Q(n5296), .DIN1(CRC_OUT_7_21), .DIN2(n3533) );
  nnd4s1 U7784 ( .Q(WX3248), .DIN1(n5304), .DIN2(n5305), .DIN3(n5306), .DIN4(
        n5307) );
  nnd2s1 U7785 ( .Q(n5307), .DIN1(n3480), .DIN2(n5036) );
  xor2s1 U7786 ( .Q(n5036), .DIN1(n5308), .DIN2(n5309) );
  xor2s1 U7787 ( .Q(n5309), .DIN1(n3569), .DIN2(WX4542) );
  xor2s1 U7788 ( .Q(n5308), .DIN1(n3019), .DIN2(n5310) );
  xor2s1 U7789 ( .Q(n5310), .DIN1(WX4734), .DIN2(WX4670) );
  nnd2s1 U7790 ( .Q(n5306), .DIN1(n3438), .DIN2(n5311) );
  nnd2s1 U7791 ( .Q(n5305), .DIN1(WX3089), .DIN2(n3501) );
  nnd2s1 U7792 ( .Q(n5304), .DIN1(CRC_OUT_7_22), .DIN2(n3533) );
  nnd4s1 U7793 ( .Q(WX3246), .DIN1(n5312), .DIN2(n5313), .DIN3(n5314), .DIN4(
        n5315) );
  nnd2s1 U7794 ( .Q(n5315), .DIN1(n3480), .DIN2(n5044) );
  xor2s1 U7795 ( .Q(n5044), .DIN1(n5316), .DIN2(n5317) );
  xor2s1 U7796 ( .Q(n5317), .DIN1(n3569), .DIN2(WX4540) );
  xor2s1 U7797 ( .Q(n5316), .DIN1(n3020), .DIN2(n5318) );
  xor2s1 U7798 ( .Q(n5318), .DIN1(WX4732), .DIN2(WX4668) );
  nnd2s1 U7799 ( .Q(n5314), .DIN1(n3438), .DIN2(n5319) );
  nnd2s1 U7800 ( .Q(n5313), .DIN1(WX3087), .DIN2(n3501) );
  nnd2s1 U7801 ( .Q(n5312), .DIN1(CRC_OUT_7_23), .DIN2(n3533) );
  nnd4s1 U7802 ( .Q(WX3244), .DIN1(n5320), .DIN2(n5321), .DIN3(n5322), .DIN4(
        n5323) );
  nnd2s1 U7803 ( .Q(n5323), .DIN1(n3480), .DIN2(n5052) );
  xor2s1 U7804 ( .Q(n5052), .DIN1(n5324), .DIN2(n5325) );
  xor2s1 U7805 ( .Q(n5325), .DIN1(n3569), .DIN2(WX4538) );
  xor2s1 U7806 ( .Q(n5324), .DIN1(n3021), .DIN2(n5326) );
  xor2s1 U7807 ( .Q(n5326), .DIN1(WX4730), .DIN2(WX4666) );
  nnd2s1 U7808 ( .Q(n5322), .DIN1(n3438), .DIN2(n5327) );
  nnd2s1 U7809 ( .Q(n5321), .DIN1(WX3085), .DIN2(n3500) );
  nnd2s1 U7810 ( .Q(n5320), .DIN1(CRC_OUT_7_24), .DIN2(n3532) );
  nnd4s1 U7811 ( .Q(WX3242), .DIN1(n5328), .DIN2(n5329), .DIN3(n5330), .DIN4(
        n5331) );
  nnd2s1 U7812 ( .Q(n5331), .DIN1(n3480), .DIN2(n5060) );
  xor2s1 U7813 ( .Q(n5060), .DIN1(n5332), .DIN2(n5333) );
  xor2s1 U7814 ( .Q(n5333), .DIN1(n3569), .DIN2(WX4536) );
  xor2s1 U7815 ( .Q(n5332), .DIN1(n3022), .DIN2(n5334) );
  xor2s1 U7816 ( .Q(n5334), .DIN1(WX4728), .DIN2(WX4664) );
  nnd2s1 U7817 ( .Q(n5330), .DIN1(n3438), .DIN2(n5335) );
  nnd2s1 U7818 ( .Q(n5329), .DIN1(WX3083), .DIN2(n3500) );
  nnd2s1 U7819 ( .Q(n5328), .DIN1(CRC_OUT_7_25), .DIN2(n3532) );
  nnd4s1 U7820 ( .Q(WX3240), .DIN1(n5336), .DIN2(n5337), .DIN3(n5338), .DIN4(
        n5339) );
  nnd2s1 U7821 ( .Q(n5339), .DIN1(n3480), .DIN2(n5068) );
  xor2s1 U7822 ( .Q(n5068), .DIN1(n5340), .DIN2(n5341) );
  xor2s1 U7823 ( .Q(n5341), .DIN1(n3569), .DIN2(WX4534) );
  xor2s1 U7824 ( .Q(n5340), .DIN1(n3023), .DIN2(n5342) );
  xor2s1 U7825 ( .Q(n5342), .DIN1(WX4726), .DIN2(WX4662) );
  nnd2s1 U7826 ( .Q(n5338), .DIN1(n3438), .DIN2(n5343) );
  nnd2s1 U7827 ( .Q(n5337), .DIN1(WX3081), .DIN2(n3500) );
  nnd2s1 U7828 ( .Q(n5336), .DIN1(CRC_OUT_7_26), .DIN2(n3532) );
  nnd4s1 U7829 ( .Q(WX3238), .DIN1(n5344), .DIN2(n5345), .DIN3(n5346), .DIN4(
        n5347) );
  nnd2s1 U7830 ( .Q(n5347), .DIN1(n3480), .DIN2(n5076) );
  xor2s1 U7831 ( .Q(n5076), .DIN1(n5348), .DIN2(n5349) );
  xor2s1 U7832 ( .Q(n5349), .DIN1(n3569), .DIN2(WX4532) );
  xor2s1 U7833 ( .Q(n5348), .DIN1(n3024), .DIN2(n5350) );
  xor2s1 U7834 ( .Q(n5350), .DIN1(WX4724), .DIN2(WX4660) );
  nnd2s1 U7835 ( .Q(n5346), .DIN1(n3438), .DIN2(n5351) );
  nnd2s1 U7836 ( .Q(n5345), .DIN1(WX3079), .DIN2(n3500) );
  nnd2s1 U7837 ( .Q(n5344), .DIN1(CRC_OUT_7_27), .DIN2(n3532) );
  nnd4s1 U7838 ( .Q(WX3236), .DIN1(n5352), .DIN2(n5353), .DIN3(n5354), .DIN4(
        n5355) );
  nnd2s1 U7839 ( .Q(n5355), .DIN1(n3480), .DIN2(n5084) );
  xor2s1 U7840 ( .Q(n5084), .DIN1(n5356), .DIN2(n5357) );
  xor2s1 U7841 ( .Q(n5357), .DIN1(n3570), .DIN2(WX4530) );
  xor2s1 U7842 ( .Q(n5356), .DIN1(n3025), .DIN2(n5358) );
  xor2s1 U7843 ( .Q(n5358), .DIN1(WX4722), .DIN2(WX4658) );
  nnd2s1 U7844 ( .Q(n5354), .DIN1(n3438), .DIN2(n5359) );
  nnd2s1 U7845 ( .Q(n5353), .DIN1(WX3077), .DIN2(n3500) );
  nnd2s1 U7846 ( .Q(n5352), .DIN1(CRC_OUT_7_28), .DIN2(n3532) );
  nnd4s1 U7847 ( .Q(WX3234), .DIN1(n5360), .DIN2(n5361), .DIN3(n5362), .DIN4(
        n5363) );
  nnd2s1 U7848 ( .Q(n5363), .DIN1(n3481), .DIN2(n5092) );
  xor2s1 U7849 ( .Q(n5092), .DIN1(n5364), .DIN2(n5365) );
  xor2s1 U7850 ( .Q(n5365), .DIN1(n3570), .DIN2(WX4528) );
  xor2s1 U7851 ( .Q(n5364), .DIN1(n3026), .DIN2(n5366) );
  xor2s1 U7852 ( .Q(n5366), .DIN1(WX4720), .DIN2(WX4656) );
  nnd2s1 U7853 ( .Q(n5362), .DIN1(n3438), .DIN2(n5367) );
  nnd2s1 U7854 ( .Q(n5361), .DIN1(WX3075), .DIN2(n3500) );
  nnd2s1 U7855 ( .Q(n5360), .DIN1(CRC_OUT_7_29), .DIN2(n3532) );
  nnd4s1 U7856 ( .Q(WX3232), .DIN1(n5368), .DIN2(n5369), .DIN3(n5370), .DIN4(
        n5371) );
  nnd2s1 U7857 ( .Q(n5371), .DIN1(n3481), .DIN2(n5100) );
  xor2s1 U7858 ( .Q(n5100), .DIN1(n5372), .DIN2(n5373) );
  xor2s1 U7859 ( .Q(n5373), .DIN1(n3570), .DIN2(WX4526) );
  xor2s1 U7860 ( .Q(n5372), .DIN1(n3027), .DIN2(n5374) );
  xor2s1 U7861 ( .Q(n5374), .DIN1(WX4718), .DIN2(WX4654) );
  nnd2s1 U7862 ( .Q(n5370), .DIN1(n3438), .DIN2(n5375) );
  nnd2s1 U7863 ( .Q(n5369), .DIN1(WX3073), .DIN2(n3500) );
  nnd2s1 U7864 ( .Q(n5368), .DIN1(CRC_OUT_7_30), .DIN2(n3532) );
  nnd4s1 U7865 ( .Q(WX3230), .DIN1(n5376), .DIN2(n5377), .DIN3(n5378), .DIN4(
        n5379) );
  nnd2s1 U7866 ( .Q(n5379), .DIN1(n3481), .DIN2(n5108) );
  xor2s1 U7867 ( .Q(n5108), .DIN1(n5380), .DIN2(n5381) );
  xor2s1 U7868 ( .Q(n5381), .DIN1(n3570), .DIN2(WX4524) );
  xor2s1 U7869 ( .Q(n5380), .DIN1(n3028), .DIN2(n5382) );
  xor2s1 U7870 ( .Q(n5382), .DIN1(WX4716), .DIN2(WX4652) );
  nnd2s1 U7871 ( .Q(n5378), .DIN1(n3437), .DIN2(n5383) );
  nnd2s1 U7872 ( .Q(n5377), .DIN1(WX3071), .DIN2(n3500) );
  nnd2s1 U7873 ( .Q(n5376), .DIN1(CRC_OUT_7_31), .DIN2(n3532) );
  nor2s1 U7874 ( .Q(WX3132), .DIN1(WX3071), .DIN2(n3363) );
  and2s1 U7875 ( .Q(WX3130), .DIN1(RESET), .DIN2(WX3133) );
  and2s1 U7876 ( .Q(WX3128), .DIN1(RESET), .DIN2(WX3131) );
  and2s1 U7877 ( .Q(WX3126), .DIN1(RESET), .DIN2(WX3129) );
  and2s1 U7878 ( .Q(WX3124), .DIN1(RESET), .DIN2(WX3127) );
  and2s1 U7879 ( .Q(WX3122), .DIN1(RESET), .DIN2(WX3125) );
  and2s1 U7880 ( .Q(WX3120), .DIN1(RESET), .DIN2(WX3123) );
  and2s1 U7881 ( .Q(WX3118), .DIN1(RESET), .DIN2(WX3121) );
  and2s1 U7882 ( .Q(WX3116), .DIN1(RESET), .DIN2(WX3119) );
  and2s1 U7883 ( .Q(WX3114), .DIN1(RESET), .DIN2(WX3117) );
  and2s1 U7884 ( .Q(WX3112), .DIN1(RESET), .DIN2(WX3115) );
  and2s1 U7885 ( .Q(WX3110), .DIN1(RESET), .DIN2(WX3113) );
  and2s1 U7886 ( .Q(WX3108), .DIN1(RESET), .DIN2(WX3111) );
  and2s1 U7887 ( .Q(WX3106), .DIN1(RESET), .DIN2(WX3109) );
  and2s1 U7888 ( .Q(WX3104), .DIN1(RESET), .DIN2(WX3107) );
  and2s1 U7889 ( .Q(WX3102), .DIN1(RESET), .DIN2(WX3105) );
  and2s1 U7890 ( .Q(WX3100), .DIN1(RESET), .DIN2(WX3103) );
  and2s1 U7891 ( .Q(WX3098), .DIN1(RESET), .DIN2(WX3101) );
  and2s1 U7892 ( .Q(WX3096), .DIN1(RESET), .DIN2(WX3099) );
  and2s1 U7893 ( .Q(WX3094), .DIN1(RESET), .DIN2(WX3097) );
  and2s1 U7894 ( .Q(WX3092), .DIN1(RESET), .DIN2(WX3095) );
  and2s1 U7895 ( .Q(WX3090), .DIN1(RESET), .DIN2(WX3093) );
  and2s1 U7896 ( .Q(WX3088), .DIN1(RESET), .DIN2(WX3091) );
  and2s1 U7897 ( .Q(WX3086), .DIN1(RESET), .DIN2(WX3089) );
  and2s1 U7898 ( .Q(WX3084), .DIN1(RESET), .DIN2(WX3087) );
  and2s1 U7899 ( .Q(WX3082), .DIN1(RESET), .DIN2(WX3085) );
  and2s1 U7900 ( .Q(WX3080), .DIN1(RESET), .DIN2(WX3083) );
  and2s1 U7901 ( .Q(WX3078), .DIN1(RESET), .DIN2(WX3081) );
  and2s1 U7902 ( .Q(WX3076), .DIN1(RESET), .DIN2(WX3079) );
  and2s1 U7903 ( .Q(WX3074), .DIN1(RESET), .DIN2(WX3077) );
  and2s1 U7904 ( .Q(WX3072), .DIN1(RESET), .DIN2(WX3075) );
  and2s1 U7905 ( .Q(WX3070), .DIN1(RESET), .DIN2(WX3073) );
  nor2s1 U7906 ( .Q(WX2619), .DIN1(n3412), .DIN2(n5384) );
  xor2s1 U7907 ( .Q(n5384), .DIN1(WX2130), .DIN2(CRC_OUT_8_30) );
  nor2s1 U7908 ( .Q(WX2617), .DIN1(n3413), .DIN2(n5385) );
  xor2s1 U7909 ( .Q(n5385), .DIN1(WX2132), .DIN2(CRC_OUT_8_29) );
  nor2s1 U7910 ( .Q(WX2615), .DIN1(n3413), .DIN2(n5386) );
  xor2s1 U7911 ( .Q(n5386), .DIN1(WX2134), .DIN2(CRC_OUT_8_28) );
  nor2s1 U7912 ( .Q(WX2613), .DIN1(n3413), .DIN2(n5387) );
  xor2s1 U7913 ( .Q(n5387), .DIN1(WX2136), .DIN2(CRC_OUT_8_27) );
  nor2s1 U7914 ( .Q(WX2611), .DIN1(n3413), .DIN2(n5388) );
  xor2s1 U7915 ( .Q(n5388), .DIN1(WX2138), .DIN2(CRC_OUT_8_26) );
  nor2s1 U7916 ( .Q(WX2609), .DIN1(n3413), .DIN2(n5389) );
  xor2s1 U7917 ( .Q(n5389), .DIN1(WX2140), .DIN2(CRC_OUT_8_25) );
  nor2s1 U7918 ( .Q(WX2607), .DIN1(n3413), .DIN2(n5390) );
  xor2s1 U7919 ( .Q(n5390), .DIN1(WX2142), .DIN2(CRC_OUT_8_24) );
  nor2s1 U7920 ( .Q(WX2605), .DIN1(n3413), .DIN2(n5391) );
  xor2s1 U7921 ( .Q(n5391), .DIN1(WX2144), .DIN2(CRC_OUT_8_23) );
  nor2s1 U7922 ( .Q(WX2603), .DIN1(n3413), .DIN2(n5392) );
  xor2s1 U7923 ( .Q(n5392), .DIN1(WX2146), .DIN2(CRC_OUT_8_22) );
  nor2s1 U7924 ( .Q(WX2601), .DIN1(n3413), .DIN2(n5393) );
  xor2s1 U7925 ( .Q(n5393), .DIN1(WX2148), .DIN2(CRC_OUT_8_21) );
  nor2s1 U7926 ( .Q(WX2599), .DIN1(n3413), .DIN2(n5394) );
  xor2s1 U7927 ( .Q(n5394), .DIN1(WX2150), .DIN2(CRC_OUT_8_20) );
  nor2s1 U7928 ( .Q(WX2597), .DIN1(n3414), .DIN2(n5395) );
  xor2s1 U7929 ( .Q(n5395), .DIN1(WX2152), .DIN2(CRC_OUT_8_19) );
  nor2s1 U7930 ( .Q(WX2595), .DIN1(n3414), .DIN2(n5396) );
  xor2s1 U7931 ( .Q(n5396), .DIN1(WX2154), .DIN2(CRC_OUT_8_18) );
  nor2s1 U7932 ( .Q(WX2593), .DIN1(n3414), .DIN2(n5397) );
  xor2s1 U7933 ( .Q(n5397), .DIN1(WX2156), .DIN2(CRC_OUT_8_17) );
  nor2s1 U7934 ( .Q(WX2591), .DIN1(n3414), .DIN2(n5398) );
  xor2s1 U7935 ( .Q(n5398), .DIN1(WX2158), .DIN2(CRC_OUT_8_16) );
  nor2s1 U7936 ( .Q(WX2589), .DIN1(n3414), .DIN2(n5399) );
  xor2s1 U7937 ( .Q(n5399), .DIN1(CRC_OUT_8_15), .DIN2(n5400) );
  xor2s1 U7938 ( .Q(n5400), .DIN1(WX2160), .DIN2(CRC_OUT_8_31) );
  nor2s1 U7939 ( .Q(WX2587), .DIN1(n3414), .DIN2(n5401) );
  xor2s1 U7940 ( .Q(n5401), .DIN1(WX2162), .DIN2(CRC_OUT_8_14) );
  nor2s1 U7941 ( .Q(WX2585), .DIN1(n3414), .DIN2(n5402) );
  xor2s1 U7942 ( .Q(n5402), .DIN1(WX2164), .DIN2(CRC_OUT_8_13) );
  nor2s1 U7943 ( .Q(WX2583), .DIN1(n3414), .DIN2(n5403) );
  xor2s1 U7944 ( .Q(n5403), .DIN1(WX2166), .DIN2(CRC_OUT_8_12) );
  nor2s1 U7945 ( .Q(WX2581), .DIN1(n3414), .DIN2(n5404) );
  xor2s1 U7946 ( .Q(n5404), .DIN1(WX2168), .DIN2(CRC_OUT_8_11) );
  nor2s1 U7947 ( .Q(WX2579), .DIN1(n3414), .DIN2(n5405) );
  xor2s1 U7948 ( .Q(n5405), .DIN1(CRC_OUT_8_10), .DIN2(n5406) );
  xor2s1 U7949 ( .Q(n5406), .DIN1(WX2170), .DIN2(CRC_OUT_8_31) );
  nor2s1 U7950 ( .Q(WX2577), .DIN1(n3415), .DIN2(n5407) );
  xor2s1 U7951 ( .Q(n5407), .DIN1(WX2172), .DIN2(CRC_OUT_8_9) );
  nor2s1 U7952 ( .Q(WX2575), .DIN1(n3415), .DIN2(n5408) );
  xor2s1 U7953 ( .Q(n5408), .DIN1(WX2174), .DIN2(CRC_OUT_8_8) );
  nor2s1 U7954 ( .Q(WX2573), .DIN1(n3415), .DIN2(n5409) );
  xor2s1 U7955 ( .Q(n5409), .DIN1(WX2176), .DIN2(CRC_OUT_8_7) );
  nor2s1 U7956 ( .Q(WX2571), .DIN1(n3415), .DIN2(n5410) );
  xor2s1 U7957 ( .Q(n5410), .DIN1(WX2178), .DIN2(CRC_OUT_8_6) );
  nor2s1 U7958 ( .Q(WX2569), .DIN1(n3415), .DIN2(n5411) );
  xor2s1 U7959 ( .Q(n5411), .DIN1(WX2180), .DIN2(CRC_OUT_8_5) );
  nor2s1 U7960 ( .Q(WX2567), .DIN1(n3415), .DIN2(n5412) );
  xor2s1 U7961 ( .Q(n5412), .DIN1(WX2182), .DIN2(CRC_OUT_8_4) );
  nor2s1 U7962 ( .Q(WX2565), .DIN1(n3415), .DIN2(n5413) );
  xor2s1 U7963 ( .Q(n5413), .DIN1(CRC_OUT_8_3), .DIN2(n5414) );
  xor2s1 U7964 ( .Q(n5414), .DIN1(WX2184), .DIN2(CRC_OUT_8_31) );
  nor2s1 U7965 ( .Q(WX2563), .DIN1(n3415), .DIN2(n5415) );
  xor2s1 U7966 ( .Q(n5415), .DIN1(WX2186), .DIN2(CRC_OUT_8_2) );
  nor2s1 U7967 ( .Q(WX2561), .DIN1(n3415), .DIN2(n5416) );
  xor2s1 U7968 ( .Q(n5416), .DIN1(WX2188), .DIN2(CRC_OUT_8_1) );
  nor2s1 U7969 ( .Q(WX2559), .DIN1(n3415), .DIN2(n5417) );
  xor2s1 U7970 ( .Q(n5417), .DIN1(WX2190), .DIN2(CRC_OUT_8_0) );
  nor2s1 U7971 ( .Q(WX2557), .DIN1(n3416), .DIN2(n5418) );
  xor2s1 U7972 ( .Q(n5418), .DIN1(WX2192), .DIN2(CRC_OUT_8_31) );
  and2s1 U7973 ( .Q(WX2191), .DIN1(RESET), .DIN2(WX2128) );
  and2s1 U7974 ( .Q(WX2189), .DIN1(RESET), .DIN2(WX2126) );
  and2s1 U7975 ( .Q(WX2187), .DIN1(RESET), .DIN2(WX2124) );
  and2s1 U7976 ( .Q(WX2185), .DIN1(RESET), .DIN2(WX2122) );
  and2s1 U7977 ( .Q(WX2183), .DIN1(RESET), .DIN2(WX2120) );
  and2s1 U7978 ( .Q(WX2181), .DIN1(RESET), .DIN2(WX2118) );
  and2s1 U7979 ( .Q(WX2179), .DIN1(RESET), .DIN2(WX2116) );
  and2s1 U7980 ( .Q(WX2177), .DIN1(RESET), .DIN2(WX2114) );
  and2s1 U7981 ( .Q(WX2175), .DIN1(RESET), .DIN2(WX2112) );
  and2s1 U7982 ( .Q(WX2173), .DIN1(RESET), .DIN2(WX2110) );
  and2s1 U7983 ( .Q(WX2171), .DIN1(RESET), .DIN2(WX2108) );
  and2s1 U7984 ( .Q(WX2169), .DIN1(RESET), .DIN2(WX2106) );
  and2s1 U7985 ( .Q(WX2167), .DIN1(RESET), .DIN2(WX2104) );
  and2s1 U7986 ( .Q(WX2165), .DIN1(RESET), .DIN2(WX2102) );
  and2s1 U7987 ( .Q(WX2163), .DIN1(RESET), .DIN2(WX2100) );
  and2s1 U7988 ( .Q(WX2161), .DIN1(RESET), .DIN2(WX2098) );
  and2s1 U7989 ( .Q(WX2159), .DIN1(RESET), .DIN2(WX2096) );
  and2s1 U7990 ( .Q(WX2157), .DIN1(RESET), .DIN2(WX2094) );
  and2s1 U7991 ( .Q(WX2155), .DIN1(RESET), .DIN2(WX2092) );
  and2s1 U7992 ( .Q(WX2153), .DIN1(RESET), .DIN2(WX2090) );
  and2s1 U7993 ( .Q(WX2151), .DIN1(RESET), .DIN2(WX2088) );
  and2s1 U7994 ( .Q(WX2149), .DIN1(RESET), .DIN2(WX2086) );
  and2s1 U7995 ( .Q(WX2147), .DIN1(RESET), .DIN2(WX2084) );
  and2s1 U7996 ( .Q(WX2145), .DIN1(RESET), .DIN2(WX2082) );
  and2s1 U7997 ( .Q(WX2143), .DIN1(RESET), .DIN2(WX2080) );
  and2s1 U7998 ( .Q(WX2141), .DIN1(RESET), .DIN2(WX2078) );
  and2s1 U7999 ( .Q(WX2139), .DIN1(RESET), .DIN2(WX2076) );
  and2s1 U8000 ( .Q(WX2137), .DIN1(RESET), .DIN2(WX2074) );
  and2s1 U8001 ( .Q(WX2135), .DIN1(RESET), .DIN2(WX2072) );
  and2s1 U8002 ( .Q(WX2133), .DIN1(RESET), .DIN2(WX2070) );
  and2s1 U8003 ( .Q(WX2131), .DIN1(RESET), .DIN2(WX2068) );
  and2s1 U8004 ( .Q(WX2129), .DIN1(RESET), .DIN2(WX2066) );
  nor2s1 U8005 ( .Q(WX2127), .DIN1(n3416), .DIN2(n3029) );
  nor2s1 U8006 ( .Q(WX2125), .DIN1(n3416), .DIN2(n3030) );
  nor2s1 U8007 ( .Q(WX2123), .DIN1(n3416), .DIN2(n3031) );
  nor2s1 U8008 ( .Q(WX2121), .DIN1(n3416), .DIN2(n3032) );
  nor2s1 U8009 ( .Q(WX2119), .DIN1(n3416), .DIN2(n3033) );
  nor2s1 U8010 ( .Q(WX2117), .DIN1(n3416), .DIN2(n3034) );
  nor2s1 U8011 ( .Q(WX2115), .DIN1(n3416), .DIN2(n3035) );
  nor2s1 U8012 ( .Q(WX2113), .DIN1(n3416), .DIN2(n3036) );
  nor2s1 U8013 ( .Q(WX2111), .DIN1(n3416), .DIN2(n3037) );
  nor2s1 U8014 ( .Q(WX2109), .DIN1(n3417), .DIN2(n3038) );
  nor2s1 U8015 ( .Q(WX2107), .DIN1(n3417), .DIN2(n3039) );
  nor2s1 U8016 ( .Q(WX2105), .DIN1(n3417), .DIN2(n3040) );
  nor2s1 U8017 ( .Q(WX2103), .DIN1(n3417), .DIN2(n3041) );
  nor2s1 U8018 ( .Q(WX2101), .DIN1(n3417), .DIN2(n3042) );
  nor2s1 U8019 ( .Q(WX2099), .DIN1(n3417), .DIN2(n3043) );
  nor2s1 U8020 ( .Q(WX2097), .DIN1(n3417), .DIN2(n3044) );
  nor2s1 U8021 ( .Q(WX2095), .DIN1(n3417), .DIN2(n3046) );
  nor2s1 U8022 ( .Q(WX2093), .DIN1(n3417), .DIN2(n3048) );
  nor2s1 U8023 ( .Q(WX2091), .DIN1(n3417), .DIN2(n3050) );
  nor2s1 U8024 ( .Q(WX2089), .DIN1(n3418), .DIN2(n3052) );
  nor2s1 U8025 ( .Q(WX2087), .DIN1(n3418), .DIN2(n3054) );
  nor2s1 U8026 ( .Q(WX2085), .DIN1(n3418), .DIN2(n3056) );
  nor2s1 U8027 ( .Q(WX2083), .DIN1(n3397), .DIN2(n3058) );
  nor2s1 U8028 ( .Q(WX2081), .DIN1(n3390), .DIN2(n3060) );
  nor2s1 U8029 ( .Q(WX2079), .DIN1(n3391), .DIN2(n3062) );
  nor2s1 U8030 ( .Q(WX2077), .DIN1(n3391), .DIN2(n3064) );
  nor2s1 U8031 ( .Q(WX2075), .DIN1(n3391), .DIN2(n3066) );
  nor2s1 U8032 ( .Q(WX2073), .DIN1(n3391), .DIN2(n3068) );
  nor2s1 U8033 ( .Q(WX2071), .DIN1(n3391), .DIN2(n3070) );
  nor2s1 U8034 ( .Q(WX2069), .DIN1(n3391), .DIN2(n3072) );
  nor2s1 U8035 ( .Q(WX2067), .DIN1(n3391), .DIN2(n3074) );
  nor2s1 U8036 ( .Q(WX2065), .DIN1(n3391), .DIN2(n3076) );
  and2s1 U8037 ( .Q(WX2063), .DIN1(RESET), .DIN2(WX2000) );
  and2s1 U8038 ( .Q(WX2061), .DIN1(RESET), .DIN2(WX1998) );
  and2s1 U8039 ( .Q(WX2059), .DIN1(RESET), .DIN2(WX1996) );
  and2s1 U8040 ( .Q(WX2057), .DIN1(RESET), .DIN2(WX1994) );
  and2s1 U8041 ( .Q(WX2055), .DIN1(RESET), .DIN2(WX1992) );
  and2s1 U8042 ( .Q(WX2053), .DIN1(RESET), .DIN2(WX1990) );
  and2s1 U8043 ( .Q(WX2051), .DIN1(RESET), .DIN2(WX1988) );
  and2s1 U8044 ( .Q(WX2049), .DIN1(RESET), .DIN2(WX1986) );
  and2s1 U8045 ( .Q(WX2047), .DIN1(RESET), .DIN2(WX1984) );
  and2s1 U8046 ( .Q(WX2045), .DIN1(RESET), .DIN2(WX1982) );
  and2s1 U8047 ( .Q(WX2043), .DIN1(RESET), .DIN2(WX1980) );
  and2s1 U8048 ( .Q(WX2041), .DIN1(RESET), .DIN2(WX1978) );
  and2s1 U8049 ( .Q(WX2039), .DIN1(RESET), .DIN2(WX1976) );
  and2s1 U8050 ( .Q(WX2037), .DIN1(RESET), .DIN2(WX1974) );
  and2s1 U8051 ( .Q(WX2035), .DIN1(RESET), .DIN2(WX1972) );
  and2s1 U8052 ( .Q(WX2033), .DIN1(RESET), .DIN2(WX1970) );
  and2s1 U8053 ( .Q(WX2031), .DIN1(RESET), .DIN2(WX1968) );
  and2s1 U8054 ( .Q(WX2029), .DIN1(RESET), .DIN2(WX1966) );
  and2s1 U8055 ( .Q(WX2027), .DIN1(RESET), .DIN2(WX1964) );
  and2s1 U8056 ( .Q(WX2025), .DIN1(RESET), .DIN2(WX1962) );
  and2s1 U8057 ( .Q(WX2023), .DIN1(RESET), .DIN2(WX1960) );
  and2s1 U8058 ( .Q(WX2021), .DIN1(RESET), .DIN2(WX1958) );
  and2s1 U8059 ( .Q(WX2019), .DIN1(RESET), .DIN2(WX1956) );
  and2s1 U8060 ( .Q(WX2017), .DIN1(RESET), .DIN2(WX1954) );
  and2s1 U8061 ( .Q(WX2015), .DIN1(RESET), .DIN2(WX1952) );
  and2s1 U8062 ( .Q(WX2013), .DIN1(RESET), .DIN2(WX1950) );
  and2s1 U8063 ( .Q(WX2011), .DIN1(RESET), .DIN2(WX1948) );
  and2s1 U8064 ( .Q(WX2009), .DIN1(RESET), .DIN2(WX1946) );
  and2s1 U8065 ( .Q(WX2007), .DIN1(RESET), .DIN2(WX1944) );
  and2s1 U8066 ( .Q(WX2005), .DIN1(RESET), .DIN2(WX1942) );
  and2s1 U8067 ( .Q(WX2003), .DIN1(RESET), .DIN2(WX1940) );
  and2s1 U8068 ( .Q(WX2001), .DIN1(RESET), .DIN2(WX1938) );
  nnd4s1 U8069 ( .Q(WX1999), .DIN1(n5419), .DIN2(n5420), .DIN3(n5421), .DIN4(
        n5422) );
  nnd2s1 U8070 ( .Q(n5422), .DIN1(n3481), .DIN2(n5150) );
  xor2s1 U8071 ( .Q(n5150), .DIN1(n5423), .DIN2(n5424) );
  xor2s1 U8072 ( .Q(n5424), .DIN1(WX3357), .DIN2(n3189) );
  xor2s1 U8073 ( .Q(n5423), .DIN1(n3285), .DIN2(WX3421) );
  nnd2s1 U8074 ( .Q(n5421), .DIN1(n3437), .DIN2(n4339) );
  xor2s1 U8075 ( .Q(n4339), .DIN1(n5425), .DIN2(n5426) );
  xor2s1 U8076 ( .Q(n5426), .DIN1(n3029), .DIN2(WX2000) );
  xor2s1 U8077 ( .Q(n5425), .DIN1(n3286), .DIN2(WX2128) );
  nnd2s1 U8078 ( .Q(n5420), .DIN1(WX1840), .DIN2(n3500) );
  nnd2s1 U8079 ( .Q(n5419), .DIN1(CRC_OUT_8_0), .DIN2(n3532) );
  nnd4s1 U8080 ( .Q(WX1997), .DIN1(n5427), .DIN2(n5428), .DIN3(n5429), .DIN4(
        n5430) );
  nnd2s1 U8081 ( .Q(n5430), .DIN1(n3481), .DIN2(n5157) );
  xor2s1 U8082 ( .Q(n5157), .DIN1(n5431), .DIN2(n5432) );
  xor2s1 U8083 ( .Q(n5432), .DIN1(WX3355), .DIN2(n3190) );
  xor2s1 U8084 ( .Q(n5431), .DIN1(n3287), .DIN2(WX3419) );
  nnd2s1 U8085 ( .Q(n5429), .DIN1(n3437), .DIN2(n4346) );
  xor2s1 U8086 ( .Q(n4346), .DIN1(n5433), .DIN2(n5434) );
  xor2s1 U8087 ( .Q(n5434), .DIN1(n3030), .DIN2(WX1998) );
  xor2s1 U8088 ( .Q(n5433), .DIN1(n3288), .DIN2(WX2126) );
  nnd2s1 U8089 ( .Q(n5428), .DIN1(WX1838), .DIN2(n3500) );
  nnd2s1 U8090 ( .Q(n5427), .DIN1(CRC_OUT_8_1), .DIN2(n3532) );
  nnd4s1 U8091 ( .Q(WX1995), .DIN1(n5435), .DIN2(n5436), .DIN3(n5437), .DIN4(
        n5438) );
  nnd2s1 U8092 ( .Q(n5438), .DIN1(n3481), .DIN2(n5164) );
  xor2s1 U8093 ( .Q(n5164), .DIN1(n5439), .DIN2(n5440) );
  xor2s1 U8094 ( .Q(n5440), .DIN1(WX3353), .DIN2(n3191) );
  xor2s1 U8095 ( .Q(n5439), .DIN1(n3289), .DIN2(WX3417) );
  nnd2s1 U8096 ( .Q(n5437), .DIN1(n3437), .DIN2(n4353) );
  xor2s1 U8097 ( .Q(n4353), .DIN1(n5441), .DIN2(n5442) );
  xor2s1 U8098 ( .Q(n5442), .DIN1(n3031), .DIN2(WX1996) );
  xor2s1 U8099 ( .Q(n5441), .DIN1(n3290), .DIN2(WX2124) );
  nnd2s1 U8100 ( .Q(n5436), .DIN1(WX1836), .DIN2(n3500) );
  nnd2s1 U8101 ( .Q(n5435), .DIN1(CRC_OUT_8_2), .DIN2(n3532) );
  nnd4s1 U8102 ( .Q(WX1993), .DIN1(n5443), .DIN2(n5444), .DIN3(n5445), .DIN4(
        n5446) );
  nnd2s1 U8103 ( .Q(n5446), .DIN1(n3481), .DIN2(n5171) );
  xor2s1 U8104 ( .Q(n5171), .DIN1(n5447), .DIN2(n5448) );
  xor2s1 U8105 ( .Q(n5448), .DIN1(WX3351), .DIN2(n3192) );
  xor2s1 U8106 ( .Q(n5447), .DIN1(n3291), .DIN2(WX3415) );
  nnd2s1 U8107 ( .Q(n5445), .DIN1(n3437), .DIN2(n4360) );
  xor2s1 U8108 ( .Q(n4360), .DIN1(n5449), .DIN2(n5450) );
  xor2s1 U8109 ( .Q(n5450), .DIN1(n3032), .DIN2(WX1994) );
  xor2s1 U8110 ( .Q(n5449), .DIN1(n3292), .DIN2(WX2122) );
  nnd2s1 U8111 ( .Q(n5444), .DIN1(WX1834), .DIN2(n3500) );
  nnd2s1 U8112 ( .Q(n5443), .DIN1(CRC_OUT_8_3), .DIN2(n3532) );
  nnd4s1 U8113 ( .Q(WX1991), .DIN1(n5451), .DIN2(n5452), .DIN3(n5453), .DIN4(
        n5454) );
  nnd2s1 U8114 ( .Q(n5454), .DIN1(n3481), .DIN2(n5178) );
  xor2s1 U8115 ( .Q(n5178), .DIN1(n5455), .DIN2(n5456) );
  xor2s1 U8116 ( .Q(n5456), .DIN1(WX3349), .DIN2(n3193) );
  xor2s1 U8117 ( .Q(n5455), .DIN1(n3293), .DIN2(WX3413) );
  nnd2s1 U8118 ( .Q(n5453), .DIN1(n3437), .DIN2(n4367) );
  xor2s1 U8119 ( .Q(n4367), .DIN1(n5457), .DIN2(n5458) );
  xor2s1 U8120 ( .Q(n5458), .DIN1(n3033), .DIN2(WX1992) );
  xor2s1 U8121 ( .Q(n5457), .DIN1(n3294), .DIN2(WX2120) );
  nnd2s1 U8122 ( .Q(n5452), .DIN1(WX1832), .DIN2(n3499) );
  nnd2s1 U8123 ( .Q(n5451), .DIN1(CRC_OUT_8_4), .DIN2(n3531) );
  nnd4s1 U8124 ( .Q(WX1989), .DIN1(n5459), .DIN2(n5460), .DIN3(n5461), .DIN4(
        n5462) );
  nnd2s1 U8125 ( .Q(n5462), .DIN1(n3481), .DIN2(n5185) );
  xor2s1 U8126 ( .Q(n5185), .DIN1(n5463), .DIN2(n5464) );
  xor2s1 U8127 ( .Q(n5464), .DIN1(WX3347), .DIN2(n3194) );
  xor2s1 U8128 ( .Q(n5463), .DIN1(n3295), .DIN2(WX3411) );
  nnd2s1 U8129 ( .Q(n5461), .DIN1(n3437), .DIN2(n4374) );
  xor2s1 U8130 ( .Q(n4374), .DIN1(n5465), .DIN2(n5466) );
  xor2s1 U8131 ( .Q(n5466), .DIN1(n3034), .DIN2(WX1990) );
  xor2s1 U8132 ( .Q(n5465), .DIN1(n3296), .DIN2(WX2118) );
  nnd2s1 U8133 ( .Q(n5460), .DIN1(WX1830), .DIN2(n3499) );
  nnd2s1 U8134 ( .Q(n5459), .DIN1(CRC_OUT_8_5), .DIN2(n3531) );
  nnd4s1 U8135 ( .Q(WX1987), .DIN1(n5467), .DIN2(n5468), .DIN3(n5469), .DIN4(
        n5470) );
  nnd2s1 U8136 ( .Q(n5470), .DIN1(n3481), .DIN2(n5192) );
  xor2s1 U8137 ( .Q(n5192), .DIN1(n5471), .DIN2(n5472) );
  xor2s1 U8138 ( .Q(n5472), .DIN1(WX3345), .DIN2(n3195) );
  xor2s1 U8139 ( .Q(n5471), .DIN1(n3297), .DIN2(WX3409) );
  nnd2s1 U8140 ( .Q(n5469), .DIN1(n3437), .DIN2(n4381) );
  xor2s1 U8141 ( .Q(n4381), .DIN1(n5473), .DIN2(n5474) );
  xor2s1 U8142 ( .Q(n5474), .DIN1(n3035), .DIN2(WX1988) );
  xor2s1 U8143 ( .Q(n5473), .DIN1(n3298), .DIN2(WX2116) );
  nnd2s1 U8144 ( .Q(n5468), .DIN1(WX1828), .DIN2(n3499) );
  nnd2s1 U8145 ( .Q(n5467), .DIN1(CRC_OUT_8_6), .DIN2(n3531) );
  nnd4s1 U8146 ( .Q(WX1985), .DIN1(n5475), .DIN2(n5476), .DIN3(n5477), .DIN4(
        n5478) );
  nnd2s1 U8147 ( .Q(n5478), .DIN1(n3481), .DIN2(n5199) );
  xor2s1 U8148 ( .Q(n5199), .DIN1(n5479), .DIN2(n5480) );
  xor2s1 U8149 ( .Q(n5480), .DIN1(WX3343), .DIN2(n3196) );
  xor2s1 U8150 ( .Q(n5479), .DIN1(n3299), .DIN2(WX3407) );
  nnd2s1 U8151 ( .Q(n5477), .DIN1(n3437), .DIN2(n4388) );
  xor2s1 U8152 ( .Q(n4388), .DIN1(n5481), .DIN2(n5482) );
  xor2s1 U8153 ( .Q(n5482), .DIN1(n3036), .DIN2(WX1986) );
  xor2s1 U8154 ( .Q(n5481), .DIN1(n3300), .DIN2(WX2114) );
  nnd2s1 U8155 ( .Q(n5476), .DIN1(WX1826), .DIN2(n3499) );
  nnd2s1 U8156 ( .Q(n5475), .DIN1(CRC_OUT_8_7), .DIN2(n3531) );
  nnd4s1 U8157 ( .Q(WX1983), .DIN1(n5483), .DIN2(n5484), .DIN3(n5485), .DIN4(
        n5486) );
  nnd2s1 U8158 ( .Q(n5486), .DIN1(n3481), .DIN2(n5206) );
  xor2s1 U8159 ( .Q(n5206), .DIN1(n5487), .DIN2(n5488) );
  xor2s1 U8160 ( .Q(n5488), .DIN1(WX3341), .DIN2(n3197) );
  xor2s1 U8161 ( .Q(n5487), .DIN1(n3301), .DIN2(WX3405) );
  nnd2s1 U8162 ( .Q(n5485), .DIN1(n3437), .DIN2(n4395) );
  xor2s1 U8163 ( .Q(n4395), .DIN1(n5489), .DIN2(n5490) );
  xor2s1 U8164 ( .Q(n5490), .DIN1(n3037), .DIN2(WX1984) );
  xor2s1 U8165 ( .Q(n5489), .DIN1(n3302), .DIN2(WX2112) );
  nnd2s1 U8166 ( .Q(n5484), .DIN1(WX1824), .DIN2(n3499) );
  nnd2s1 U8167 ( .Q(n5483), .DIN1(CRC_OUT_8_8), .DIN2(n3531) );
  nnd4s1 U8168 ( .Q(WX1981), .DIN1(n5491), .DIN2(n5492), .DIN3(n5493), .DIN4(
        n5494) );
  nnd2s1 U8169 ( .Q(n5494), .DIN1(n3481), .DIN2(n5213) );
  xor2s1 U8170 ( .Q(n5213), .DIN1(n5495), .DIN2(n5496) );
  xor2s1 U8171 ( .Q(n5496), .DIN1(WX3339), .DIN2(n3198) );
  xor2s1 U8172 ( .Q(n5495), .DIN1(n3303), .DIN2(WX3403) );
  nnd2s1 U8173 ( .Q(n5493), .DIN1(n3437), .DIN2(n4402) );
  xor2s1 U8174 ( .Q(n4402), .DIN1(n5497), .DIN2(n5498) );
  xor2s1 U8175 ( .Q(n5498), .DIN1(n3038), .DIN2(WX1982) );
  xor2s1 U8176 ( .Q(n5497), .DIN1(n3304), .DIN2(WX2110) );
  nnd2s1 U8177 ( .Q(n5492), .DIN1(WX1822), .DIN2(n3499) );
  nnd2s1 U8178 ( .Q(n5491), .DIN1(CRC_OUT_8_9), .DIN2(n3531) );
  nnd4s1 U8179 ( .Q(WX1979), .DIN1(n5499), .DIN2(n5500), .DIN3(n5501), .DIN4(
        n5502) );
  nnd2s1 U8180 ( .Q(n5502), .DIN1(n3482), .DIN2(n5220) );
  xor2s1 U8181 ( .Q(n5220), .DIN1(n5503), .DIN2(n5504) );
  xor2s1 U8182 ( .Q(n5504), .DIN1(WX3337), .DIN2(n3199) );
  xor2s1 U8183 ( .Q(n5503), .DIN1(n3305), .DIN2(WX3401) );
  nnd2s1 U8184 ( .Q(n5501), .DIN1(n3437), .DIN2(n4409) );
  xor2s1 U8185 ( .Q(n4409), .DIN1(n5505), .DIN2(n5506) );
  xor2s1 U8186 ( .Q(n5506), .DIN1(n3039), .DIN2(WX1980) );
  xor2s1 U8187 ( .Q(n5505), .DIN1(n3306), .DIN2(WX2108) );
  nnd2s1 U8188 ( .Q(n5500), .DIN1(WX1820), .DIN2(n3499) );
  nnd2s1 U8189 ( .Q(n5499), .DIN1(CRC_OUT_8_10), .DIN2(n3531) );
  nnd4s1 U8190 ( .Q(WX1977), .DIN1(n5507), .DIN2(n5508), .DIN3(n5509), .DIN4(
        n5510) );
  nnd2s1 U8191 ( .Q(n5510), .DIN1(n3482), .DIN2(n5227) );
  xor2s1 U8192 ( .Q(n5227), .DIN1(n5511), .DIN2(n5512) );
  xor2s1 U8193 ( .Q(n5512), .DIN1(WX3335), .DIN2(n3200) );
  xor2s1 U8194 ( .Q(n5511), .DIN1(n3307), .DIN2(WX3399) );
  nnd2s1 U8195 ( .Q(n5509), .DIN1(n3437), .DIN2(n4416) );
  xor2s1 U8196 ( .Q(n4416), .DIN1(n5513), .DIN2(n5514) );
  xor2s1 U8197 ( .Q(n5514), .DIN1(n3040), .DIN2(WX1978) );
  xor2s1 U8198 ( .Q(n5513), .DIN1(n3308), .DIN2(WX2106) );
  nnd2s1 U8199 ( .Q(n5508), .DIN1(WX1818), .DIN2(n3499) );
  nnd2s1 U8200 ( .Q(n5507), .DIN1(CRC_OUT_8_11), .DIN2(n3531) );
  nnd4s1 U8201 ( .Q(WX1975), .DIN1(n5515), .DIN2(n5516), .DIN3(n5517), .DIN4(
        n5518) );
  nnd2s1 U8202 ( .Q(n5518), .DIN1(n3482), .DIN2(n5234) );
  xor2s1 U8203 ( .Q(n5234), .DIN1(n5519), .DIN2(n5520) );
  xor2s1 U8204 ( .Q(n5520), .DIN1(WX3333), .DIN2(n3201) );
  xor2s1 U8205 ( .Q(n5519), .DIN1(n3309), .DIN2(WX3397) );
  nnd2s1 U8206 ( .Q(n5517), .DIN1(n3436), .DIN2(n4423) );
  xor2s1 U8207 ( .Q(n4423), .DIN1(n5521), .DIN2(n5522) );
  xor2s1 U8208 ( .Q(n5522), .DIN1(n3041), .DIN2(WX1976) );
  xor2s1 U8209 ( .Q(n5521), .DIN1(n3310), .DIN2(WX2104) );
  nnd2s1 U8210 ( .Q(n5516), .DIN1(WX1816), .DIN2(n3499) );
  nnd2s1 U8211 ( .Q(n5515), .DIN1(CRC_OUT_8_12), .DIN2(n3531) );
  nnd4s1 U8212 ( .Q(WX1973), .DIN1(n5523), .DIN2(n5524), .DIN3(n5525), .DIN4(
        n5526) );
  nnd2s1 U8213 ( .Q(n5526), .DIN1(n3482), .DIN2(n5241) );
  xor2s1 U8214 ( .Q(n5241), .DIN1(n5527), .DIN2(n5528) );
  xor2s1 U8215 ( .Q(n5528), .DIN1(WX3331), .DIN2(n3202) );
  xor2s1 U8216 ( .Q(n5527), .DIN1(n3311), .DIN2(WX3395) );
  nnd2s1 U8217 ( .Q(n5525), .DIN1(n3436), .DIN2(n4430) );
  xor2s1 U8218 ( .Q(n4430), .DIN1(n5529), .DIN2(n5530) );
  xor2s1 U8219 ( .Q(n5530), .DIN1(n3042), .DIN2(WX1974) );
  xor2s1 U8220 ( .Q(n5529), .DIN1(n3312), .DIN2(WX2102) );
  nnd2s1 U8221 ( .Q(n5524), .DIN1(WX1814), .DIN2(n3499) );
  nnd2s1 U8222 ( .Q(n5523), .DIN1(CRC_OUT_8_13), .DIN2(n3531) );
  nnd4s1 U8223 ( .Q(WX1971), .DIN1(n5531), .DIN2(n5532), .DIN3(n5533), .DIN4(
        n5534) );
  nnd2s1 U8224 ( .Q(n5534), .DIN1(n3482), .DIN2(n5248) );
  xor2s1 U8225 ( .Q(n5248), .DIN1(n5535), .DIN2(n5536) );
  xor2s1 U8226 ( .Q(n5536), .DIN1(WX3329), .DIN2(n3203) );
  xor2s1 U8227 ( .Q(n5535), .DIN1(n3313), .DIN2(WX3393) );
  nnd2s1 U8228 ( .Q(n5533), .DIN1(n3436), .DIN2(n4437) );
  xor2s1 U8229 ( .Q(n4437), .DIN1(n5537), .DIN2(n5538) );
  xor2s1 U8230 ( .Q(n5538), .DIN1(n3043), .DIN2(WX1972) );
  xor2s1 U8231 ( .Q(n5537), .DIN1(n3314), .DIN2(WX2100) );
  nnd2s1 U8232 ( .Q(n5532), .DIN1(WX1812), .DIN2(n3499) );
  nnd2s1 U8233 ( .Q(n5531), .DIN1(CRC_OUT_8_14), .DIN2(n3531) );
  nnd4s1 U8234 ( .Q(WX1969), .DIN1(n5539), .DIN2(n5540), .DIN3(n5541), .DIN4(
        n5542) );
  nnd2s1 U8235 ( .Q(n5542), .DIN1(n3482), .DIN2(n5255) );
  xor2s1 U8236 ( .Q(n5255), .DIN1(n5543), .DIN2(n5544) );
  xor2s1 U8237 ( .Q(n5544), .DIN1(WX3327), .DIN2(n3204) );
  xor2s1 U8238 ( .Q(n5543), .DIN1(n3315), .DIN2(WX3391) );
  nnd2s1 U8239 ( .Q(n5541), .DIN1(n3436), .DIN2(n4444) );
  xor2s1 U8240 ( .Q(n4444), .DIN1(n5545), .DIN2(n5546) );
  xor2s1 U8241 ( .Q(n5546), .DIN1(n3044), .DIN2(WX1970) );
  xor2s1 U8242 ( .Q(n5545), .DIN1(n3316), .DIN2(WX2098) );
  nnd2s1 U8243 ( .Q(n5540), .DIN1(WX1810), .DIN2(n3499) );
  nnd2s1 U8244 ( .Q(n5539), .DIN1(CRC_OUT_8_15), .DIN2(n3531) );
  nnd4s1 U8245 ( .Q(WX1967), .DIN1(n5547), .DIN2(n5548), .DIN3(n5549), .DIN4(
        n5550) );
  nnd2s1 U8246 ( .Q(n5550), .DIN1(n3482), .DIN2(n5263) );
  xor2s1 U8247 ( .Q(n5263), .DIN1(n5551), .DIN2(n5552) );
  xor2s1 U8248 ( .Q(n5552), .DIN1(n3570), .DIN2(WX3261) );
  xor2s1 U8249 ( .Q(n5551), .DIN1(n3045), .DIN2(n5553) );
  xor2s1 U8250 ( .Q(n5553), .DIN1(WX3453), .DIN2(WX3389) );
  nnd2s1 U8251 ( .Q(n5549), .DIN1(n3436), .DIN2(n4451) );
  xor2s1 U8252 ( .Q(n4451), .DIN1(n5554), .DIN2(n5555) );
  xor2s1 U8253 ( .Q(n5555), .DIN1(n3570), .DIN2(WX1968) );
  xor2s1 U8254 ( .Q(n5554), .DIN1(n3046), .DIN2(n5556) );
  xor2s1 U8255 ( .Q(n5556), .DIN1(WX2160), .DIN2(WX2096) );
  nnd2s1 U8256 ( .Q(n5548), .DIN1(WX1808), .DIN2(n3498) );
  nnd2s1 U8257 ( .Q(n5547), .DIN1(CRC_OUT_8_16), .DIN2(n3530) );
  nnd4s1 U8258 ( .Q(WX1965), .DIN1(n5557), .DIN2(n5558), .DIN3(n5559), .DIN4(
        n5560) );
  nnd2s1 U8259 ( .Q(n5560), .DIN1(n3482), .DIN2(n5271) );
  xor2s1 U8260 ( .Q(n5271), .DIN1(n5561), .DIN2(n5562) );
  xor2s1 U8261 ( .Q(n5562), .DIN1(n3570), .DIN2(WX3259) );
  xor2s1 U8262 ( .Q(n5561), .DIN1(n3047), .DIN2(n5563) );
  xor2s1 U8263 ( .Q(n5563), .DIN1(WX3451), .DIN2(WX3387) );
  nnd2s1 U8264 ( .Q(n5559), .DIN1(n3436), .DIN2(n4458) );
  xor2s1 U8265 ( .Q(n4458), .DIN1(n5564), .DIN2(n5565) );
  xor2s1 U8266 ( .Q(n5565), .DIN1(n3571), .DIN2(WX1966) );
  xor2s1 U8267 ( .Q(n5564), .DIN1(n3048), .DIN2(n5566) );
  xor2s1 U8268 ( .Q(n5566), .DIN1(WX2158), .DIN2(WX2094) );
  nnd2s1 U8269 ( .Q(n5558), .DIN1(WX1806), .DIN2(n3498) );
  nnd2s1 U8270 ( .Q(n5557), .DIN1(CRC_OUT_8_17), .DIN2(n3530) );
  nnd4s1 U8271 ( .Q(WX1963), .DIN1(n5567), .DIN2(n5568), .DIN3(n5569), .DIN4(
        n5570) );
  nnd2s1 U8272 ( .Q(n5570), .DIN1(n3482), .DIN2(n5279) );
  xor2s1 U8273 ( .Q(n5279), .DIN1(n5571), .DIN2(n5572) );
  xor2s1 U8274 ( .Q(n5572), .DIN1(n3571), .DIN2(WX3257) );
  xor2s1 U8275 ( .Q(n5571), .DIN1(n3049), .DIN2(n5573) );
  xor2s1 U8276 ( .Q(n5573), .DIN1(WX3449), .DIN2(WX3385) );
  nnd2s1 U8277 ( .Q(n5569), .DIN1(n3436), .DIN2(n4465) );
  xor2s1 U8278 ( .Q(n4465), .DIN1(n5574), .DIN2(n5575) );
  xor2s1 U8279 ( .Q(n5575), .DIN1(n3571), .DIN2(WX1964) );
  xor2s1 U8280 ( .Q(n5574), .DIN1(n3050), .DIN2(n5576) );
  xor2s1 U8281 ( .Q(n5576), .DIN1(WX2156), .DIN2(WX2092) );
  nnd2s1 U8282 ( .Q(n5568), .DIN1(WX1804), .DIN2(n3498) );
  nnd2s1 U8283 ( .Q(n5567), .DIN1(CRC_OUT_8_18), .DIN2(n3530) );
  nnd4s1 U8284 ( .Q(WX1961), .DIN1(n5577), .DIN2(n5578), .DIN3(n5579), .DIN4(
        n5580) );
  nnd2s1 U8285 ( .Q(n5580), .DIN1(n3482), .DIN2(n5287) );
  xor2s1 U8286 ( .Q(n5287), .DIN1(n5581), .DIN2(n5582) );
  xor2s1 U8287 ( .Q(n5582), .DIN1(n3571), .DIN2(WX3255) );
  xor2s1 U8288 ( .Q(n5581), .DIN1(n3051), .DIN2(n5583) );
  xor2s1 U8289 ( .Q(n5583), .DIN1(WX3447), .DIN2(WX3383) );
  nnd2s1 U8290 ( .Q(n5579), .DIN1(n3436), .DIN2(n4472) );
  xor2s1 U8291 ( .Q(n4472), .DIN1(n5584), .DIN2(n5585) );
  xor2s1 U8292 ( .Q(n5585), .DIN1(n3571), .DIN2(WX1962) );
  xor2s1 U8293 ( .Q(n5584), .DIN1(n3052), .DIN2(n5586) );
  xor2s1 U8294 ( .Q(n5586), .DIN1(WX2154), .DIN2(WX2090) );
  nnd2s1 U8295 ( .Q(n5578), .DIN1(WX1802), .DIN2(n3498) );
  nnd2s1 U8296 ( .Q(n5577), .DIN1(CRC_OUT_8_19), .DIN2(n3530) );
  nnd4s1 U8297 ( .Q(WX1959), .DIN1(n5587), .DIN2(n5588), .DIN3(n5589), .DIN4(
        n5590) );
  nnd2s1 U8298 ( .Q(n5590), .DIN1(n3482), .DIN2(n5295) );
  xor2s1 U8299 ( .Q(n5295), .DIN1(n5591), .DIN2(n5592) );
  xor2s1 U8300 ( .Q(n5592), .DIN1(n3571), .DIN2(WX3253) );
  xor2s1 U8301 ( .Q(n5591), .DIN1(n3053), .DIN2(n5593) );
  xor2s1 U8302 ( .Q(n5593), .DIN1(WX3445), .DIN2(WX3381) );
  nnd2s1 U8303 ( .Q(n5589), .DIN1(n3436), .DIN2(n4479) );
  xor2s1 U8304 ( .Q(n4479), .DIN1(n5594), .DIN2(n5595) );
  xor2s1 U8305 ( .Q(n5595), .DIN1(n3571), .DIN2(WX1960) );
  xor2s1 U8306 ( .Q(n5594), .DIN1(n3054), .DIN2(n5596) );
  xor2s1 U8307 ( .Q(n5596), .DIN1(WX2152), .DIN2(WX2088) );
  nnd2s1 U8308 ( .Q(n5588), .DIN1(WX1800), .DIN2(n3498) );
  nnd2s1 U8309 ( .Q(n5587), .DIN1(CRC_OUT_8_20), .DIN2(n3530) );
  nnd4s1 U8310 ( .Q(WX1957), .DIN1(n5597), .DIN2(n5598), .DIN3(n5599), .DIN4(
        n5600) );
  nnd2s1 U8311 ( .Q(n5600), .DIN1(n3482), .DIN2(n5303) );
  xor2s1 U8312 ( .Q(n5303), .DIN1(n5601), .DIN2(n5602) );
  xor2s1 U8313 ( .Q(n5602), .DIN1(n3572), .DIN2(WX3251) );
  xor2s1 U8314 ( .Q(n5601), .DIN1(n3055), .DIN2(n5603) );
  xor2s1 U8315 ( .Q(n5603), .DIN1(WX3443), .DIN2(WX3379) );
  nnd2s1 U8316 ( .Q(n5599), .DIN1(n3436), .DIN2(n4486) );
  xor2s1 U8317 ( .Q(n4486), .DIN1(n5604), .DIN2(n5605) );
  xor2s1 U8318 ( .Q(n5605), .DIN1(n3572), .DIN2(WX1958) );
  xor2s1 U8319 ( .Q(n5604), .DIN1(n3056), .DIN2(n5606) );
  xor2s1 U8320 ( .Q(n5606), .DIN1(WX2150), .DIN2(WX2086) );
  nnd2s1 U8321 ( .Q(n5598), .DIN1(WX1798), .DIN2(n3498) );
  nnd2s1 U8322 ( .Q(n5597), .DIN1(CRC_OUT_8_21), .DIN2(n3530) );
  nnd4s1 U8323 ( .Q(WX1955), .DIN1(n5607), .DIN2(n5608), .DIN3(n5609), .DIN4(
        n5610) );
  nnd2s1 U8324 ( .Q(n5610), .DIN1(n3482), .DIN2(n5311) );
  xor2s1 U8325 ( .Q(n5311), .DIN1(n5611), .DIN2(n5612) );
  xor2s1 U8326 ( .Q(n5612), .DIN1(n3572), .DIN2(WX3249) );
  xor2s1 U8327 ( .Q(n5611), .DIN1(n3057), .DIN2(n5613) );
  xor2s1 U8328 ( .Q(n5613), .DIN1(WX3441), .DIN2(WX3377) );
  nnd2s1 U8329 ( .Q(n5609), .DIN1(n3436), .DIN2(n4493) );
  xor2s1 U8330 ( .Q(n4493), .DIN1(n5614), .DIN2(n5615) );
  xor2s1 U8331 ( .Q(n5615), .DIN1(n3572), .DIN2(WX1956) );
  xor2s1 U8332 ( .Q(n5614), .DIN1(n3058), .DIN2(n5616) );
  xor2s1 U8333 ( .Q(n5616), .DIN1(WX2148), .DIN2(WX2084) );
  nnd2s1 U8334 ( .Q(n5608), .DIN1(WX1796), .DIN2(n3498) );
  nnd2s1 U8335 ( .Q(n5607), .DIN1(CRC_OUT_8_22), .DIN2(n3530) );
  nnd4s1 U8336 ( .Q(WX1953), .DIN1(n5617), .DIN2(n5618), .DIN3(n5619), .DIN4(
        n5620) );
  nnd2s1 U8337 ( .Q(n5620), .DIN1(n3483), .DIN2(n5319) );
  xor2s1 U8338 ( .Q(n5319), .DIN1(n5621), .DIN2(n5622) );
  xor2s1 U8339 ( .Q(n5622), .DIN1(n3572), .DIN2(WX3247) );
  xor2s1 U8340 ( .Q(n5621), .DIN1(n3059), .DIN2(n5623) );
  xor2s1 U8341 ( .Q(n5623), .DIN1(WX3439), .DIN2(WX3375) );
  nnd2s1 U8342 ( .Q(n5619), .DIN1(n3436), .DIN2(n4500) );
  xor2s1 U8343 ( .Q(n4500), .DIN1(n5624), .DIN2(n5625) );
  xor2s1 U8344 ( .Q(n5625), .DIN1(n3572), .DIN2(WX1954) );
  xor2s1 U8345 ( .Q(n5624), .DIN1(n3060), .DIN2(n5626) );
  xor2s1 U8346 ( .Q(n5626), .DIN1(WX2146), .DIN2(WX2082) );
  nnd2s1 U8347 ( .Q(n5618), .DIN1(WX1794), .DIN2(n3498) );
  nnd2s1 U8348 ( .Q(n5617), .DIN1(CRC_OUT_8_23), .DIN2(n3530) );
  nnd4s1 U8349 ( .Q(WX1951), .DIN1(n5627), .DIN2(n5628), .DIN3(n5629), .DIN4(
        n5630) );
  nnd2s1 U8350 ( .Q(n5630), .DIN1(n3483), .DIN2(n5327) );
  xor2s1 U8351 ( .Q(n5327), .DIN1(n5631), .DIN2(n5632) );
  xor2s1 U8352 ( .Q(n5632), .DIN1(n3572), .DIN2(WX3245) );
  xor2s1 U8353 ( .Q(n5631), .DIN1(n3061), .DIN2(n5633) );
  xor2s1 U8354 ( .Q(n5633), .DIN1(WX3437), .DIN2(WX3373) );
  nnd2s1 U8355 ( .Q(n5629), .DIN1(n3436), .DIN2(n4507) );
  xor2s1 U8356 ( .Q(n4507), .DIN1(n5634), .DIN2(n5635) );
  xor2s1 U8357 ( .Q(n5635), .DIN1(n3573), .DIN2(WX1952) );
  xor2s1 U8358 ( .Q(n5634), .DIN1(n3062), .DIN2(n5636) );
  xor2s1 U8359 ( .Q(n5636), .DIN1(WX2144), .DIN2(WX2080) );
  nnd2s1 U8360 ( .Q(n5628), .DIN1(WX1792), .DIN2(n3498) );
  nnd2s1 U8361 ( .Q(n5627), .DIN1(CRC_OUT_8_24), .DIN2(n3530) );
  nnd4s1 U8362 ( .Q(WX1949), .DIN1(n5637), .DIN2(n5638), .DIN3(n5639), .DIN4(
        n5640) );
  nnd2s1 U8363 ( .Q(n5640), .DIN1(n3483), .DIN2(n5335) );
  xor2s1 U8364 ( .Q(n5335), .DIN1(n5641), .DIN2(n5642) );
  xor2s1 U8365 ( .Q(n5642), .DIN1(n3573), .DIN2(WX3243) );
  xor2s1 U8366 ( .Q(n5641), .DIN1(n3063), .DIN2(n5643) );
  xor2s1 U8367 ( .Q(n5643), .DIN1(WX3435), .DIN2(WX3371) );
  nnd2s1 U8368 ( .Q(n5639), .DIN1(n3435), .DIN2(n4514) );
  xor2s1 U8369 ( .Q(n4514), .DIN1(n5644), .DIN2(n5645) );
  xor2s1 U8370 ( .Q(n5645), .DIN1(n3573), .DIN2(WX1950) );
  xor2s1 U8371 ( .Q(n5644), .DIN1(n3064), .DIN2(n5646) );
  xor2s1 U8372 ( .Q(n5646), .DIN1(WX2142), .DIN2(WX2078) );
  nnd2s1 U8373 ( .Q(n5638), .DIN1(WX1790), .DIN2(n3498) );
  nnd2s1 U8374 ( .Q(n5637), .DIN1(CRC_OUT_8_25), .DIN2(n3530) );
  nnd4s1 U8375 ( .Q(WX1947), .DIN1(n5647), .DIN2(n5648), .DIN3(n5649), .DIN4(
        n5650) );
  nnd2s1 U8376 ( .Q(n5650), .DIN1(n3483), .DIN2(n5343) );
  xor2s1 U8377 ( .Q(n5343), .DIN1(n5651), .DIN2(n5652) );
  xor2s1 U8378 ( .Q(n5652), .DIN1(n3573), .DIN2(WX3241) );
  xor2s1 U8379 ( .Q(n5651), .DIN1(n3065), .DIN2(n5653) );
  xor2s1 U8380 ( .Q(n5653), .DIN1(WX3433), .DIN2(WX3369) );
  nnd2s1 U8381 ( .Q(n5649), .DIN1(n3435), .DIN2(n4521) );
  xor2s1 U8382 ( .Q(n4521), .DIN1(n5654), .DIN2(n5655) );
  xor2s1 U8383 ( .Q(n5655), .DIN1(n3573), .DIN2(WX1948) );
  xor2s1 U8384 ( .Q(n5654), .DIN1(n3066), .DIN2(n5656) );
  xor2s1 U8385 ( .Q(n5656), .DIN1(WX2140), .DIN2(WX2076) );
  nnd2s1 U8386 ( .Q(n5648), .DIN1(WX1788), .DIN2(n3498) );
  nnd2s1 U8387 ( .Q(n5647), .DIN1(CRC_OUT_8_26), .DIN2(n3530) );
  nnd4s1 U8388 ( .Q(WX1945), .DIN1(n5657), .DIN2(n5658), .DIN3(n5659), .DIN4(
        n5660) );
  nnd2s1 U8389 ( .Q(n5660), .DIN1(n3483), .DIN2(n5351) );
  xor2s1 U8390 ( .Q(n5351), .DIN1(n5661), .DIN2(n5662) );
  xor2s1 U8391 ( .Q(n5662), .DIN1(n3573), .DIN2(WX3239) );
  xor2s1 U8392 ( .Q(n5661), .DIN1(n3067), .DIN2(n5663) );
  xor2s1 U8393 ( .Q(n5663), .DIN1(WX3431), .DIN2(WX3367) );
  nnd2s1 U8394 ( .Q(n5659), .DIN1(n3435), .DIN2(n4528) );
  xor2s1 U8395 ( .Q(n4528), .DIN1(n5664), .DIN2(n5665) );
  xor2s1 U8396 ( .Q(n5665), .DIN1(n3573), .DIN2(WX1946) );
  xor2s1 U8397 ( .Q(n5664), .DIN1(n3068), .DIN2(n5666) );
  xor2s1 U8398 ( .Q(n5666), .DIN1(WX2138), .DIN2(WX2074) );
  nnd2s1 U8399 ( .Q(n5658), .DIN1(WX1786), .DIN2(n3498) );
  nnd2s1 U8400 ( .Q(n5657), .DIN1(CRC_OUT_8_27), .DIN2(n3530) );
  nnd4s1 U8401 ( .Q(WX1943), .DIN1(n5667), .DIN2(n5668), .DIN3(n5669), .DIN4(
        n5670) );
  nnd2s1 U8402 ( .Q(n5670), .DIN1(n3483), .DIN2(n5359) );
  xor2s1 U8403 ( .Q(n5359), .DIN1(n5671), .DIN2(n5672) );
  xor2s1 U8404 ( .Q(n5672), .DIN1(n3574), .DIN2(WX3237) );
  xor2s1 U8405 ( .Q(n5671), .DIN1(n3069), .DIN2(n5673) );
  xor2s1 U8406 ( .Q(n5673), .DIN1(WX3429), .DIN2(WX3365) );
  nnd2s1 U8407 ( .Q(n5669), .DIN1(n3435), .DIN2(n4535) );
  xor2s1 U8408 ( .Q(n4535), .DIN1(n5674), .DIN2(n5675) );
  xor2s1 U8409 ( .Q(n5675), .DIN1(n3574), .DIN2(WX1944) );
  xor2s1 U8410 ( .Q(n5674), .DIN1(n3070), .DIN2(n5676) );
  xor2s1 U8411 ( .Q(n5676), .DIN1(WX2136), .DIN2(WX2072) );
  nnd2s1 U8412 ( .Q(n5668), .DIN1(WX1784), .DIN2(n3497) );
  nnd2s1 U8413 ( .Q(n5667), .DIN1(CRC_OUT_8_28), .DIN2(n3529) );
  nnd4s1 U8414 ( .Q(WX1941), .DIN1(n5677), .DIN2(n5678), .DIN3(n5679), .DIN4(
        n5680) );
  nnd2s1 U8415 ( .Q(n5680), .DIN1(n3483), .DIN2(n5367) );
  xor2s1 U8416 ( .Q(n5367), .DIN1(n5681), .DIN2(n5682) );
  xor2s1 U8417 ( .Q(n5682), .DIN1(n3574), .DIN2(WX3235) );
  xor2s1 U8418 ( .Q(n5681), .DIN1(n3071), .DIN2(n5683) );
  xor2s1 U8419 ( .Q(n5683), .DIN1(WX3427), .DIN2(WX3363) );
  nnd2s1 U8420 ( .Q(n5679), .DIN1(n3435), .DIN2(n4552) );
  xor2s1 U8421 ( .Q(n4552), .DIN1(n5684), .DIN2(n5685) );
  xor2s1 U8422 ( .Q(n5685), .DIN1(n3574), .DIN2(WX1942) );
  xor2s1 U8423 ( .Q(n5684), .DIN1(n3072), .DIN2(n5686) );
  xor2s1 U8424 ( .Q(n5686), .DIN1(WX2134), .DIN2(WX2070) );
  nnd2s1 U8425 ( .Q(n5678), .DIN1(WX1782), .DIN2(n3497) );
  nnd2s1 U8426 ( .Q(n5677), .DIN1(CRC_OUT_8_29), .DIN2(n3529) );
  nnd4s1 U8427 ( .Q(WX1939), .DIN1(n5687), .DIN2(n5688), .DIN3(n5689), .DIN4(
        n5690) );
  nnd2s1 U8428 ( .Q(n5690), .DIN1(n3483), .DIN2(n5375) );
  xor2s1 U8429 ( .Q(n5375), .DIN1(n5691), .DIN2(n5692) );
  xor2s1 U8430 ( .Q(n5692), .DIN1(n3574), .DIN2(WX3233) );
  xor2s1 U8431 ( .Q(n5691), .DIN1(n3073), .DIN2(n5693) );
  xor2s1 U8432 ( .Q(n5693), .DIN1(WX3425), .DIN2(WX3361) );
  nnd2s1 U8433 ( .Q(n5689), .DIN1(n3435), .DIN2(n4570) );
  xor2s1 U8434 ( .Q(n4570), .DIN1(n5694), .DIN2(n5695) );
  xor2s1 U8435 ( .Q(n5695), .DIN1(n3574), .DIN2(WX1940) );
  xor2s1 U8436 ( .Q(n5694), .DIN1(n3074), .DIN2(n5696) );
  xor2s1 U8437 ( .Q(n5696), .DIN1(WX2132), .DIN2(WX2068) );
  nnd2s1 U8438 ( .Q(n5688), .DIN1(WX1780), .DIN2(n3497) );
  nnd2s1 U8439 ( .Q(n5687), .DIN1(CRC_OUT_8_30), .DIN2(n3529) );
  nnd4s1 U8440 ( .Q(WX1937), .DIN1(n5697), .DIN2(n5698), .DIN3(n5699), .DIN4(
        n5700) );
  nnd2s1 U8441 ( .Q(n5700), .DIN1(n3483), .DIN2(n5383) );
  xor2s1 U8442 ( .Q(n5383), .DIN1(n5701), .DIN2(n5702) );
  xor2s1 U8443 ( .Q(n5702), .DIN1(n3574), .DIN2(WX3231) );
  xor2s1 U8444 ( .Q(n5701), .DIN1(n3075), .DIN2(n5703) );
  xor2s1 U8445 ( .Q(n5703), .DIN1(WX3423), .DIN2(WX3359) );
  nnd2s1 U8446 ( .Q(n5699), .DIN1(n3435), .DIN2(n4589) );
  xor2s1 U8447 ( .Q(n4589), .DIN1(n5704), .DIN2(n5705) );
  xor2s1 U8448 ( .Q(n5705), .DIN1(n3575), .DIN2(WX1938) );
  xor2s1 U8449 ( .Q(n5704), .DIN1(n3076), .DIN2(n5706) );
  xor2s1 U8450 ( .Q(n5706), .DIN1(WX2130), .DIN2(WX2066) );
  nnd2s1 U8451 ( .Q(n5698), .DIN1(WX1778), .DIN2(n3497) );
  nnd2s1 U8452 ( .Q(n5697), .DIN1(CRC_OUT_8_31), .DIN2(n3529) );
  nor2s1 U8453 ( .Q(WX1839), .DIN1(WX1778), .DIN2(n3363) );
  and2s1 U8454 ( .Q(WX1837), .DIN1(RESET), .DIN2(WX1840) );
  and2s1 U8455 ( .Q(WX1835), .DIN1(RESET), .DIN2(WX1838) );
  and2s1 U8456 ( .Q(WX1833), .DIN1(RESET), .DIN2(WX1836) );
  and2s1 U8457 ( .Q(WX1831), .DIN1(RESET), .DIN2(WX1834) );
  and2s1 U8458 ( .Q(WX1829), .DIN1(RESET), .DIN2(WX1832) );
  and2s1 U8459 ( .Q(WX1827), .DIN1(RESET), .DIN2(WX1830) );
  and2s1 U8460 ( .Q(WX1825), .DIN1(RESET), .DIN2(WX1828) );
  and2s1 U8461 ( .Q(WX1823), .DIN1(RESET), .DIN2(WX1826) );
  and2s1 U8462 ( .Q(WX1821), .DIN1(RESET), .DIN2(WX1824) );
  and2s1 U8463 ( .Q(WX1819), .DIN1(RESET), .DIN2(WX1822) );
  and2s1 U8464 ( .Q(WX1817), .DIN1(RESET), .DIN2(WX1820) );
  and2s1 U8465 ( .Q(WX1815), .DIN1(RESET), .DIN2(WX1818) );
  and2s1 U8466 ( .Q(WX1813), .DIN1(RESET), .DIN2(WX1816) );
  and2s1 U8467 ( .Q(WX1811), .DIN1(RESET), .DIN2(WX1814) );
  and2s1 U8468 ( .Q(WX1809), .DIN1(RESET), .DIN2(WX1812) );
  and2s1 U8469 ( .Q(WX1807), .DIN1(RESET), .DIN2(WX1810) );
  and2s1 U8470 ( .Q(WX1805), .DIN1(RESET), .DIN2(WX1808) );
  and2s1 U8471 ( .Q(WX1803), .DIN1(RESET), .DIN2(WX1806) );
  and2s1 U8472 ( .Q(WX1801), .DIN1(RESET), .DIN2(WX1804) );
  and2s1 U8473 ( .Q(WX1799), .DIN1(RESET), .DIN2(WX1802) );
  and2s1 U8474 ( .Q(WX1797), .DIN1(RESET), .DIN2(WX1800) );
  and2s1 U8475 ( .Q(WX1795), .DIN1(RESET), .DIN2(WX1798) );
  and2s1 U8476 ( .Q(WX1793), .DIN1(RESET), .DIN2(WX1796) );
  and2s1 U8477 ( .Q(WX1791), .DIN1(RESET), .DIN2(WX1794) );
  and2s1 U8478 ( .Q(WX1789), .DIN1(RESET), .DIN2(WX1792) );
  and2s1 U8479 ( .Q(WX1787), .DIN1(RESET), .DIN2(WX1790) );
  and2s1 U8480 ( .Q(WX1785), .DIN1(RESET), .DIN2(WX1788) );
  and2s1 U8481 ( .Q(WX1783), .DIN1(RESET), .DIN2(WX1786) );
  and2s1 U8482 ( .Q(WX1781), .DIN1(RESET), .DIN2(WX1784) );
  and2s1 U8483 ( .Q(WX1779), .DIN1(RESET), .DIN2(WX1782) );
  and2s1 U8484 ( .Q(WX1777), .DIN1(RESET), .DIN2(WX1780) );
  nor2s1 U8485 ( .Q(WX1326), .DIN1(n3391), .DIN2(n5707) );
  xor2s1 U8486 ( .Q(n5707), .DIN1(WX837), .DIN2(CRC_OUT_9_30) );
  nor2s1 U8487 ( .Q(WX1324), .DIN1(n3391), .DIN2(n5708) );
  xor2s1 U8488 ( .Q(n5708), .DIN1(WX839), .DIN2(CRC_OUT_9_29) );
  nor2s1 U8489 ( .Q(WX1322), .DIN1(n3392), .DIN2(n5709) );
  xor2s1 U8490 ( .Q(n5709), .DIN1(WX841), .DIN2(CRC_OUT_9_28) );
  nor2s1 U8491 ( .Q(WX1320), .DIN1(n3392), .DIN2(n5710) );
  xor2s1 U8492 ( .Q(n5710), .DIN1(WX843), .DIN2(CRC_OUT_9_27) );
  nor2s1 U8493 ( .Q(WX1318), .DIN1(n3392), .DIN2(n5711) );
  xor2s1 U8494 ( .Q(n5711), .DIN1(WX845), .DIN2(CRC_OUT_9_26) );
  nor2s1 U8495 ( .Q(WX1316), .DIN1(n3392), .DIN2(n5712) );
  xor2s1 U8496 ( .Q(n5712), .DIN1(WX847), .DIN2(CRC_OUT_9_25) );
  nor2s1 U8497 ( .Q(WX1314), .DIN1(n3392), .DIN2(n5713) );
  xor2s1 U8498 ( .Q(n5713), .DIN1(WX849), .DIN2(CRC_OUT_9_24) );
  nor2s1 U8499 ( .Q(WX1312), .DIN1(n3392), .DIN2(n5714) );
  xor2s1 U8500 ( .Q(n5714), .DIN1(WX851), .DIN2(CRC_OUT_9_23) );
  nor2s1 U8501 ( .Q(WX1310), .DIN1(n3392), .DIN2(n5715) );
  xor2s1 U8502 ( .Q(n5715), .DIN1(WX853), .DIN2(CRC_OUT_9_22) );
  nor2s1 U8503 ( .Q(WX1308), .DIN1(n3392), .DIN2(n5716) );
  xor2s1 U8504 ( .Q(n5716), .DIN1(WX855), .DIN2(CRC_OUT_9_21) );
  nor2s1 U8505 ( .Q(WX1306), .DIN1(n3392), .DIN2(n5717) );
  xor2s1 U8506 ( .Q(n5717), .DIN1(WX857), .DIN2(CRC_OUT_9_20) );
  nor2s1 U8507 ( .Q(WX1304), .DIN1(n3392), .DIN2(n5718) );
  xor2s1 U8508 ( .Q(n5718), .DIN1(WX859), .DIN2(CRC_OUT_9_19) );
  nor2s1 U8509 ( .Q(WX1302), .DIN1(n3393), .DIN2(n5719) );
  xor2s1 U8510 ( .Q(n5719), .DIN1(WX861), .DIN2(CRC_OUT_9_18) );
  nor2s1 U8511 ( .Q(WX1300), .DIN1(n3393), .DIN2(n5720) );
  xor2s1 U8512 ( .Q(n5720), .DIN1(WX863), .DIN2(CRC_OUT_9_17) );
  nor2s1 U8513 ( .Q(WX1298), .DIN1(n3393), .DIN2(n5721) );
  xor2s1 U8514 ( .Q(n5721), .DIN1(WX865), .DIN2(CRC_OUT_9_16) );
  nor2s1 U8515 ( .Q(WX1296), .DIN1(n3393), .DIN2(n5722) );
  xor2s1 U8516 ( .Q(n5722), .DIN1(CRC_OUT_9_15), .DIN2(n5723) );
  xor2s1 U8517 ( .Q(n5723), .DIN1(WX867), .DIN2(CRC_OUT_9_31) );
  nor2s1 U8518 ( .Q(WX1294), .DIN1(n3393), .DIN2(n5724) );
  xor2s1 U8519 ( .Q(n5724), .DIN1(WX869), .DIN2(CRC_OUT_9_14) );
  nor2s1 U8520 ( .Q(WX1292), .DIN1(n3393), .DIN2(n5725) );
  xor2s1 U8521 ( .Q(n5725), .DIN1(WX871), .DIN2(CRC_OUT_9_13) );
  nor2s1 U8522 ( .Q(WX1290), .DIN1(n3393), .DIN2(n5726) );
  xor2s1 U8523 ( .Q(n5726), .DIN1(WX873), .DIN2(CRC_OUT_9_12) );
  nor2s1 U8524 ( .Q(WX1288), .DIN1(n3393), .DIN2(n5727) );
  xor2s1 U8525 ( .Q(n5727), .DIN1(WX875), .DIN2(CRC_OUT_9_11) );
  nor2s1 U8526 ( .Q(WX1286), .DIN1(n3393), .DIN2(n5728) );
  xor2s1 U8527 ( .Q(n5728), .DIN1(CRC_OUT_9_10), .DIN2(n5729) );
  xor2s1 U8528 ( .Q(n5729), .DIN1(WX877), .DIN2(CRC_OUT_9_31) );
  nor2s1 U8529 ( .Q(WX1284), .DIN1(n3393), .DIN2(n5730) );
  xor2s1 U8530 ( .Q(n5730), .DIN1(WX879), .DIN2(CRC_OUT_9_9) );
  nor2s1 U8531 ( .Q(WX1282), .DIN1(n3394), .DIN2(n5731) );
  xor2s1 U8532 ( .Q(n5731), .DIN1(WX881), .DIN2(CRC_OUT_9_8) );
  nor2s1 U8533 ( .Q(WX1280), .DIN1(n3394), .DIN2(n5732) );
  xor2s1 U8534 ( .Q(n5732), .DIN1(WX883), .DIN2(CRC_OUT_9_7) );
  nor2s1 U8535 ( .Q(WX1278), .DIN1(n3394), .DIN2(n5733) );
  xor2s1 U8536 ( .Q(n5733), .DIN1(WX885), .DIN2(CRC_OUT_9_6) );
  nor2s1 U8537 ( .Q(WX1276), .DIN1(n3394), .DIN2(n5734) );
  xor2s1 U8538 ( .Q(n5734), .DIN1(WX887), .DIN2(CRC_OUT_9_5) );
  nor2s1 U8539 ( .Q(WX1274), .DIN1(n3394), .DIN2(n5735) );
  xor2s1 U8540 ( .Q(n5735), .DIN1(WX889), .DIN2(CRC_OUT_9_4) );
  nor2s1 U8541 ( .Q(WX1272), .DIN1(n3394), .DIN2(n5736) );
  xor2s1 U8542 ( .Q(n5736), .DIN1(CRC_OUT_9_3), .DIN2(n5737) );
  xor2s1 U8543 ( .Q(n5737), .DIN1(WX891), .DIN2(CRC_OUT_9_31) );
  nor2s1 U8544 ( .Q(WX1270), .DIN1(n3394), .DIN2(n5738) );
  xor2s1 U8545 ( .Q(n5738), .DIN1(WX893), .DIN2(CRC_OUT_9_2) );
  nor2s1 U8546 ( .Q(WX1268), .DIN1(n3394), .DIN2(n5739) );
  xor2s1 U8547 ( .Q(n5739), .DIN1(WX895), .DIN2(CRC_OUT_9_1) );
  nor2s1 U8548 ( .Q(WX1266), .DIN1(n3394), .DIN2(n5740) );
  xor2s1 U8549 ( .Q(n5740), .DIN1(WX897), .DIN2(CRC_OUT_9_0) );
  nor2s1 U8550 ( .Q(WX1264), .DIN1(n3394), .DIN2(n5741) );
  xor2s1 U8551 ( .Q(n5741), .DIN1(WX899), .DIN2(CRC_OUT_9_31) );
  xor2s1 U8552 ( .Q(WX1227), .DIN1(n4341), .DIN2(n5742) );
  nnd2s1 U8553 ( .Q(n5742), .DIN1(WX547), .DIN2(TM0) );
  xor2s1 U8554 ( .Q(n4341), .DIN1(n5743), .DIN2(n5744) );
  xor2s1 U8555 ( .Q(n5744), .DIN1(n3362), .DIN2(WX707) );
  xor2s1 U8556 ( .Q(n5743), .DIN1(WX771), .DIN2(n5746) );
  xor2s1 U8557 ( .Q(n5746), .DIN1(WX899), .DIN2(WX835) );
  xor2s1 U8558 ( .Q(WX1220), .DIN1(n4348), .DIN2(n5747) );
  nnd2s1 U8559 ( .Q(n5747), .DIN1(WX545), .DIN2(TM0) );
  xor2s1 U8560 ( .Q(n4348), .DIN1(n5748), .DIN2(n5749) );
  xor2s1 U8561 ( .Q(n5749), .DIN1(n3361), .DIN2(WX705) );
  xor2s1 U8562 ( .Q(n5748), .DIN1(WX769), .DIN2(n5750) );
  xor2s1 U8563 ( .Q(n5750), .DIN1(WX897), .DIN2(WX833) );
  xor2s1 U8564 ( .Q(WX1213), .DIN1(n4355), .DIN2(n5751) );
  nnd2s1 U8565 ( .Q(n5751), .DIN1(WX543), .DIN2(TM0) );
  xor2s1 U8566 ( .Q(n4355), .DIN1(n5752), .DIN2(n5753) );
  xor2s1 U8567 ( .Q(n5753), .DIN1(n3361), .DIN2(WX703) );
  xor2s1 U8568 ( .Q(n5752), .DIN1(WX767), .DIN2(n5754) );
  xor2s1 U8569 ( .Q(n5754), .DIN1(WX895), .DIN2(WX831) );
  xor2s1 U8570 ( .Q(WX1206), .DIN1(n4362), .DIN2(n5755) );
  nnd2s1 U8571 ( .Q(n5755), .DIN1(WX541), .DIN2(TM0) );
  xor2s1 U8572 ( .Q(n4362), .DIN1(n5756), .DIN2(n5757) );
  xor2s1 U8573 ( .Q(n5757), .DIN1(n3361), .DIN2(WX701) );
  xor2s1 U8574 ( .Q(n5756), .DIN1(WX765), .DIN2(n5758) );
  xor2s1 U8575 ( .Q(n5758), .DIN1(WX893), .DIN2(WX829) );
  xor2s1 U8576 ( .Q(WX1199), .DIN1(n4369), .DIN2(n5759) );
  nnd2s1 U8577 ( .Q(n5759), .DIN1(WX539), .DIN2(TM0) );
  xor2s1 U8578 ( .Q(n4369), .DIN1(n5760), .DIN2(n5761) );
  xor2s1 U8579 ( .Q(n5761), .DIN1(n5745), .DIN2(WX699) );
  xor2s1 U8580 ( .Q(n5760), .DIN1(WX763), .DIN2(n5762) );
  xor2s1 U8581 ( .Q(n5762), .DIN1(WX891), .DIN2(WX827) );
  xor2s1 U8582 ( .Q(WX1192), .DIN1(n4376), .DIN2(n5763) );
  nnd2s1 U8583 ( .Q(n5763), .DIN1(WX537), .DIN2(TM0) );
  xor2s1 U8584 ( .Q(n4376), .DIN1(n5764), .DIN2(n5765) );
  xor2s1 U8585 ( .Q(n5765), .DIN1(n5745), .DIN2(WX697) );
  xor2s1 U8586 ( .Q(n5764), .DIN1(WX761), .DIN2(n5766) );
  xor2s1 U8587 ( .Q(n5766), .DIN1(WX889), .DIN2(WX825) );
  xor2s1 U8588 ( .Q(WX1185), .DIN1(n4383), .DIN2(n5767) );
  nnd2s1 U8589 ( .Q(n5767), .DIN1(WX535), .DIN2(TM0) );
  xor2s1 U8590 ( .Q(n4383), .DIN1(n5768), .DIN2(n5769) );
  xor2s1 U8591 ( .Q(n5769), .DIN1(n3361), .DIN2(WX695) );
  xor2s1 U8592 ( .Q(n5768), .DIN1(WX759), .DIN2(n5770) );
  xor2s1 U8593 ( .Q(n5770), .DIN1(WX887), .DIN2(WX823) );
  xor2s1 U8594 ( .Q(WX1178), .DIN1(n4390), .DIN2(n5771) );
  nnd2s1 U8595 ( .Q(n5771), .DIN1(WX533), .DIN2(TM0) );
  xor2s1 U8596 ( .Q(n4390), .DIN1(n5772), .DIN2(n5773) );
  xor2s1 U8597 ( .Q(n5773), .DIN1(n3362), .DIN2(WX693) );
  xor2s1 U8598 ( .Q(n5772), .DIN1(WX757), .DIN2(n5774) );
  xor2s1 U8599 ( .Q(n5774), .DIN1(WX885), .DIN2(WX821) );
  xor2s1 U8600 ( .Q(WX1171), .DIN1(n4397), .DIN2(n5775) );
  nnd2s1 U8601 ( .Q(n5775), .DIN1(WX531), .DIN2(TM0) );
  xor2s1 U8602 ( .Q(n4397), .DIN1(n5776), .DIN2(n5777) );
  xor2s1 U8603 ( .Q(n5777), .DIN1(n3362), .DIN2(WX691) );
  xor2s1 U8604 ( .Q(n5776), .DIN1(WX755), .DIN2(n5778) );
  xor2s1 U8605 ( .Q(n5778), .DIN1(WX883), .DIN2(WX819) );
  nor2s1 U8606 ( .Q(WX11670), .DIN1(n3395), .DIN2(n5779) );
  xor2s1 U8607 ( .Q(n5779), .DIN1(WX11181), .DIN2(CRC_OUT_1_30) );
  nor2s1 U8608 ( .Q(WX11668), .DIN1(n3395), .DIN2(n5780) );
  xor2s1 U8609 ( .Q(n5780), .DIN1(WX11183), .DIN2(CRC_OUT_1_29) );
  nor2s1 U8610 ( .Q(WX11666), .DIN1(n3395), .DIN2(n5781) );
  xor2s1 U8611 ( .Q(n5781), .DIN1(WX11185), .DIN2(CRC_OUT_1_28) );
  nor2s1 U8612 ( .Q(WX11664), .DIN1(n3395), .DIN2(n5782) );
  xor2s1 U8613 ( .Q(n5782), .DIN1(WX11187), .DIN2(CRC_OUT_1_27) );
  nor2s1 U8614 ( .Q(WX11662), .DIN1(n3395), .DIN2(n5783) );
  xor2s1 U8615 ( .Q(n5783), .DIN1(WX11189), .DIN2(CRC_OUT_1_26) );
  nor2s1 U8616 ( .Q(WX11660), .DIN1(n3395), .DIN2(n5784) );
  xor2s1 U8617 ( .Q(n5784), .DIN1(WX11191), .DIN2(CRC_OUT_1_25) );
  nor2s1 U8618 ( .Q(WX11658), .DIN1(n3395), .DIN2(n5785) );
  xor2s1 U8619 ( .Q(n5785), .DIN1(WX11193), .DIN2(CRC_OUT_1_24) );
  nor2s1 U8620 ( .Q(WX11656), .DIN1(n3395), .DIN2(n5786) );
  xor2s1 U8621 ( .Q(n5786), .DIN1(WX11195), .DIN2(CRC_OUT_1_23) );
  nor2s1 U8622 ( .Q(WX11654), .DIN1(n3395), .DIN2(n5787) );
  xor2s1 U8623 ( .Q(n5787), .DIN1(WX11197), .DIN2(CRC_OUT_1_22) );
  nor2s1 U8624 ( .Q(WX11652), .DIN1(n3395), .DIN2(n5788) );
  xor2s1 U8625 ( .Q(n5788), .DIN1(WX11199), .DIN2(CRC_OUT_1_21) );
  nor2s1 U8626 ( .Q(WX11650), .DIN1(n3396), .DIN2(n5789) );
  xor2s1 U8627 ( .Q(n5789), .DIN1(WX11201), .DIN2(CRC_OUT_1_20) );
  nor2s1 U8628 ( .Q(WX11648), .DIN1(n3396), .DIN2(n5790) );
  xor2s1 U8629 ( .Q(n5790), .DIN1(WX11203), .DIN2(CRC_OUT_1_19) );
  nor2s1 U8630 ( .Q(WX11646), .DIN1(n3396), .DIN2(n5791) );
  xor2s1 U8631 ( .Q(n5791), .DIN1(WX11205), .DIN2(CRC_OUT_1_18) );
  nor2s1 U8632 ( .Q(WX11644), .DIN1(n3396), .DIN2(n5792) );
  xor2s1 U8633 ( .Q(n5792), .DIN1(WX11207), .DIN2(CRC_OUT_1_17) );
  nor2s1 U8634 ( .Q(WX11642), .DIN1(n3396), .DIN2(n5793) );
  xor2s1 U8635 ( .Q(n5793), .DIN1(WX11209), .DIN2(CRC_OUT_1_16) );
  nor2s1 U8636 ( .Q(WX11640), .DIN1(n3396), .DIN2(n5794) );
  xor2s1 U8637 ( .Q(n5794), .DIN1(CRC_OUT_1_15), .DIN2(n5795) );
  xor2s1 U8638 ( .Q(n5795), .DIN1(WX11211), .DIN2(CRC_OUT_1_31) );
  xor2s1 U8639 ( .Q(WX1164), .DIN1(n4404), .DIN2(n5796) );
  nnd2s1 U8640 ( .Q(n5796), .DIN1(WX529), .DIN2(TM0) );
  xor2s1 U8641 ( .Q(n4404), .DIN1(n5797), .DIN2(n5798) );
  xor2s1 U8642 ( .Q(n5798), .DIN1(n3361), .DIN2(WX689) );
  xor2s1 U8643 ( .Q(n5797), .DIN1(WX753), .DIN2(n5799) );
  xor2s1 U8644 ( .Q(n5799), .DIN1(WX881), .DIN2(WX817) );
  nor2s1 U8645 ( .Q(WX11638), .DIN1(n3396), .DIN2(n5800) );
  xor2s1 U8646 ( .Q(n5800), .DIN1(WX11213), .DIN2(CRC_OUT_1_14) );
  nor2s1 U8647 ( .Q(WX11636), .DIN1(n3396), .DIN2(n5801) );
  xor2s1 U8648 ( .Q(n5801), .DIN1(WX11215), .DIN2(CRC_OUT_1_13) );
  nor2s1 U8649 ( .Q(WX11634), .DIN1(n3396), .DIN2(n5802) );
  xor2s1 U8650 ( .Q(n5802), .DIN1(WX11217), .DIN2(CRC_OUT_1_12) );
  nor2s1 U8651 ( .Q(WX11632), .DIN1(n3396), .DIN2(n5803) );
  xor2s1 U8652 ( .Q(n5803), .DIN1(WX11219), .DIN2(CRC_OUT_1_11) );
  nor2s1 U8653 ( .Q(WX11630), .DIN1(n3397), .DIN2(n5804) );
  xor2s1 U8654 ( .Q(n5804), .DIN1(CRC_OUT_1_10), .DIN2(n5805) );
  xor2s1 U8655 ( .Q(n5805), .DIN1(WX11221), .DIN2(CRC_OUT_1_31) );
  nor2s1 U8656 ( .Q(WX11628), .DIN1(n3397), .DIN2(n5806) );
  xor2s1 U8657 ( .Q(n5806), .DIN1(WX11223), .DIN2(CRC_OUT_1_9) );
  nor2s1 U8658 ( .Q(WX11626), .DIN1(n3397), .DIN2(n5807) );
  xor2s1 U8659 ( .Q(n5807), .DIN1(WX11225), .DIN2(CRC_OUT_1_8) );
  nor2s1 U8660 ( .Q(WX11624), .DIN1(n3397), .DIN2(n5808) );
  xor2s1 U8661 ( .Q(n5808), .DIN1(WX11227), .DIN2(CRC_OUT_1_7) );
  nor2s1 U8662 ( .Q(WX11622), .DIN1(n3397), .DIN2(n5809) );
  xor2s1 U8663 ( .Q(n5809), .DIN1(WX11229), .DIN2(CRC_OUT_1_6) );
  nor2s1 U8664 ( .Q(WX11620), .DIN1(n3397), .DIN2(n5810) );
  xor2s1 U8665 ( .Q(n5810), .DIN1(WX11231), .DIN2(CRC_OUT_1_5) );
  nor2s1 U8666 ( .Q(WX11618), .DIN1(n3397), .DIN2(n5811) );
  xor2s1 U8667 ( .Q(n5811), .DIN1(WX11233), .DIN2(CRC_OUT_1_4) );
  nor2s1 U8668 ( .Q(WX11616), .DIN1(n3397), .DIN2(n5812) );
  xor2s1 U8669 ( .Q(n5812), .DIN1(CRC_OUT_1_3), .DIN2(n5813) );
  xor2s1 U8670 ( .Q(n5813), .DIN1(WX11235), .DIN2(CRC_OUT_1_31) );
  nor2s1 U8671 ( .Q(WX11614), .DIN1(n3397), .DIN2(n5814) );
  xor2s1 U8672 ( .Q(n5814), .DIN1(WX11237), .DIN2(CRC_OUT_1_2) );
  nor2s1 U8673 ( .Q(WX11612), .DIN1(n3398), .DIN2(n5815) );
  xor2s1 U8674 ( .Q(n5815), .DIN1(WX11239), .DIN2(CRC_OUT_1_1) );
  nor2s1 U8675 ( .Q(WX11610), .DIN1(n3398), .DIN2(n5816) );
  xor2s1 U8676 ( .Q(n5816), .DIN1(WX11241), .DIN2(CRC_OUT_1_0) );
  nor2s1 U8677 ( .Q(WX11608), .DIN1(n3398), .DIN2(n5817) );
  xor2s1 U8678 ( .Q(n5817), .DIN1(WX11243), .DIN2(CRC_OUT_1_31) );
  xor2s1 U8679 ( .Q(WX1157), .DIN1(n4411), .DIN2(n5818) );
  nnd2s1 U8680 ( .Q(n5818), .DIN1(WX527), .DIN2(TM0) );
  xor2s1 U8681 ( .Q(n4411), .DIN1(n5819), .DIN2(n5820) );
  xor2s1 U8682 ( .Q(n5820), .DIN1(n5745), .DIN2(WX687) );
  xor2s1 U8683 ( .Q(n5819), .DIN1(WX751), .DIN2(n5821) );
  xor2s1 U8684 ( .Q(n5821), .DIN1(WX879), .DIN2(WX815) );
  xor2s1 U8685 ( .Q(WX1150), .DIN1(n4418), .DIN2(n5822) );
  nnd2s1 U8686 ( .Q(n5822), .DIN1(WX525), .DIN2(TM0) );
  xor2s1 U8687 ( .Q(n4418), .DIN1(n5823), .DIN2(n5824) );
  xor2s1 U8688 ( .Q(n5824), .DIN1(n3362), .DIN2(WX685) );
  xor2s1 U8689 ( .Q(n5823), .DIN1(WX749), .DIN2(n5825) );
  xor2s1 U8690 ( .Q(n5825), .DIN1(WX877), .DIN2(WX813) );
  xor2s1 U8691 ( .Q(WX1143), .DIN1(n4425), .DIN2(n5826) );
  nnd2s1 U8692 ( .Q(n5826), .DIN1(WX523), .DIN2(TM0) );
  xor2s1 U8693 ( .Q(n4425), .DIN1(n5827), .DIN2(n5828) );
  xor2s1 U8694 ( .Q(n5828), .DIN1(n5745), .DIN2(WX683) );
  xor2s1 U8695 ( .Q(n5827), .DIN1(WX747), .DIN2(n5829) );
  xor2s1 U8696 ( .Q(n5829), .DIN1(WX875), .DIN2(WX811) );
  xor2s1 U8697 ( .Q(WX1136), .DIN1(n4432), .DIN2(n5830) );
  nnd2s1 U8698 ( .Q(n5830), .DIN1(WX521), .DIN2(TM0) );
  xor2s1 U8699 ( .Q(n4432), .DIN1(n5831), .DIN2(n5832) );
  xor2s1 U8700 ( .Q(n5832), .DIN1(n3361), .DIN2(WX681) );
  xor2s1 U8701 ( .Q(n5831), .DIN1(WX745), .DIN2(n5833) );
  xor2s1 U8702 ( .Q(n5833), .DIN1(WX873), .DIN2(WX809) );
  xor2s1 U8703 ( .Q(WX1129), .DIN1(n4439), .DIN2(n5834) );
  nnd2s1 U8704 ( .Q(n5834), .DIN1(WX519), .DIN2(TM0) );
  xor2s1 U8705 ( .Q(n4439), .DIN1(n5835), .DIN2(n5836) );
  xor2s1 U8706 ( .Q(n5836), .DIN1(n3362), .DIN2(WX679) );
  xor2s1 U8707 ( .Q(n5835), .DIN1(WX743), .DIN2(n5837) );
  xor2s1 U8708 ( .Q(n5837), .DIN1(WX871), .DIN2(WX807) );
  and2s1 U8709 ( .Q(WX11242), .DIN1(RESET), .DIN2(WX11179) );
  and2s1 U8710 ( .Q(WX11240), .DIN1(RESET), .DIN2(WX11177) );
  and2s1 U8711 ( .Q(WX11238), .DIN1(RESET), .DIN2(WX11175) );
  and2s1 U8712 ( .Q(WX11236), .DIN1(RESET), .DIN2(WX11173) );
  and2s1 U8713 ( .Q(WX11234), .DIN1(RESET), .DIN2(WX11171) );
  and2s1 U8714 ( .Q(WX11232), .DIN1(RESET), .DIN2(WX11169) );
  and2s1 U8715 ( .Q(WX11230), .DIN1(RESET), .DIN2(WX11167) );
  and2s1 U8716 ( .Q(WX11228), .DIN1(RESET), .DIN2(WX11165) );
  and2s1 U8717 ( .Q(WX11226), .DIN1(RESET), .DIN2(WX11163) );
  and2s1 U8718 ( .Q(WX11224), .DIN1(RESET), .DIN2(WX11161) );
  and2s1 U8719 ( .Q(WX11222), .DIN1(RESET), .DIN2(WX11159) );
  and2s1 U8720 ( .Q(WX11220), .DIN1(RESET), .DIN2(WX11157) );
  xor2s1 U8721 ( .Q(WX1122), .DIN1(n4446), .DIN2(n5838) );
  nnd2s1 U8722 ( .Q(n5838), .DIN1(WX517), .DIN2(TM0) );
  xor2s1 U8723 ( .Q(n4446), .DIN1(n5839), .DIN2(n5840) );
  xor2s1 U8724 ( .Q(n5840), .DIN1(n5745), .DIN2(WX677) );
  xor2s1 U8725 ( .Q(n5839), .DIN1(WX741), .DIN2(n5841) );
  xor2s1 U8726 ( .Q(n5841), .DIN1(WX869), .DIN2(WX805) );
  and2s1 U8727 ( .Q(WX11218), .DIN1(RESET), .DIN2(WX11155) );
  and2s1 U8728 ( .Q(WX11216), .DIN1(RESET), .DIN2(WX11153) );
  and2s1 U8729 ( .Q(WX11214), .DIN1(RESET), .DIN2(WX11151) );
  and2s1 U8730 ( .Q(WX11212), .DIN1(RESET), .DIN2(WX11149) );
  and2s1 U8731 ( .Q(WX11210), .DIN1(RESET), .DIN2(WX11147) );
  and2s1 U8732 ( .Q(WX11208), .DIN1(RESET), .DIN2(WX11145) );
  and2s1 U8733 ( .Q(WX11206), .DIN1(RESET), .DIN2(WX11143) );
  and2s1 U8734 ( .Q(WX11204), .DIN1(RESET), .DIN2(WX11141) );
  and2s1 U8735 ( .Q(WX11202), .DIN1(RESET), .DIN2(WX11139) );
  and2s1 U8736 ( .Q(WX11200), .DIN1(RESET), .DIN2(WX11137) );
  and2s1 U8737 ( .Q(WX11198), .DIN1(RESET), .DIN2(WX11135) );
  and2s1 U8738 ( .Q(WX11196), .DIN1(RESET), .DIN2(WX11133) );
  and2s1 U8739 ( .Q(WX11194), .DIN1(RESET), .DIN2(WX11131) );
  and2s1 U8740 ( .Q(WX11192), .DIN1(RESET), .DIN2(WX11129) );
  and2s1 U8741 ( .Q(WX11190), .DIN1(RESET), .DIN2(WX11127) );
  and2s1 U8742 ( .Q(WX11188), .DIN1(RESET), .DIN2(WX11125) );
  and2s1 U8743 ( .Q(WX11186), .DIN1(RESET), .DIN2(WX11123) );
  and2s1 U8744 ( .Q(WX11184), .DIN1(RESET), .DIN2(WX11121) );
  and2s1 U8745 ( .Q(WX11182), .DIN1(RESET), .DIN2(WX11119) );
  and2s1 U8746 ( .Q(WX11180), .DIN1(RESET), .DIN2(WX11117) );
  nor2s1 U8747 ( .Q(WX11178), .DIN1(n3398), .DIN2(n3077) );
  nor2s1 U8748 ( .Q(WX11176), .DIN1(n3398), .DIN2(n3078) );
  nor2s1 U8749 ( .Q(WX11174), .DIN1(n3398), .DIN2(n3079) );
  nor2s1 U8750 ( .Q(WX11172), .DIN1(n3398), .DIN2(n3080) );
  nor2s1 U8751 ( .Q(WX11170), .DIN1(n3398), .DIN2(n3081) );
  nor2s1 U8752 ( .Q(WX11168), .DIN1(n3398), .DIN2(n3082) );
  nor2s1 U8753 ( .Q(WX11166), .DIN1(n3398), .DIN2(n3083) );
  nor2s1 U8754 ( .Q(WX11164), .DIN1(n3399), .DIN2(n3084) );
  nor2s1 U8755 ( .Q(WX11162), .DIN1(n3399), .DIN2(n3085) );
  nor2s1 U8756 ( .Q(WX11160), .DIN1(n3399), .DIN2(n3086) );
  nor2s1 U8757 ( .Q(WX11158), .DIN1(n3399), .DIN2(n3087) );
  nor2s1 U8758 ( .Q(WX11156), .DIN1(n3399), .DIN2(n3088) );
  nor2s1 U8759 ( .Q(WX11154), .DIN1(n3399), .DIN2(n3089) );
  nor2s1 U8760 ( .Q(WX11152), .DIN1(n3399), .DIN2(n3090) );
  nor2s1 U8761 ( .Q(WX11150), .DIN1(n3399), .DIN2(n3091) );
  xor2s1 U8762 ( .Q(WX1115), .DIN1(n4453), .DIN2(n5842) );
  nnd2s1 U8763 ( .Q(n5842), .DIN1(WX515), .DIN2(TM0) );
  xor2s1 U8764 ( .Q(n4453), .DIN1(n5843), .DIN2(n5844) );
  xor2s1 U8765 ( .Q(n5844), .DIN1(n3575), .DIN2(WX675) );
  xor2s1 U8766 ( .Q(n5843), .DIN1(WX739), .DIN2(n5845) );
  xor2s1 U8767 ( .Q(n5845), .DIN1(WX867), .DIN2(WX803) );
  nor2s1 U8768 ( .Q(WX11148), .DIN1(n3399), .DIN2(n3092) );
  nor2s1 U8769 ( .Q(WX11146), .DIN1(n3399), .DIN2(n3093) );
  nor2s1 U8770 ( .Q(WX11144), .DIN1(n3400), .DIN2(n3094) );
  nor2s1 U8771 ( .Q(WX11142), .DIN1(n3400), .DIN2(n3095) );
  nor2s1 U8772 ( .Q(WX11140), .DIN1(n3400), .DIN2(n3096) );
  nor2s1 U8773 ( .Q(WX11138), .DIN1(n3400), .DIN2(n3097) );
  nor2s1 U8774 ( .Q(WX11136), .DIN1(n3400), .DIN2(n3098) );
  nor2s1 U8775 ( .Q(WX11134), .DIN1(n3400), .DIN2(n3099) );
  nor2s1 U8776 ( .Q(WX11132), .DIN1(n3400), .DIN2(n3100) );
  nor2s1 U8777 ( .Q(WX11130), .DIN1(n3400), .DIN2(n3101) );
  nor2s1 U8778 ( .Q(WX11128), .DIN1(n3400), .DIN2(n3102) );
  nor2s1 U8779 ( .Q(WX11126), .DIN1(n3400), .DIN2(n3103) );
  nor2s1 U8780 ( .Q(WX11124), .DIN1(n3401), .DIN2(n3104) );
  nor2s1 U8781 ( .Q(WX11122), .DIN1(n3401), .DIN2(n3105) );
  nor2s1 U8782 ( .Q(WX11120), .DIN1(n3401), .DIN2(n3106) );
  nor2s1 U8783 ( .Q(WX11118), .DIN1(n3401), .DIN2(n3107) );
  nor2s1 U8784 ( .Q(WX11116), .DIN1(n3401), .DIN2(n3108) );
  and2s1 U8785 ( .Q(WX11114), .DIN1(RESET), .DIN2(WX11051) );
  and2s1 U8786 ( .Q(WX11112), .DIN1(RESET), .DIN2(WX11049) );
  and2s1 U8787 ( .Q(WX11110), .DIN1(RESET), .DIN2(WX11047) );
  and2s1 U8788 ( .Q(WX11108), .DIN1(RESET), .DIN2(WX11045) );
  and2s1 U8789 ( .Q(WX11106), .DIN1(RESET), .DIN2(WX11043) );
  and2s1 U8790 ( .Q(WX11104), .DIN1(RESET), .DIN2(WX11041) );
  and2s1 U8791 ( .Q(WX11102), .DIN1(RESET), .DIN2(WX11039) );
  and2s1 U8792 ( .Q(WX11100), .DIN1(RESET), .DIN2(WX11037) );
  and2s1 U8793 ( .Q(WX11098), .DIN1(RESET), .DIN2(WX11035) );
  and2s1 U8794 ( .Q(WX11096), .DIN1(RESET), .DIN2(WX11033) );
  and2s1 U8795 ( .Q(WX11094), .DIN1(RESET), .DIN2(WX11031) );
  and2s1 U8796 ( .Q(WX11092), .DIN1(RESET), .DIN2(WX11029) );
  and2s1 U8797 ( .Q(WX11090), .DIN1(RESET), .DIN2(WX11027) );
  and2s1 U8798 ( .Q(WX11088), .DIN1(RESET), .DIN2(WX11025) );
  and2s1 U8799 ( .Q(WX11086), .DIN1(RESET), .DIN2(WX11023) );
  and2s1 U8800 ( .Q(WX11084), .DIN1(RESET), .DIN2(WX11021) );
  and2s1 U8801 ( .Q(WX11082), .DIN1(RESET), .DIN2(WX11019) );
  and2s1 U8802 ( .Q(WX11080), .DIN1(RESET), .DIN2(WX11017) );
  xor2s1 U8803 ( .Q(WX1108), .DIN1(n4460), .DIN2(n5846) );
  nnd2s1 U8804 ( .Q(n5846), .DIN1(WX513), .DIN2(TM0) );
  xor2s1 U8805 ( .Q(n4460), .DIN1(n5847), .DIN2(n5848) );
  xor2s1 U8806 ( .Q(n5848), .DIN1(n3575), .DIN2(WX673) );
  xor2s1 U8807 ( .Q(n5847), .DIN1(WX737), .DIN2(n5849) );
  xor2s1 U8808 ( .Q(n5849), .DIN1(WX865), .DIN2(WX801) );
  and2s1 U8809 ( .Q(WX11078), .DIN1(RESET), .DIN2(WX11015) );
  and2s1 U8810 ( .Q(WX11076), .DIN1(RESET), .DIN2(WX11013) );
  and2s1 U8811 ( .Q(WX11074), .DIN1(RESET), .DIN2(WX11011) );
  and2s1 U8812 ( .Q(WX11072), .DIN1(RESET), .DIN2(WX11009) );
  and2s1 U8813 ( .Q(WX11070), .DIN1(RESET), .DIN2(WX11007) );
  and2s1 U8814 ( .Q(WX11068), .DIN1(RESET), .DIN2(WX11005) );
  and2s1 U8815 ( .Q(WX11066), .DIN1(RESET), .DIN2(WX11003) );
  and2s1 U8816 ( .Q(WX11064), .DIN1(RESET), .DIN2(WX11001) );
  and2s1 U8817 ( .Q(WX11062), .DIN1(RESET), .DIN2(WX10999) );
  and2s1 U8818 ( .Q(WX11060), .DIN1(RESET), .DIN2(WX10997) );
  and2s1 U8819 ( .Q(WX11058), .DIN1(RESET), .DIN2(WX10995) );
  and2s1 U8820 ( .Q(WX11056), .DIN1(RESET), .DIN2(WX10993) );
  and2s1 U8821 ( .Q(WX11054), .DIN1(RESET), .DIN2(WX10991) );
  and2s1 U8822 ( .Q(WX11052), .DIN1(RESET), .DIN2(WX10989) );
  nnd4s1 U8823 ( .Q(WX11050), .DIN1(n5850), .DIN2(n5851), .DIN3(n5852), .DIN4(
        n5853) );
  nnd2s1 U8824 ( .Q(n5853), .DIN1(n3435), .DIN2(n3595) );
  xor2s1 U8825 ( .Q(n3595), .DIN1(n5854), .DIN2(n5855) );
  xor2s1 U8826 ( .Q(n5855), .DIN1(n3077), .DIN2(WX11051) );
  xor2s1 U8827 ( .Q(n5854), .DIN1(n3317), .DIN2(WX11179) );
  nnd2s1 U8828 ( .Q(n5852), .DIN1(WX10891), .DIN2(n3497) );
  nnd2s1 U8829 ( .Q(n5851), .DIN1(DATA_0_0), .DIN2(n3483) );
  nnd2s1 U8830 ( .Q(n5850), .DIN1(CRC_OUT_1_0), .DIN2(n3529) );
  nnd4s1 U8831 ( .Q(WX11048), .DIN1(n5856), .DIN2(n5857), .DIN3(n5858), .DIN4(
        n5859) );
  nnd2s1 U8832 ( .Q(n5859), .DIN1(n3435), .DIN2(n3603) );
  xor2s1 U8833 ( .Q(n3603), .DIN1(n5860), .DIN2(n5861) );
  xor2s1 U8834 ( .Q(n5861), .DIN1(n3078), .DIN2(WX11049) );
  xor2s1 U8835 ( .Q(n5860), .DIN1(n3318), .DIN2(WX11177) );
  nnd2s1 U8836 ( .Q(n5858), .DIN1(WX10889), .DIN2(n3497) );
  nnd2s1 U8837 ( .Q(n5857), .DIN1(DATA_0_1), .DIN2(n3483) );
  nnd2s1 U8838 ( .Q(n5856), .DIN1(CRC_OUT_1_1), .DIN2(n3529) );
  nnd4s1 U8839 ( .Q(WX11046), .DIN1(n5862), .DIN2(n5863), .DIN3(n5864), .DIN4(
        n5865) );
  nnd2s1 U8840 ( .Q(n5865), .DIN1(n3435), .DIN2(n3609) );
  xor2s1 U8841 ( .Q(n3609), .DIN1(n5866), .DIN2(n5867) );
  xor2s1 U8842 ( .Q(n5867), .DIN1(n3079), .DIN2(WX11047) );
  xor2s1 U8843 ( .Q(n5866), .DIN1(n3319), .DIN2(WX11175) );
  nnd2s1 U8844 ( .Q(n5864), .DIN1(WX10887), .DIN2(n3497) );
  nnd2s1 U8845 ( .Q(n5863), .DIN1(DATA_0_2), .DIN2(n3483) );
  nnd2s1 U8846 ( .Q(n5862), .DIN1(CRC_OUT_1_2), .DIN2(n3529) );
  nnd4s1 U8847 ( .Q(WX11044), .DIN1(n5868), .DIN2(n5869), .DIN3(n5870), .DIN4(
        n5871) );
  nnd2s1 U8848 ( .Q(n5871), .DIN1(n3435), .DIN2(n3615) );
  xor2s1 U8849 ( .Q(n3615), .DIN1(n5872), .DIN2(n5873) );
  xor2s1 U8850 ( .Q(n5873), .DIN1(n3080), .DIN2(WX11045) );
  xor2s1 U8851 ( .Q(n5872), .DIN1(n3320), .DIN2(WX11173) );
  nnd2s1 U8852 ( .Q(n5870), .DIN1(WX10885), .DIN2(n3497) );
  nnd2s1 U8853 ( .Q(n5869), .DIN1(DATA_0_3), .DIN2(n3483) );
  nnd2s1 U8854 ( .Q(n5868), .DIN1(CRC_OUT_1_3), .DIN2(n3529) );
  nnd4s1 U8855 ( .Q(WX11042), .DIN1(n5874), .DIN2(n5875), .DIN3(n5876), .DIN4(
        n5877) );
  nnd2s1 U8856 ( .Q(n5877), .DIN1(n3435), .DIN2(n3621) );
  xor2s1 U8857 ( .Q(n3621), .DIN1(n5878), .DIN2(n5879) );
  xor2s1 U8858 ( .Q(n5879), .DIN1(n3081), .DIN2(WX11043) );
  xor2s1 U8859 ( .Q(n5878), .DIN1(n3321), .DIN2(WX11171) );
  nnd2s1 U8860 ( .Q(n5876), .DIN1(WX10883), .DIN2(n3497) );
  nnd2s1 U8861 ( .Q(n5875), .DIN1(DATA_0_4), .DIN2(n3484) );
  nnd2s1 U8862 ( .Q(n5874), .DIN1(CRC_OUT_1_4), .DIN2(n3529) );
  nnd4s1 U8863 ( .Q(WX11040), .DIN1(n5880), .DIN2(n5881), .DIN3(n5882), .DIN4(
        n5883) );
  nnd2s1 U8864 ( .Q(n5883), .DIN1(n3435), .DIN2(n3627) );
  xor2s1 U8865 ( .Q(n3627), .DIN1(n5884), .DIN2(n5885) );
  xor2s1 U8866 ( .Q(n5885), .DIN1(n3082), .DIN2(WX11041) );
  xor2s1 U8867 ( .Q(n5884), .DIN1(n3322), .DIN2(WX11169) );
  nnd2s1 U8868 ( .Q(n5882), .DIN1(WX10881), .DIN2(n3497) );
  nnd2s1 U8869 ( .Q(n5881), .DIN1(DATA_0_5), .DIN2(n3484) );
  nnd2s1 U8870 ( .Q(n5880), .DIN1(CRC_OUT_1_5), .DIN2(n3529) );
  nnd4s1 U8871 ( .Q(WX11038), .DIN1(n5886), .DIN2(n5887), .DIN3(n5888), .DIN4(
        n5889) );
  nnd2s1 U8872 ( .Q(n5889), .DIN1(n3434), .DIN2(n3633) );
  xor2s1 U8873 ( .Q(n3633), .DIN1(n5890), .DIN2(n5891) );
  xor2s1 U8874 ( .Q(n5891), .DIN1(n3083), .DIN2(WX11039) );
  xor2s1 U8875 ( .Q(n5890), .DIN1(n3323), .DIN2(WX11167) );
  nnd2s1 U8876 ( .Q(n5888), .DIN1(WX10879), .DIN2(n3497) );
  nnd2s1 U8877 ( .Q(n5887), .DIN1(DATA_0_6), .DIN2(n3484) );
  nnd2s1 U8878 ( .Q(n5886), .DIN1(CRC_OUT_1_6), .DIN2(n3529) );
  nnd4s1 U8879 ( .Q(WX11036), .DIN1(n5892), .DIN2(n5893), .DIN3(n5894), .DIN4(
        n5895) );
  nnd2s1 U8880 ( .Q(n5895), .DIN1(n3434), .DIN2(n3639) );
  xor2s1 U8881 ( .Q(n3639), .DIN1(n5896), .DIN2(n5897) );
  xor2s1 U8882 ( .Q(n5897), .DIN1(n3084), .DIN2(WX11037) );
  xor2s1 U8883 ( .Q(n5896), .DIN1(n3324), .DIN2(WX11165) );
  nnd2s1 U8884 ( .Q(n5894), .DIN1(WX10877), .DIN2(n3497) );
  nnd2s1 U8885 ( .Q(n5893), .DIN1(DATA_0_7), .DIN2(n3484) );
  nnd2s1 U8886 ( .Q(n5892), .DIN1(CRC_OUT_1_7), .DIN2(n3529) );
  nnd4s1 U8887 ( .Q(WX11034), .DIN1(n5898), .DIN2(n5899), .DIN3(n5900), .DIN4(
        n5901) );
  nnd2s1 U8888 ( .Q(n5901), .DIN1(n3434), .DIN2(n3645) );
  xor2s1 U8889 ( .Q(n3645), .DIN1(n5902), .DIN2(n5903) );
  xor2s1 U8890 ( .Q(n5903), .DIN1(n3085), .DIN2(WX11035) );
  xor2s1 U8891 ( .Q(n5902), .DIN1(n3325), .DIN2(WX11163) );
  nnd2s1 U8892 ( .Q(n5900), .DIN1(WX10875), .DIN2(n3496) );
  nnd2s1 U8893 ( .Q(n5899), .DIN1(DATA_0_8), .DIN2(n3484) );
  nnd2s1 U8894 ( .Q(n5898), .DIN1(CRC_OUT_1_8), .DIN2(n3528) );
  nnd4s1 U8895 ( .Q(WX11032), .DIN1(n5904), .DIN2(n5905), .DIN3(n5906), .DIN4(
        n5907) );
  nnd2s1 U8896 ( .Q(n5907), .DIN1(n3434), .DIN2(n3651) );
  xor2s1 U8897 ( .Q(n3651), .DIN1(n5908), .DIN2(n5909) );
  xor2s1 U8898 ( .Q(n5909), .DIN1(n3086), .DIN2(WX11033) );
  xor2s1 U8899 ( .Q(n5908), .DIN1(n3326), .DIN2(WX11161) );
  nnd2s1 U8900 ( .Q(n5906), .DIN1(WX10873), .DIN2(n3496) );
  nnd2s1 U8901 ( .Q(n5905), .DIN1(DATA_0_9), .DIN2(n3484) );
  nnd2s1 U8902 ( .Q(n5904), .DIN1(CRC_OUT_1_9), .DIN2(n3528) );
  nnd4s1 U8903 ( .Q(WX11030), .DIN1(n5910), .DIN2(n5911), .DIN3(n5912), .DIN4(
        n5913) );
  nnd2s1 U8904 ( .Q(n5913), .DIN1(n3434), .DIN2(n3657) );
  xor2s1 U8905 ( .Q(n3657), .DIN1(n5914), .DIN2(n5915) );
  xor2s1 U8906 ( .Q(n5915), .DIN1(n3087), .DIN2(WX11031) );
  xor2s1 U8907 ( .Q(n5914), .DIN1(n3327), .DIN2(WX11159) );
  nnd2s1 U8908 ( .Q(n5912), .DIN1(WX10871), .DIN2(n3496) );
  nnd2s1 U8909 ( .Q(n5911), .DIN1(DATA_0_10), .DIN2(n3484) );
  nnd2s1 U8910 ( .Q(n5910), .DIN1(CRC_OUT_1_10), .DIN2(n3528) );
  nnd4s1 U8911 ( .Q(WX11028), .DIN1(n5916), .DIN2(n5917), .DIN3(n5918), .DIN4(
        n5919) );
  nnd2s1 U8912 ( .Q(n5919), .DIN1(n3434), .DIN2(n3663) );
  xor2s1 U8913 ( .Q(n3663), .DIN1(n5920), .DIN2(n5921) );
  xor2s1 U8914 ( .Q(n5921), .DIN1(n3088), .DIN2(WX11029) );
  xor2s1 U8915 ( .Q(n5920), .DIN1(n3328), .DIN2(WX11157) );
  nnd2s1 U8916 ( .Q(n5918), .DIN1(WX10869), .DIN2(n3496) );
  nnd2s1 U8917 ( .Q(n5917), .DIN1(DATA_0_11), .DIN2(n3484) );
  nnd2s1 U8918 ( .Q(n5916), .DIN1(CRC_OUT_1_11), .DIN2(n3528) );
  nnd4s1 U8919 ( .Q(WX11026), .DIN1(n5922), .DIN2(n5923), .DIN3(n5924), .DIN4(
        n5925) );
  nnd2s1 U8920 ( .Q(n5925), .DIN1(n3434), .DIN2(n3669) );
  xor2s1 U8921 ( .Q(n3669), .DIN1(n5926), .DIN2(n5927) );
  xor2s1 U8922 ( .Q(n5927), .DIN1(n3089), .DIN2(WX11027) );
  xor2s1 U8923 ( .Q(n5926), .DIN1(n3329), .DIN2(WX11155) );
  nnd2s1 U8924 ( .Q(n5924), .DIN1(WX10867), .DIN2(n3496) );
  nnd2s1 U8925 ( .Q(n5923), .DIN1(DATA_0_12), .DIN2(n3484) );
  nnd2s1 U8926 ( .Q(n5922), .DIN1(CRC_OUT_1_12), .DIN2(n3528) );
  nnd4s1 U8927 ( .Q(WX11024), .DIN1(n5928), .DIN2(n5929), .DIN3(n5930), .DIN4(
        n5931) );
  nnd2s1 U8928 ( .Q(n5931), .DIN1(n3434), .DIN2(n3675) );
  xor2s1 U8929 ( .Q(n3675), .DIN1(n5932), .DIN2(n5933) );
  xor2s1 U8930 ( .Q(n5933), .DIN1(n3090), .DIN2(WX11025) );
  xor2s1 U8931 ( .Q(n5932), .DIN1(n3330), .DIN2(WX11153) );
  nnd2s1 U8932 ( .Q(n5930), .DIN1(WX10865), .DIN2(n3496) );
  nnd2s1 U8933 ( .Q(n5929), .DIN1(DATA_0_13), .DIN2(n3484) );
  nnd2s1 U8934 ( .Q(n5928), .DIN1(CRC_OUT_1_13), .DIN2(n3528) );
  nnd4s1 U8935 ( .Q(WX11022), .DIN1(n5934), .DIN2(n5935), .DIN3(n5936), .DIN4(
        n5937) );
  nnd2s1 U8936 ( .Q(n5937), .DIN1(n3434), .DIN2(n3681) );
  xor2s1 U8937 ( .Q(n3681), .DIN1(n5938), .DIN2(n5939) );
  xor2s1 U8938 ( .Q(n5939), .DIN1(n3091), .DIN2(WX11023) );
  xor2s1 U8939 ( .Q(n5938), .DIN1(n3331), .DIN2(WX11151) );
  nnd2s1 U8940 ( .Q(n5936), .DIN1(WX10863), .DIN2(n3496) );
  nnd2s1 U8941 ( .Q(n5935), .DIN1(DATA_0_14), .DIN2(n3484) );
  nnd2s1 U8942 ( .Q(n5934), .DIN1(CRC_OUT_1_14), .DIN2(n3528) );
  nnd4s1 U8943 ( .Q(WX11020), .DIN1(n5940), .DIN2(n5941), .DIN3(n5942), .DIN4(
        n5943) );
  nnd2s1 U8944 ( .Q(n5943), .DIN1(n3434), .DIN2(n3687) );
  xor2s1 U8945 ( .Q(n3687), .DIN1(n5944), .DIN2(n5945) );
  xor2s1 U8946 ( .Q(n5945), .DIN1(n3092), .DIN2(WX11021) );
  xor2s1 U8947 ( .Q(n5944), .DIN1(n3332), .DIN2(WX11149) );
  nnd2s1 U8948 ( .Q(n5942), .DIN1(WX10861), .DIN2(n3496) );
  nnd2s1 U8949 ( .Q(n5941), .DIN1(DATA_0_15), .DIN2(n3484) );
  nnd2s1 U8950 ( .Q(n5940), .DIN1(CRC_OUT_1_15), .DIN2(n3528) );
  nnd4s1 U8951 ( .Q(WX11018), .DIN1(n5946), .DIN2(n5947), .DIN3(n5948), .DIN4(
        n5949) );
  nnd2s1 U8952 ( .Q(n5949), .DIN1(n3434), .DIN2(n3693) );
  xor2s1 U8953 ( .Q(n3693), .DIN1(n5950), .DIN2(n5951) );
  xor2s1 U8954 ( .Q(n5951), .DIN1(n3575), .DIN2(WX11019) );
  xor2s1 U8955 ( .Q(n5950), .DIN1(n3093), .DIN2(n5952) );
  xor2s1 U8956 ( .Q(n5952), .DIN1(WX11211), .DIN2(WX11147) );
  nnd2s1 U8957 ( .Q(n5948), .DIN1(WX10859), .DIN2(n3496) );
  nnd2s1 U8958 ( .Q(n5947), .DIN1(DATA_0_16), .DIN2(n3484) );
  nnd2s1 U8959 ( .Q(n5946), .DIN1(CRC_OUT_1_16), .DIN2(n3528) );
  nnd4s1 U8960 ( .Q(WX11016), .DIN1(n5953), .DIN2(n5954), .DIN3(n5955), .DIN4(
        n5956) );
  nnd2s1 U8961 ( .Q(n5956), .DIN1(n3434), .DIN2(n3699) );
  xor2s1 U8962 ( .Q(n3699), .DIN1(n5957), .DIN2(n5958) );
  xor2s1 U8963 ( .Q(n5958), .DIN1(n3575), .DIN2(WX11017) );
  xor2s1 U8964 ( .Q(n5957), .DIN1(n3094), .DIN2(n5959) );
  xor2s1 U8965 ( .Q(n5959), .DIN1(WX11209), .DIN2(WX11145) );
  nnd2s1 U8966 ( .Q(n5955), .DIN1(WX10857), .DIN2(n3496) );
  nnd2s1 U8967 ( .Q(n5954), .DIN1(DATA_0_17), .DIN2(n3485) );
  nnd2s1 U8968 ( .Q(n5953), .DIN1(CRC_OUT_1_17), .DIN2(n3528) );
  nnd4s1 U8969 ( .Q(WX11014), .DIN1(n5960), .DIN2(n5961), .DIN3(n5962), .DIN4(
        n5963) );
  nnd2s1 U8970 ( .Q(n5963), .DIN1(n3434), .DIN2(n3705) );
  xor2s1 U8971 ( .Q(n3705), .DIN1(n5964), .DIN2(n5965) );
  xor2s1 U8972 ( .Q(n5965), .DIN1(n3575), .DIN2(WX11015) );
  xor2s1 U8973 ( .Q(n5964), .DIN1(n3095), .DIN2(n5966) );
  xor2s1 U8974 ( .Q(n5966), .DIN1(WX11207), .DIN2(WX11143) );
  nnd2s1 U8975 ( .Q(n5962), .DIN1(WX10855), .DIN2(n3496) );
  nnd2s1 U8976 ( .Q(n5961), .DIN1(DATA_0_18), .DIN2(n3485) );
  nnd2s1 U8977 ( .Q(n5960), .DIN1(CRC_OUT_1_18), .DIN2(n3528) );
  nnd4s1 U8978 ( .Q(WX11012), .DIN1(n5967), .DIN2(n5968), .DIN3(n5969), .DIN4(
        n5970) );
  nnd2s1 U8979 ( .Q(n5970), .DIN1(n3433), .DIN2(n3711) );
  xor2s1 U8980 ( .Q(n3711), .DIN1(n5971), .DIN2(n5972) );
  xor2s1 U8981 ( .Q(n5972), .DIN1(n3575), .DIN2(WX11013) );
  xor2s1 U8982 ( .Q(n5971), .DIN1(n3096), .DIN2(n5973) );
  xor2s1 U8983 ( .Q(n5973), .DIN1(WX11205), .DIN2(WX11141) );
  nnd2s1 U8984 ( .Q(n5969), .DIN1(WX10853), .DIN2(n3496) );
  nnd2s1 U8985 ( .Q(n5968), .DIN1(DATA_0_19), .DIN2(n3485) );
  nnd2s1 U8986 ( .Q(n5967), .DIN1(CRC_OUT_1_19), .DIN2(n3528) );
  nnd4s1 U8987 ( .Q(WX11010), .DIN1(n5974), .DIN2(n5975), .DIN3(n5976), .DIN4(
        n5977) );
  nnd2s1 U8988 ( .Q(n5977), .DIN1(n3433), .DIN2(n3717) );
  xor2s1 U8989 ( .Q(n3717), .DIN1(n5978), .DIN2(n5979) );
  xor2s1 U8990 ( .Q(n5979), .DIN1(n3576), .DIN2(WX11011) );
  xor2s1 U8991 ( .Q(n5978), .DIN1(n3097), .DIN2(n5980) );
  xor2s1 U8992 ( .Q(n5980), .DIN1(WX11203), .DIN2(WX11139) );
  nnd2s1 U8993 ( .Q(n5976), .DIN1(WX10851), .DIN2(n3495) );
  nnd2s1 U8994 ( .Q(n5975), .DIN1(DATA_0_20), .DIN2(n3485) );
  nnd2s1 U8995 ( .Q(n5974), .DIN1(CRC_OUT_1_20), .DIN2(n3527) );
  xor2s1 U8996 ( .Q(WX1101), .DIN1(n4467), .DIN2(n5981) );
  nnd2s1 U8997 ( .Q(n5981), .DIN1(WX511), .DIN2(TM0) );
  xor2s1 U8998 ( .Q(n4467), .DIN1(n5982), .DIN2(n5983) );
  xor2s1 U8999 ( .Q(n5983), .DIN1(n3576), .DIN2(WX671) );
  xor2s1 U9000 ( .Q(n5982), .DIN1(WX735), .DIN2(n5984) );
  xor2s1 U9001 ( .Q(n5984), .DIN1(WX863), .DIN2(WX799) );
  nnd4s1 U9002 ( .Q(WX11008), .DIN1(n5985), .DIN2(n5986), .DIN3(n5987), .DIN4(
        n5988) );
  nnd2s1 U9003 ( .Q(n5988), .DIN1(n3433), .DIN2(n3723) );
  xor2s1 U9004 ( .Q(n3723), .DIN1(n5989), .DIN2(n5990) );
  xor2s1 U9005 ( .Q(n5990), .DIN1(n3576), .DIN2(WX11009) );
  xor2s1 U9006 ( .Q(n5989), .DIN1(n3098), .DIN2(n5991) );
  xor2s1 U9007 ( .Q(n5991), .DIN1(WX11201), .DIN2(WX11137) );
  nnd2s1 U9008 ( .Q(n5987), .DIN1(WX10849), .DIN2(n3495) );
  nnd2s1 U9009 ( .Q(n5986), .DIN1(DATA_0_21), .DIN2(n3485) );
  nnd2s1 U9010 ( .Q(n5985), .DIN1(CRC_OUT_1_21), .DIN2(n3527) );
  nnd4s1 U9011 ( .Q(WX11006), .DIN1(n5992), .DIN2(n5993), .DIN3(n5994), .DIN4(
        n5995) );
  nnd2s1 U9012 ( .Q(n5995), .DIN1(n3433), .DIN2(n3729) );
  xor2s1 U9013 ( .Q(n3729), .DIN1(n5996), .DIN2(n5997) );
  xor2s1 U9014 ( .Q(n5997), .DIN1(n3576), .DIN2(WX11007) );
  xor2s1 U9015 ( .Q(n5996), .DIN1(n3099), .DIN2(n5998) );
  xor2s1 U9016 ( .Q(n5998), .DIN1(WX11199), .DIN2(WX11135) );
  nnd2s1 U9017 ( .Q(n5994), .DIN1(WX10847), .DIN2(n3495) );
  nnd2s1 U9018 ( .Q(n5993), .DIN1(DATA_0_22), .DIN2(n3485) );
  nnd2s1 U9019 ( .Q(n5992), .DIN1(CRC_OUT_1_22), .DIN2(n3527) );
  nnd4s1 U9020 ( .Q(WX11004), .DIN1(n5999), .DIN2(n6000), .DIN3(n6001), .DIN4(
        n6002) );
  nnd2s1 U9021 ( .Q(n6002), .DIN1(n3433), .DIN2(n3735) );
  xor2s1 U9022 ( .Q(n3735), .DIN1(n6003), .DIN2(n6004) );
  xor2s1 U9023 ( .Q(n6004), .DIN1(n3576), .DIN2(WX11005) );
  xor2s1 U9024 ( .Q(n6003), .DIN1(n3100), .DIN2(n6005) );
  xor2s1 U9025 ( .Q(n6005), .DIN1(WX11197), .DIN2(WX11133) );
  nnd2s1 U9026 ( .Q(n6001), .DIN1(WX10845), .DIN2(n3495) );
  nnd2s1 U9027 ( .Q(n6000), .DIN1(DATA_0_23), .DIN2(n3485) );
  nnd2s1 U9028 ( .Q(n5999), .DIN1(CRC_OUT_1_23), .DIN2(n3527) );
  nnd4s1 U9029 ( .Q(WX11002), .DIN1(n6006), .DIN2(n6007), .DIN3(n6008), .DIN4(
        n6009) );
  nnd2s1 U9030 ( .Q(n6009), .DIN1(n3433), .DIN2(n3741) );
  xor2s1 U9031 ( .Q(n3741), .DIN1(n6010), .DIN2(n6011) );
  xor2s1 U9032 ( .Q(n6011), .DIN1(n3576), .DIN2(WX11003) );
  xor2s1 U9033 ( .Q(n6010), .DIN1(n3101), .DIN2(n6012) );
  xor2s1 U9034 ( .Q(n6012), .DIN1(WX11195), .DIN2(WX11131) );
  nnd2s1 U9035 ( .Q(n6008), .DIN1(WX10843), .DIN2(n3495) );
  nnd2s1 U9036 ( .Q(n6007), .DIN1(DATA_0_24), .DIN2(n3485) );
  nnd2s1 U9037 ( .Q(n6006), .DIN1(CRC_OUT_1_24), .DIN2(n3527) );
  nnd4s1 U9038 ( .Q(WX11000), .DIN1(n6013), .DIN2(n6014), .DIN3(n6015), .DIN4(
        n6016) );
  nnd2s1 U9039 ( .Q(n6016), .DIN1(n3433), .DIN2(n3747) );
  xor2s1 U9040 ( .Q(n3747), .DIN1(n6017), .DIN2(n6018) );
  xor2s1 U9041 ( .Q(n6018), .DIN1(n3576), .DIN2(WX11001) );
  xor2s1 U9042 ( .Q(n6017), .DIN1(n3102), .DIN2(n6019) );
  xor2s1 U9043 ( .Q(n6019), .DIN1(WX11193), .DIN2(WX11129) );
  nnd2s1 U9044 ( .Q(n6015), .DIN1(WX10841), .DIN2(n3495) );
  nnd2s1 U9045 ( .Q(n6014), .DIN1(DATA_0_25), .DIN2(n3485) );
  nnd2s1 U9046 ( .Q(n6013), .DIN1(CRC_OUT_1_25), .DIN2(n3527) );
  nnd4s1 U9047 ( .Q(WX10998), .DIN1(n6020), .DIN2(n6021), .DIN3(n6022), .DIN4(
        n6023) );
  nnd2s1 U9048 ( .Q(n6023), .DIN1(n3433), .DIN2(n3753) );
  xor2s1 U9049 ( .Q(n3753), .DIN1(n6024), .DIN2(n6025) );
  xor2s1 U9050 ( .Q(n6025), .DIN1(n3577), .DIN2(WX10999) );
  xor2s1 U9051 ( .Q(n6024), .DIN1(n3103), .DIN2(n6026) );
  xor2s1 U9052 ( .Q(n6026), .DIN1(WX11191), .DIN2(WX11127) );
  nnd2s1 U9053 ( .Q(n6022), .DIN1(WX10839), .DIN2(n3495) );
  nnd2s1 U9054 ( .Q(n6021), .DIN1(DATA_0_26), .DIN2(n3485) );
  nnd2s1 U9055 ( .Q(n6020), .DIN1(CRC_OUT_1_26), .DIN2(n3527) );
  nnd4s1 U9056 ( .Q(WX10996), .DIN1(n6027), .DIN2(n6028), .DIN3(n6029), .DIN4(
        n6030) );
  nnd2s1 U9057 ( .Q(n6030), .DIN1(n3433), .DIN2(n3759) );
  xor2s1 U9058 ( .Q(n3759), .DIN1(n6031), .DIN2(n6032) );
  xor2s1 U9059 ( .Q(n6032), .DIN1(n3577), .DIN2(WX10997) );
  xor2s1 U9060 ( .Q(n6031), .DIN1(n3104), .DIN2(n6033) );
  xor2s1 U9061 ( .Q(n6033), .DIN1(WX11189), .DIN2(WX11125) );
  nnd2s1 U9062 ( .Q(n6029), .DIN1(WX10837), .DIN2(n3495) );
  nnd2s1 U9063 ( .Q(n6028), .DIN1(DATA_0_27), .DIN2(n3485) );
  nnd2s1 U9064 ( .Q(n6027), .DIN1(CRC_OUT_1_27), .DIN2(n3527) );
  nnd4s1 U9065 ( .Q(WX10994), .DIN1(n6034), .DIN2(n6035), .DIN3(n6036), .DIN4(
        n6037) );
  nnd2s1 U9066 ( .Q(n6037), .DIN1(n3433), .DIN2(n3765) );
  xor2s1 U9067 ( .Q(n3765), .DIN1(n6038), .DIN2(n6039) );
  xor2s1 U9068 ( .Q(n6039), .DIN1(n3577), .DIN2(WX10995) );
  xor2s1 U9069 ( .Q(n6038), .DIN1(n3105), .DIN2(n6040) );
  xor2s1 U9070 ( .Q(n6040), .DIN1(WX11187), .DIN2(WX11123) );
  nnd2s1 U9071 ( .Q(n6036), .DIN1(WX10835), .DIN2(n3495) );
  nnd2s1 U9072 ( .Q(n6035), .DIN1(DATA_0_28), .DIN2(n3485) );
  nnd2s1 U9073 ( .Q(n6034), .DIN1(CRC_OUT_1_28), .DIN2(n3527) );
  nnd4s1 U9074 ( .Q(WX10992), .DIN1(n6041), .DIN2(n6042), .DIN3(n6043), .DIN4(
        n6044) );
  nnd2s1 U9075 ( .Q(n6044), .DIN1(n3433), .DIN2(n3771) );
  xor2s1 U9076 ( .Q(n3771), .DIN1(n6045), .DIN2(n6046) );
  xor2s1 U9077 ( .Q(n6046), .DIN1(n3577), .DIN2(WX10993) );
  xor2s1 U9078 ( .Q(n6045), .DIN1(n3106), .DIN2(n6047) );
  xor2s1 U9079 ( .Q(n6047), .DIN1(WX11185), .DIN2(WX11121) );
  nnd2s1 U9080 ( .Q(n6043), .DIN1(WX10833), .DIN2(n3495) );
  nnd2s1 U9081 ( .Q(n6042), .DIN1(DATA_0_29), .DIN2(n3485) );
  nnd2s1 U9082 ( .Q(n6041), .DIN1(CRC_OUT_1_29), .DIN2(n3527) );
  nnd4s1 U9083 ( .Q(WX10990), .DIN1(n6048), .DIN2(n6049), .DIN3(n6050), .DIN4(
        n6051) );
  nnd2s1 U9084 ( .Q(n6051), .DIN1(n3433), .DIN2(n3777) );
  xor2s1 U9085 ( .Q(n3777), .DIN1(n6052), .DIN2(n6053) );
  xor2s1 U9086 ( .Q(n6053), .DIN1(n3577), .DIN2(WX10991) );
  xor2s1 U9087 ( .Q(n6052), .DIN1(n3107), .DIN2(n6054) );
  xor2s1 U9088 ( .Q(n6054), .DIN1(WX11183), .DIN2(WX11119) );
  nnd2s1 U9089 ( .Q(n6050), .DIN1(WX10831), .DIN2(n3495) );
  nnd2s1 U9090 ( .Q(n6049), .DIN1(DATA_0_30), .DIN2(n3486) );
  nnd2s1 U9091 ( .Q(n6048), .DIN1(CRC_OUT_1_30), .DIN2(n3527) );
  nnd4s1 U9092 ( .Q(WX10988), .DIN1(n6055), .DIN2(n6056), .DIN3(n6057), .DIN4(
        n6058) );
  nnd2s1 U9093 ( .Q(n6058), .DIN1(WX10829), .DIN2(n3495) );
  and3s1 U9094 ( .Q(n3596), .DIN1(TM1), .DIN2(RESET), .DIN3(TM0) );
  nnd2s1 U9095 ( .Q(n6057), .DIN1(DATA_0_31), .DIN2(n3486) );
  and3s1 U9096 ( .Q(n3594), .DIN1(n3362), .DIN2(n3560), .DIN3(RESET) );
  nnd2s1 U9097 ( .Q(n6056), .DIN1(CRC_OUT_1_31), .DIN2(n3527) );
  and3s1 U9098 ( .Q(n3597), .DIN1(RESET), .DIN2(n3559), .DIN3(TM0) );
  nnd2s1 U9099 ( .Q(n6055), .DIN1(n3433), .DIN2(n3783) );
  xor2s1 U9100 ( .Q(n3783), .DIN1(n6059), .DIN2(n6060) );
  xor2s1 U9101 ( .Q(n6060), .DIN1(n3577), .DIN2(WX10989) );
  xor2s1 U9102 ( .Q(n6059), .DIN1(n3108), .DIN2(n6061) );
  xor2s1 U9103 ( .Q(n6061), .DIN1(WX11181), .DIN2(WX11117) );
  and3s1 U9104 ( .Q(n3592), .DIN1(RESET), .DIN2(n5745), .DIN3(TM1) );
  hi1s1 U9105 ( .Q(n5745), .DIN(TM0) );
  xor2s1 U9106 ( .Q(WX1094), .DIN1(n4474), .DIN2(n6062) );
  nnd2s1 U9107 ( .Q(n6062), .DIN1(WX509), .DIN2(TM0) );
  xor2s1 U9108 ( .Q(n4474), .DIN1(n6063), .DIN2(n6064) );
  xor2s1 U9109 ( .Q(n6064), .DIN1(n3578), .DIN2(WX669) );
  xor2s1 U9110 ( .Q(n6063), .DIN1(WX733), .DIN2(n6065) );
  xor2s1 U9111 ( .Q(n6065), .DIN1(WX861), .DIN2(WX797) );
  nor2s1 U9112 ( .Q(WX10890), .DIN1(WX10829), .DIN2(n3363) );
  and2s1 U9113 ( .Q(WX10888), .DIN1(RESET), .DIN2(WX10891) );
  and2s1 U9114 ( .Q(WX10886), .DIN1(RESET), .DIN2(WX10889) );
  and2s1 U9115 ( .Q(WX10884), .DIN1(RESET), .DIN2(WX10887) );
  and2s1 U9116 ( .Q(WX10882), .DIN1(RESET), .DIN2(WX10885) );
  and2s1 U9117 ( .Q(WX10880), .DIN1(RESET), .DIN2(WX10883) );
  and2s1 U9118 ( .Q(WX10878), .DIN1(RESET), .DIN2(WX10881) );
  and2s1 U9119 ( .Q(WX10876), .DIN1(RESET), .DIN2(WX10879) );
  and2s1 U9120 ( .Q(WX10874), .DIN1(RESET), .DIN2(WX10877) );
  and2s1 U9121 ( .Q(WX10872), .DIN1(RESET), .DIN2(WX10875) );
  and2s1 U9122 ( .Q(WX10870), .DIN1(RESET), .DIN2(WX10873) );
  xor2s1 U9123 ( .Q(WX1087), .DIN1(n4481), .DIN2(n6066) );
  nnd2s1 U9124 ( .Q(n6066), .DIN1(WX507), .DIN2(TM0) );
  xor2s1 U9125 ( .Q(n4481), .DIN1(n6067), .DIN2(n6068) );
  xor2s1 U9126 ( .Q(n6068), .DIN1(n3578), .DIN2(WX667) );
  xor2s1 U9127 ( .Q(n6067), .DIN1(WX731), .DIN2(n6069) );
  xor2s1 U9128 ( .Q(n6069), .DIN1(WX859), .DIN2(WX795) );
  and2s1 U9129 ( .Q(WX10868), .DIN1(RESET), .DIN2(WX10871) );
  and2s1 U9130 ( .Q(WX10866), .DIN1(RESET), .DIN2(WX10869) );
  and2s1 U9131 ( .Q(WX10864), .DIN1(RESET), .DIN2(WX10867) );
  and2s1 U9132 ( .Q(WX10862), .DIN1(RESET), .DIN2(WX10865) );
  and2s1 U9133 ( .Q(WX10860), .DIN1(RESET), .DIN2(WX10863) );
  and2s1 U9134 ( .Q(WX10858), .DIN1(RESET), .DIN2(WX10861) );
  and2s1 U9135 ( .Q(WX10856), .DIN1(RESET), .DIN2(WX10859) );
  and2s1 U9136 ( .Q(WX10854), .DIN1(RESET), .DIN2(WX10857) );
  and2s1 U9137 ( .Q(WX10852), .DIN1(RESET), .DIN2(WX10855) );
  and2s1 U9138 ( .Q(WX10850), .DIN1(RESET), .DIN2(WX10853) );
  and2s1 U9139 ( .Q(WX10848), .DIN1(RESET), .DIN2(WX10851) );
  and2s1 U9140 ( .Q(WX10846), .DIN1(RESET), .DIN2(WX10849) );
  and2s1 U9141 ( .Q(WX10844), .DIN1(RESET), .DIN2(WX10847) );
  and2s1 U9142 ( .Q(WX10842), .DIN1(RESET), .DIN2(WX10845) );
  and2s1 U9143 ( .Q(WX10840), .DIN1(RESET), .DIN2(WX10843) );
  and2s1 U9144 ( .Q(WX10838), .DIN1(RESET), .DIN2(WX10841) );
  and2s1 U9145 ( .Q(WX10836), .DIN1(RESET), .DIN2(WX10839) );
  and2s1 U9146 ( .Q(WX10834), .DIN1(RESET), .DIN2(WX10837) );
  and2s1 U9147 ( .Q(WX10832), .DIN1(RESET), .DIN2(WX10835) );
  and2s1 U9148 ( .Q(WX10830), .DIN1(RESET), .DIN2(WX10833) );
  and2s1 U9149 ( .Q(WX10828), .DIN1(RESET), .DIN2(WX10831) );
  xor2s1 U9150 ( .Q(WX1080), .DIN1(n4488), .DIN2(n6070) );
  nnd2s1 U9151 ( .Q(n6070), .DIN1(WX505), .DIN2(TM0) );
  xor2s1 U9152 ( .Q(n4488), .DIN1(n6071), .DIN2(n6072) );
  xor2s1 U9153 ( .Q(n6072), .DIN1(n3578), .DIN2(WX665) );
  xor2s1 U9154 ( .Q(n6071), .DIN1(WX729), .DIN2(n6073) );
  xor2s1 U9155 ( .Q(n6073), .DIN1(WX857), .DIN2(WX793) );
  xor2s1 U9156 ( .Q(WX1073), .DIN1(n4495), .DIN2(n6074) );
  nnd2s1 U9157 ( .Q(n6074), .DIN1(WX503), .DIN2(TM0) );
  xor2s1 U9158 ( .Q(n4495), .DIN1(n6075), .DIN2(n6076) );
  xor2s1 U9159 ( .Q(n6076), .DIN1(n3578), .DIN2(WX663) );
  xor2s1 U9160 ( .Q(n6075), .DIN1(WX727), .DIN2(n6077) );
  xor2s1 U9161 ( .Q(n6077), .DIN1(WX855), .DIN2(WX791) );
  xor2s1 U9162 ( .Q(WX1066), .DIN1(n4502), .DIN2(n6078) );
  nnd2s1 U9163 ( .Q(n6078), .DIN1(WX501), .DIN2(TM0) );
  xor2s1 U9164 ( .Q(n4502), .DIN1(n6079), .DIN2(n6080) );
  xor2s1 U9165 ( .Q(n6080), .DIN1(n3578), .DIN2(WX661) );
  xor2s1 U9166 ( .Q(n6079), .DIN1(WX725), .DIN2(n6081) );
  xor2s1 U9167 ( .Q(n6081), .DIN1(WX853), .DIN2(WX789) );
  xor2s1 U9168 ( .Q(WX1059), .DIN1(n4509), .DIN2(n6082) );
  nnd2s1 U9169 ( .Q(n6082), .DIN1(WX499), .DIN2(TM0) );
  xor2s1 U9170 ( .Q(n4509), .DIN1(n6083), .DIN2(n6084) );
  xor2s1 U9171 ( .Q(n6084), .DIN1(n3578), .DIN2(WX659) );
  xor2s1 U9172 ( .Q(n6083), .DIN1(WX723), .DIN2(n6085) );
  xor2s1 U9173 ( .Q(n6085), .DIN1(WX851), .DIN2(WX787) );
  xor2s1 U9174 ( .Q(WX1052), .DIN1(n4516), .DIN2(n6086) );
  nnd2s1 U9175 ( .Q(n6086), .DIN1(WX497), .DIN2(TM0) );
  xor2s1 U9176 ( .Q(n4516), .DIN1(n6087), .DIN2(n6088) );
  xor2s1 U9177 ( .Q(n6088), .DIN1(n3578), .DIN2(WX657) );
  xor2s1 U9178 ( .Q(n6087), .DIN1(WX721), .DIN2(n6089) );
  xor2s1 U9179 ( .Q(n6089), .DIN1(WX849), .DIN2(WX785) );
  xor2s1 U9180 ( .Q(WX1045), .DIN1(n4523), .DIN2(n6090) );
  nnd2s1 U9181 ( .Q(n6090), .DIN1(WX495), .DIN2(TM0) );
  xor2s1 U9182 ( .Q(n4523), .DIN1(n6091), .DIN2(n6092) );
  xor2s1 U9183 ( .Q(n6092), .DIN1(n3579), .DIN2(WX655) );
  xor2s1 U9184 ( .Q(n6091), .DIN1(WX719), .DIN2(n6093) );
  xor2s1 U9185 ( .Q(n6093), .DIN1(WX847), .DIN2(WX783) );
  xor2s1 U9186 ( .Q(WX1038), .DIN1(n4530), .DIN2(n6094) );
  nnd2s1 U9187 ( .Q(n6094), .DIN1(WX493), .DIN2(TM0) );
  xor2s1 U9188 ( .Q(n4530), .DIN1(n6095), .DIN2(n6096) );
  xor2s1 U9189 ( .Q(n6096), .DIN1(n3579), .DIN2(WX653) );
  xor2s1 U9190 ( .Q(n6095), .DIN1(WX717), .DIN2(n6097) );
  xor2s1 U9191 ( .Q(n6097), .DIN1(WX845), .DIN2(WX781) );
  nor2s1 U9192 ( .Q(WX10377), .DIN1(n3401), .DIN2(n6098) );
  xor2s1 U9193 ( .Q(n6098), .DIN1(WX9888), .DIN2(CRC_OUT_2_30) );
  nor2s1 U9194 ( .Q(WX10375), .DIN1(n3401), .DIN2(n6099) );
  xor2s1 U9195 ( .Q(n6099), .DIN1(WX9890), .DIN2(CRC_OUT_2_29) );
  nor2s1 U9196 ( .Q(WX10373), .DIN1(n3401), .DIN2(n6100) );
  xor2s1 U9197 ( .Q(n6100), .DIN1(WX9892), .DIN2(CRC_OUT_2_28) );
  nor2s1 U9198 ( .Q(WX10371), .DIN1(n3401), .DIN2(n6101) );
  xor2s1 U9199 ( .Q(n6101), .DIN1(WX9894), .DIN2(CRC_OUT_2_27) );
  nor2s1 U9200 ( .Q(WX10369), .DIN1(n3401), .DIN2(n6102) );
  xor2s1 U9201 ( .Q(n6102), .DIN1(WX9896), .DIN2(CRC_OUT_2_26) );
  nor2s1 U9202 ( .Q(WX10367), .DIN1(n3402), .DIN2(n6103) );
  xor2s1 U9203 ( .Q(n6103), .DIN1(WX9898), .DIN2(CRC_OUT_2_25) );
  nor2s1 U9204 ( .Q(WX10365), .DIN1(n3402), .DIN2(n6104) );
  xor2s1 U9205 ( .Q(n6104), .DIN1(WX9900), .DIN2(CRC_OUT_2_24) );
  nor2s1 U9206 ( .Q(WX10363), .DIN1(n3402), .DIN2(n6105) );
  xor2s1 U9207 ( .Q(n6105), .DIN1(WX9902), .DIN2(CRC_OUT_2_23) );
  nor2s1 U9208 ( .Q(WX10361), .DIN1(n3402), .DIN2(n6106) );
  xor2s1 U9209 ( .Q(n6106), .DIN1(WX9904), .DIN2(CRC_OUT_2_22) );
  nor2s1 U9210 ( .Q(WX10359), .DIN1(n3402), .DIN2(n6107) );
  xor2s1 U9211 ( .Q(n6107), .DIN1(WX9906), .DIN2(CRC_OUT_2_21) );
  nor2s1 U9212 ( .Q(WX10357), .DIN1(n3402), .DIN2(n6108) );
  xor2s1 U9213 ( .Q(n6108), .DIN1(WX9908), .DIN2(CRC_OUT_2_20) );
  nor2s1 U9214 ( .Q(WX10355), .DIN1(n3402), .DIN2(n6109) );
  xor2s1 U9215 ( .Q(n6109), .DIN1(WX9910), .DIN2(CRC_OUT_2_19) );
  nor2s1 U9216 ( .Q(WX10353), .DIN1(n3402), .DIN2(n6110) );
  xor2s1 U9217 ( .Q(n6110), .DIN1(WX9912), .DIN2(CRC_OUT_2_18) );
  nor2s1 U9218 ( .Q(WX10351), .DIN1(n3402), .DIN2(n6111) );
  xor2s1 U9219 ( .Q(n6111), .DIN1(WX9914), .DIN2(CRC_OUT_2_17) );
  nor2s1 U9220 ( .Q(WX10349), .DIN1(n3402), .DIN2(n6112) );
  xor2s1 U9221 ( .Q(n6112), .DIN1(WX9916), .DIN2(CRC_OUT_2_16) );
  nor2s1 U9222 ( .Q(WX10347), .DIN1(n3403), .DIN2(n6113) );
  xor2s1 U9223 ( .Q(n6113), .DIN1(CRC_OUT_2_15), .DIN2(n6114) );
  xor2s1 U9224 ( .Q(n6114), .DIN1(WX9918), .DIN2(CRC_OUT_2_31) );
  nor2s1 U9225 ( .Q(WX10345), .DIN1(n3403), .DIN2(n6115) );
  xor2s1 U9226 ( .Q(n6115), .DIN1(WX9920), .DIN2(CRC_OUT_2_14) );
  nor2s1 U9227 ( .Q(WX10343), .DIN1(n3403), .DIN2(n6116) );
  xor2s1 U9228 ( .Q(n6116), .DIN1(WX9922), .DIN2(CRC_OUT_2_13) );
  nor2s1 U9229 ( .Q(WX10341), .DIN1(n3403), .DIN2(n6117) );
  xor2s1 U9230 ( .Q(n6117), .DIN1(WX9924), .DIN2(CRC_OUT_2_12) );
  nor2s1 U9231 ( .Q(WX10339), .DIN1(n3403), .DIN2(n6118) );
  xor2s1 U9232 ( .Q(n6118), .DIN1(WX9926), .DIN2(CRC_OUT_2_11) );
  nor2s1 U9233 ( .Q(WX10337), .DIN1(n3403), .DIN2(n6119) );
  xor2s1 U9234 ( .Q(n6119), .DIN1(CRC_OUT_2_10), .DIN2(n6120) );
  xor2s1 U9235 ( .Q(n6120), .DIN1(WX9928), .DIN2(CRC_OUT_2_31) );
  nor2s1 U9236 ( .Q(WX10335), .DIN1(n3403), .DIN2(n6121) );
  xor2s1 U9237 ( .Q(n6121), .DIN1(WX9930), .DIN2(CRC_OUT_2_9) );
  nor2s1 U9238 ( .Q(WX10333), .DIN1(n3403), .DIN2(n6122) );
  xor2s1 U9239 ( .Q(n6122), .DIN1(WX9932), .DIN2(CRC_OUT_2_8) );
  nor2s1 U9240 ( .Q(WX10331), .DIN1(n3403), .DIN2(n6123) );
  xor2s1 U9241 ( .Q(n6123), .DIN1(WX9934), .DIN2(CRC_OUT_2_7) );
  nor2s1 U9242 ( .Q(WX10329), .DIN1(n3403), .DIN2(n6124) );
  xor2s1 U9243 ( .Q(n6124), .DIN1(WX9936), .DIN2(CRC_OUT_2_6) );
  nor2s1 U9244 ( .Q(WX10327), .DIN1(n3404), .DIN2(n6125) );
  xor2s1 U9245 ( .Q(n6125), .DIN1(WX9938), .DIN2(CRC_OUT_2_5) );
  nor2s1 U9246 ( .Q(WX10325), .DIN1(n3404), .DIN2(n6126) );
  xor2s1 U9247 ( .Q(n6126), .DIN1(WX9940), .DIN2(CRC_OUT_2_4) );
  nor2s1 U9248 ( .Q(WX10323), .DIN1(n3404), .DIN2(n6127) );
  xor2s1 U9249 ( .Q(n6127), .DIN1(CRC_OUT_2_3), .DIN2(n6128) );
  xor2s1 U9250 ( .Q(n6128), .DIN1(WX9942), .DIN2(CRC_OUT_2_31) );
  nor2s1 U9251 ( .Q(WX10321), .DIN1(n3404), .DIN2(n6129) );
  xor2s1 U9252 ( .Q(n6129), .DIN1(WX9944), .DIN2(CRC_OUT_2_2) );
  nor2s1 U9253 ( .Q(WX10319), .DIN1(n3404), .DIN2(n6130) );
  xor2s1 U9254 ( .Q(n6130), .DIN1(WX9946), .DIN2(CRC_OUT_2_1) );
  nor2s1 U9255 ( .Q(WX10317), .DIN1(n3404), .DIN2(n6131) );
  xor2s1 U9256 ( .Q(n6131), .DIN1(WX9948), .DIN2(CRC_OUT_2_0) );
  nor2s1 U9257 ( .Q(WX10315), .DIN1(n3365), .DIN2(n6132) );
  xor2s1 U9258 ( .Q(n6132), .DIN1(WX9950), .DIN2(CRC_OUT_2_31) );
  hi1s1 U9259 ( .Q(n3587), .DIN(RESET) );
  xor2s1 U9260 ( .Q(WX1031), .DIN1(n4537), .DIN2(n6133) );
  nnd2s1 U9261 ( .Q(n6133), .DIN1(WX491), .DIN2(TM0) );
  xor2s1 U9262 ( .Q(n4537), .DIN1(n6134), .DIN2(n6135) );
  xor2s1 U9263 ( .Q(n6135), .DIN1(n3579), .DIN2(WX651) );
  xor2s1 U9264 ( .Q(n6134), .DIN1(WX715), .DIN2(n6136) );
  xor2s1 U9265 ( .Q(n6136), .DIN1(WX843), .DIN2(WX779) );
  xor2s1 U9266 ( .Q(WX1024), .DIN1(n4554), .DIN2(n6137) );
  nnd2s1 U9267 ( .Q(n6137), .DIN1(WX489), .DIN2(TM0) );
  xor2s1 U9268 ( .Q(n4554), .DIN1(n6138), .DIN2(n6139) );
  xor2s1 U9269 ( .Q(n6139), .DIN1(n3579), .DIN2(WX649) );
  xor2s1 U9270 ( .Q(n6138), .DIN1(WX713), .DIN2(n6140) );
  xor2s1 U9271 ( .Q(n6140), .DIN1(WX841), .DIN2(WX777) );
  xor2s1 U9272 ( .Q(WX1017), .DIN1(n4572), .DIN2(n6141) );
  nnd2s1 U9273 ( .Q(n6141), .DIN1(WX487), .DIN2(TM0) );
  xor2s1 U9274 ( .Q(n4572), .DIN1(n6142), .DIN2(n6143) );
  xor2s1 U9275 ( .Q(n6143), .DIN1(n3577), .DIN2(WX647) );
  xor2s1 U9276 ( .Q(n6142), .DIN1(WX711), .DIN2(n6144) );
  xor2s1 U9277 ( .Q(n6144), .DIN1(WX839), .DIN2(WX775) );
  xor2s1 U9278 ( .Q(WX1010), .DIN1(n4591), .DIN2(n6145) );
  nnd2s1 U9279 ( .Q(n6145), .DIN1(WX485), .DIN2(TM0) );
  xor2s1 U9280 ( .Q(n4591), .DIN1(n6146), .DIN2(n3358) );
  xor2s1 U9281 ( .Q(n6147), .DIN1(n3559), .DIN2(WX645) );
  hi1s1 U9282 ( .Q(n3937), .DIN(TM1) );
  xor2s1 U9283 ( .Q(n6146), .DIN1(WX709), .DIN2(n6148) );
  xor2s1 U9284 ( .Q(n6148), .DIN1(WX837), .DIN2(WX773) );
  dffs1 \DFF_1727/Q_reg  ( .Q(CRC_OUT_1_31), .CLK(CK), .DIN(WX11670) );
  dffs1 \DFF_1726/Q_reg  ( .Q(CRC_OUT_1_30), .CLK(CK), .DIN(WX11668) );
  dffs1 \DFF_1725/Q_reg  ( .Q(CRC_OUT_1_29), .CLK(CK), .DIN(WX11666) );
  dffs1 \DFF_1724/Q_reg  ( .Q(CRC_OUT_1_28), .CLK(CK), .DIN(WX11664) );
  dffs1 \DFF_1723/Q_reg  ( .Q(CRC_OUT_1_27), .CLK(CK), .DIN(WX11662) );
  dffs1 \DFF_1722/Q_reg  ( .Q(CRC_OUT_1_26), .CLK(CK), .DIN(WX11660) );
  dffs1 \DFF_1721/Q_reg  ( .Q(CRC_OUT_1_25), .CLK(CK), .DIN(WX11658) );
  dffs1 \DFF_1720/Q_reg  ( .Q(CRC_OUT_1_24), .CLK(CK), .DIN(WX11656) );
  dffs1 \DFF_1719/Q_reg  ( .Q(CRC_OUT_1_23), .CLK(CK), .DIN(WX11654) );
  dffs1 \DFF_1718/Q_reg  ( .Q(CRC_OUT_1_22), .CLK(CK), .DIN(WX11652) );
  dffs1 \DFF_1717/Q_reg  ( .Q(CRC_OUT_1_21), .CLK(CK), .DIN(WX11650) );
  dffs1 \DFF_1716/Q_reg  ( .Q(CRC_OUT_1_20), .CLK(CK), .DIN(WX11648) );
  dffs1 \DFF_1715/Q_reg  ( .Q(CRC_OUT_1_19), .CLK(CK), .DIN(WX11646) );
  dffs1 \DFF_1714/Q_reg  ( .Q(CRC_OUT_1_18), .CLK(CK), .DIN(WX11644) );
  dffs1 \DFF_1713/Q_reg  ( .Q(CRC_OUT_1_17), .CLK(CK), .DIN(WX11642) );
  dffs1 \DFF_1712/Q_reg  ( .Q(CRC_OUT_1_16), .CLK(CK), .DIN(WX11640) );
  dffs1 \DFF_1711/Q_reg  ( .Q(CRC_OUT_1_15), .CLK(CK), .DIN(WX11638) );
  dffs1 \DFF_1710/Q_reg  ( .Q(CRC_OUT_1_14), .CLK(CK), .DIN(WX11636) );
  dffs1 \DFF_1709/Q_reg  ( .Q(CRC_OUT_1_13), .CLK(CK), .DIN(WX11634) );
  dffs1 \DFF_1708/Q_reg  ( .Q(CRC_OUT_1_12), .CLK(CK), .DIN(WX11632) );
  dffs1 \DFF_1707/Q_reg  ( .Q(CRC_OUT_1_11), .CLK(CK), .DIN(WX11630) );
  dffs1 \DFF_1706/Q_reg  ( .Q(CRC_OUT_1_10), .CLK(CK), .DIN(WX11628) );
  dffs1 \DFF_1705/Q_reg  ( .Q(CRC_OUT_1_9), .CLK(CK), .DIN(WX11626) );
  dffs1 \DFF_1704/Q_reg  ( .Q(CRC_OUT_1_8), .CLK(CK), .DIN(WX11624) );
  dffs1 \DFF_1703/Q_reg  ( .Q(CRC_OUT_1_7), .CLK(CK), .DIN(WX11622) );
  dffs1 \DFF_1702/Q_reg  ( .Q(CRC_OUT_1_6), .CLK(CK), .DIN(WX11620) );
  dffs1 \DFF_1701/Q_reg  ( .Q(CRC_OUT_1_5), .CLK(CK), .DIN(WX11618) );
  dffs1 \DFF_1700/Q_reg  ( .Q(CRC_OUT_1_4), .CLK(CK), .DIN(WX11616) );
  dffs1 \DFF_1699/Q_reg  ( .Q(CRC_OUT_1_3), .CLK(CK), .DIN(WX11614) );
  dffs1 \DFF_1698/Q_reg  ( .Q(CRC_OUT_1_2), .CLK(CK), .DIN(WX11612) );
  dffs1 \DFF_1697/Q_reg  ( .Q(CRC_OUT_1_1), .CLK(CK), .DIN(WX11610) );
  dffs1 \DFF_1696/Q_reg  ( .Q(CRC_OUT_1_0), .CLK(CK), .DIN(WX11608) );
  dffs1 \DFF_1695/Q_reg  ( .QN(n3317), .Q(WX11243), .CLK(CK), .DIN(WX11242) );
  dffs1 \DFF_1694/Q_reg  ( .QN(n3318), .Q(WX11241), .CLK(CK), .DIN(WX11240) );
  dffs1 \DFF_1693/Q_reg  ( .QN(n3319), .Q(WX11239), .CLK(CK), .DIN(WX11238) );
  dffs1 \DFF_1692/Q_reg  ( .QN(n3320), .Q(WX11237), .CLK(CK), .DIN(WX11236) );
  dffs1 \DFF_1691/Q_reg  ( .QN(n3321), .Q(WX11235), .CLK(CK), .DIN(WX11234) );
  dffs1 \DFF_1690/Q_reg  ( .QN(n3322), .Q(WX11233), .CLK(CK), .DIN(WX11232) );
  dffs1 \DFF_1689/Q_reg  ( .QN(n3323), .Q(WX11231), .CLK(CK), .DIN(WX11230) );
  dffs1 \DFF_1688/Q_reg  ( .QN(n3324), .Q(WX11229), .CLK(CK), .DIN(WX11228) );
  dffs1 \DFF_1687/Q_reg  ( .QN(n3325), .Q(WX11227), .CLK(CK), .DIN(WX11226) );
  dffs1 \DFF_1686/Q_reg  ( .QN(n3326), .Q(WX11225), .CLK(CK), .DIN(WX11224) );
  dffs1 \DFF_1685/Q_reg  ( .QN(n3327), .Q(WX11223), .CLK(CK), .DIN(WX11222) );
  dffs1 \DFF_1684/Q_reg  ( .QN(n3328), .Q(WX11221), .CLK(CK), .DIN(WX11220) );
  dffs1 \DFF_1683/Q_reg  ( .QN(n3329), .Q(WX11219), .CLK(CK), .DIN(WX11218) );
  dffs1 \DFF_1682/Q_reg  ( .QN(n3330), .Q(WX11217), .CLK(CK), .DIN(WX11216) );
  dffs1 \DFF_1681/Q_reg  ( .QN(n3331), .Q(WX11215), .CLK(CK), .DIN(WX11214) );
  dffs1 \DFF_1680/Q_reg  ( .QN(n3332), .Q(WX11213), .CLK(CK), .DIN(WX11212) );
  dffs1 \DFF_1679/Q_reg  ( .Q(WX11211), .CLK(CK), .DIN(WX11210) );
  dffs1 \DFF_1678/Q_reg  ( .Q(WX11209), .CLK(CK), .DIN(WX11208) );
  dffs1 \DFF_1677/Q_reg  ( .Q(WX11207), .CLK(CK), .DIN(WX11206) );
  dffs1 \DFF_1676/Q_reg  ( .Q(WX11205), .CLK(CK), .DIN(WX11204) );
  dffs1 \DFF_1675/Q_reg  ( .Q(WX11203), .CLK(CK), .DIN(WX11202) );
  dffs1 \DFF_1674/Q_reg  ( .Q(WX11201), .CLK(CK), .DIN(WX11200) );
  dffs1 \DFF_1673/Q_reg  ( .Q(WX11199), .CLK(CK), .DIN(WX11198) );
  dffs1 \DFF_1672/Q_reg  ( .Q(WX11197), .CLK(CK), .DIN(WX11196) );
  dffs1 \DFF_1671/Q_reg  ( .Q(WX11195), .CLK(CK), .DIN(WX11194) );
  dffs1 \DFF_1670/Q_reg  ( .Q(WX11193), .CLK(CK), .DIN(WX11192) );
  dffs1 \DFF_1669/Q_reg  ( .Q(WX11191), .CLK(CK), .DIN(WX11190) );
  dffs1 \DFF_1668/Q_reg  ( .Q(WX11189), .CLK(CK), .DIN(WX11188) );
  dffs1 \DFF_1667/Q_reg  ( .Q(WX11187), .CLK(CK), .DIN(WX11186) );
  dffs1 \DFF_1666/Q_reg  ( .Q(WX11185), .CLK(CK), .DIN(WX11184) );
  dffs1 \DFF_1665/Q_reg  ( .Q(WX11183), .CLK(CK), .DIN(WX11182) );
  dffs1 \DFF_1664/Q_reg  ( .Q(WX11181), .CLK(CK), .DIN(WX11180) );
  dffs1 \DFF_1663/Q_reg  ( .Q(WX11179), .CLK(CK), .DIN(WX11178) );
  dffs1 \DFF_1662/Q_reg  ( .Q(WX11177), .CLK(CK), .DIN(WX11176) );
  dffs1 \DFF_1661/Q_reg  ( .Q(WX11175), .CLK(CK), .DIN(WX11174) );
  dffs1 \DFF_1660/Q_reg  ( .Q(WX11173), .CLK(CK), .DIN(WX11172) );
  dffs1 \DFF_1659/Q_reg  ( .Q(WX11171), .CLK(CK), .DIN(WX11170) );
  dffs1 \DFF_1658/Q_reg  ( .Q(WX11169), .CLK(CK), .DIN(WX11168) );
  dffs1 \DFF_1657/Q_reg  ( .Q(WX11167), .CLK(CK), .DIN(WX11166) );
  dffs1 \DFF_1656/Q_reg  ( .Q(WX11165), .CLK(CK), .DIN(WX11164) );
  dffs1 \DFF_1655/Q_reg  ( .Q(WX11163), .CLK(CK), .DIN(WX11162) );
  dffs1 \DFF_1654/Q_reg  ( .Q(WX11161), .CLK(CK), .DIN(WX11160) );
  dffs1 \DFF_1653/Q_reg  ( .Q(WX11159), .CLK(CK), .DIN(WX11158) );
  dffs1 \DFF_1652/Q_reg  ( .Q(WX11157), .CLK(CK), .DIN(WX11156) );
  dffs1 \DFF_1651/Q_reg  ( .Q(WX11155), .CLK(CK), .DIN(WX11154) );
  dffs1 \DFF_1650/Q_reg  ( .Q(WX11153), .CLK(CK), .DIN(WX11152) );
  dffs1 \DFF_1649/Q_reg  ( .Q(WX11151), .CLK(CK), .DIN(WX11150) );
  dffs1 \DFF_1648/Q_reg  ( .Q(WX11149), .CLK(CK), .DIN(WX11148) );
  dffs1 \DFF_1647/Q_reg  ( .Q(WX11147), .CLK(CK), .DIN(WX11146) );
  dffs1 \DFF_1646/Q_reg  ( .Q(WX11145), .CLK(CK), .DIN(WX11144) );
  dffs1 \DFF_1645/Q_reg  ( .Q(WX11143), .CLK(CK), .DIN(WX11142) );
  dffs1 \DFF_1644/Q_reg  ( .Q(WX11141), .CLK(CK), .DIN(WX11140) );
  dffs1 \DFF_1643/Q_reg  ( .Q(WX11139), .CLK(CK), .DIN(WX11138) );
  dffs1 \DFF_1642/Q_reg  ( .Q(WX11137), .CLK(CK), .DIN(WX11136) );
  dffs1 \DFF_1641/Q_reg  ( .Q(WX11135), .CLK(CK), .DIN(WX11134) );
  dffs1 \DFF_1640/Q_reg  ( .Q(WX11133), .CLK(CK), .DIN(WX11132) );
  dffs1 \DFF_1639/Q_reg  ( .Q(WX11131), .CLK(CK), .DIN(WX11130) );
  dffs1 \DFF_1638/Q_reg  ( .Q(WX11129), .CLK(CK), .DIN(WX11128) );
  dffs1 \DFF_1637/Q_reg  ( .Q(WX11127), .CLK(CK), .DIN(WX11126) );
  dffs1 \DFF_1636/Q_reg  ( .Q(WX11125), .CLK(CK), .DIN(WX11124) );
  dffs1 \DFF_1635/Q_reg  ( .Q(WX11123), .CLK(CK), .DIN(WX11122) );
  dffs1 \DFF_1634/Q_reg  ( .Q(WX11121), .CLK(CK), .DIN(WX11120) );
  dffs1 \DFF_1633/Q_reg  ( .Q(WX11119), .CLK(CK), .DIN(WX11118) );
  dffs1 \DFF_1632/Q_reg  ( .Q(WX11117), .CLK(CK), .DIN(WX11116) );
  dffs1 \DFF_1631/Q_reg  ( .QN(n3077), .CLK(CK), .DIN(WX11114) );
  dffs1 \DFF_1630/Q_reg  ( .QN(n3078), .CLK(CK), .DIN(WX11112) );
  dffs1 \DFF_1629/Q_reg  ( .QN(n3079), .CLK(CK), .DIN(WX11110) );
  dffs1 \DFF_1628/Q_reg  ( .QN(n3080), .CLK(CK), .DIN(WX11108) );
  dffs1 \DFF_1627/Q_reg  ( .QN(n3081), .CLK(CK), .DIN(WX11106) );
  dffs1 \DFF_1626/Q_reg  ( .QN(n3082), .CLK(CK), .DIN(WX11104) );
  dffs1 \DFF_1625/Q_reg  ( .QN(n3083), .CLK(CK), .DIN(WX11102) );
  dffs1 \DFF_1624/Q_reg  ( .QN(n3084), .CLK(CK), .DIN(WX11100) );
  dffs1 \DFF_1623/Q_reg  ( .QN(n3085), .CLK(CK), .DIN(WX11098) );
  dffs1 \DFF_1622/Q_reg  ( .QN(n3086), .CLK(CK), .DIN(WX11096) );
  dffs1 \DFF_1621/Q_reg  ( .QN(n3087), .CLK(CK), .DIN(WX11094) );
  dffs1 \DFF_1620/Q_reg  ( .QN(n3088), .CLK(CK), .DIN(WX11092) );
  dffs1 \DFF_1619/Q_reg  ( .QN(n3089), .CLK(CK), .DIN(WX11090) );
  dffs1 \DFF_1618/Q_reg  ( .QN(n3090), .CLK(CK), .DIN(WX11088) );
  dffs1 \DFF_1617/Q_reg  ( .QN(n3091), .CLK(CK), .DIN(WX11086) );
  dffs1 \DFF_1616/Q_reg  ( .QN(n3092), .CLK(CK), .DIN(WX11084) );
  dffs1 \DFF_1615/Q_reg  ( .QN(n3093), .CLK(CK), .DIN(WX11082) );
  dffs1 \DFF_1614/Q_reg  ( .QN(n3094), .CLK(CK), .DIN(WX11080) );
  dffs1 \DFF_1613/Q_reg  ( .QN(n3095), .CLK(CK), .DIN(WX11078) );
  dffs1 \DFF_1612/Q_reg  ( .QN(n3096), .CLK(CK), .DIN(WX11076) );
  dffs1 \DFF_1611/Q_reg  ( .QN(n3097), .CLK(CK), .DIN(WX11074) );
  dffs1 \DFF_1610/Q_reg  ( .QN(n3098), .CLK(CK), .DIN(WX11072) );
  dffs1 \DFF_1609/Q_reg  ( .QN(n3099), .CLK(CK), .DIN(WX11070) );
  dffs1 \DFF_1608/Q_reg  ( .QN(n3100), .CLK(CK), .DIN(WX11068) );
  dffs1 \DFF_1607/Q_reg  ( .QN(n3101), .CLK(CK), .DIN(WX11066) );
  dffs1 \DFF_1606/Q_reg  ( .QN(n3102), .CLK(CK), .DIN(WX11064) );
  dffs1 \DFF_1605/Q_reg  ( .QN(n3103), .CLK(CK), .DIN(WX11062) );
  dffs1 \DFF_1604/Q_reg  ( .QN(n3104), .CLK(CK), .DIN(WX11060) );
  dffs1 \DFF_1603/Q_reg  ( .QN(n3105), .CLK(CK), .DIN(WX11058) );
  dffs1 \DFF_1602/Q_reg  ( .QN(n3106), .CLK(CK), .DIN(WX11056) );
  dffs1 \DFF_1601/Q_reg  ( .QN(n3107), .CLK(CK), .DIN(WX11054) );
  dffs1 \DFF_1600/Q_reg  ( .QN(n3108), .CLK(CK), .DIN(WX11052) );
  dffs1 \DFF_1599/Q_reg  ( .Q(WX11051), .CLK(CK), .DIN(WX11050) );
  dffs1 \DFF_1598/Q_reg  ( .Q(WX11049), .CLK(CK), .DIN(WX11048) );
  dffs1 \DFF_1597/Q_reg  ( .Q(WX11047), .CLK(CK), .DIN(WX11046) );
  dffs1 \DFF_1596/Q_reg  ( .Q(WX11045), .CLK(CK), .DIN(WX11044) );
  dffs1 \DFF_1595/Q_reg  ( .Q(WX11043), .CLK(CK), .DIN(WX11042) );
  dffs1 \DFF_1594/Q_reg  ( .Q(WX11041), .CLK(CK), .DIN(WX11040) );
  dffs1 \DFF_1593/Q_reg  ( .Q(WX11039), .CLK(CK), .DIN(WX11038) );
  dffs1 \DFF_1592/Q_reg  ( .Q(WX11037), .CLK(CK), .DIN(WX11036) );
  dffs1 \DFF_1591/Q_reg  ( .Q(WX11035), .CLK(CK), .DIN(WX11034) );
  dffs1 \DFF_1590/Q_reg  ( .Q(WX11033), .CLK(CK), .DIN(WX11032) );
  dffs1 \DFF_1589/Q_reg  ( .Q(WX11031), .CLK(CK), .DIN(WX11030) );
  dffs1 \DFF_1588/Q_reg  ( .Q(WX11029), .CLK(CK), .DIN(WX11028) );
  dffs1 \DFF_1587/Q_reg  ( .Q(WX11027), .CLK(CK), .DIN(WX11026) );
  dffs1 \DFF_1586/Q_reg  ( .Q(WX11025), .CLK(CK), .DIN(WX11024) );
  dffs1 \DFF_1585/Q_reg  ( .Q(WX11023), .CLK(CK), .DIN(WX11022) );
  dffs1 \DFF_1584/Q_reg  ( .Q(WX11021), .CLK(CK), .DIN(WX11020) );
  dffs1 \DFF_1583/Q_reg  ( .Q(WX11019), .CLK(CK), .DIN(WX11018) );
  dffs1 \DFF_1582/Q_reg  ( .Q(WX11017), .CLK(CK), .DIN(WX11016) );
  dffs1 \DFF_1581/Q_reg  ( .Q(WX11015), .CLK(CK), .DIN(WX11014) );
  dffs1 \DFF_1580/Q_reg  ( .Q(WX11013), .CLK(CK), .DIN(WX11012) );
  dffs1 \DFF_1579/Q_reg  ( .Q(WX11011), .CLK(CK), .DIN(WX11010) );
  dffs1 \DFF_1578/Q_reg  ( .Q(WX11009), .CLK(CK), .DIN(WX11008) );
  dffs1 \DFF_1577/Q_reg  ( .Q(WX11007), .CLK(CK), .DIN(WX11006) );
  dffs1 \DFF_1576/Q_reg  ( .Q(WX11005), .CLK(CK), .DIN(WX11004) );
  dffs1 \DFF_1575/Q_reg  ( .Q(WX11003), .CLK(CK), .DIN(WX11002) );
  dffs1 \DFF_1574/Q_reg  ( .Q(WX11001), .CLK(CK), .DIN(WX11000) );
  dffs1 \DFF_1573/Q_reg  ( .Q(WX10999), .CLK(CK), .DIN(WX10998) );
  dffs1 \DFF_1572/Q_reg  ( .Q(WX10997), .CLK(CK), .DIN(WX10996) );
  dffs1 \DFF_1571/Q_reg  ( .Q(WX10995), .CLK(CK), .DIN(WX10994) );
  dffs1 \DFF_1570/Q_reg  ( .Q(WX10993), .CLK(CK), .DIN(WX10992) );
  dffs1 \DFF_1569/Q_reg  ( .Q(WX10991), .CLK(CK), .DIN(WX10990) );
  dffs1 \DFF_1568/Q_reg  ( .Q(WX10989), .CLK(CK), .DIN(WX10988) );
  dffs1 \DFF_1567/Q_reg  ( .Q(WX10891), .CLK(CK), .DIN(WX10890) );
  dffs1 \DFF_1566/Q_reg  ( .Q(WX10889), .CLK(CK), .DIN(WX10888) );
  dffs1 \DFF_1565/Q_reg  ( .Q(WX10887), .CLK(CK), .DIN(WX10886) );
  dffs1 \DFF_1564/Q_reg  ( .Q(WX10885), .CLK(CK), .DIN(WX10884) );
  dffs1 \DFF_1563/Q_reg  ( .Q(WX10883), .CLK(CK), .DIN(WX10882) );
  dffs1 \DFF_1562/Q_reg  ( .Q(WX10881), .CLK(CK), .DIN(WX10880) );
  dffs1 \DFF_1561/Q_reg  ( .Q(WX10879), .CLK(CK), .DIN(WX10878) );
  dffs1 \DFF_1560/Q_reg  ( .Q(WX10877), .CLK(CK), .DIN(WX10876) );
  dffs1 \DFF_1559/Q_reg  ( .Q(WX10875), .CLK(CK), .DIN(WX10874) );
  dffs1 \DFF_1558/Q_reg  ( .Q(WX10873), .CLK(CK), .DIN(WX10872) );
  dffs1 \DFF_1557/Q_reg  ( .Q(WX10871), .CLK(CK), .DIN(WX10870) );
  dffs1 \DFF_1556/Q_reg  ( .Q(WX10869), .CLK(CK), .DIN(WX10868) );
  dffs1 \DFF_1555/Q_reg  ( .Q(WX10867), .CLK(CK), .DIN(WX10866) );
  dffs1 \DFF_1554/Q_reg  ( .Q(WX10865), .CLK(CK), .DIN(WX10864) );
  dffs1 \DFF_1553/Q_reg  ( .Q(WX10863), .CLK(CK), .DIN(WX10862) );
  dffs1 \DFF_1552/Q_reg  ( .Q(WX10861), .CLK(CK), .DIN(WX10860) );
  dffs1 \DFF_1551/Q_reg  ( .Q(WX10859), .CLK(CK), .DIN(WX10858) );
  dffs1 \DFF_1550/Q_reg  ( .Q(WX10857), .CLK(CK), .DIN(WX10856) );
  dffs1 \DFF_1549/Q_reg  ( .Q(WX10855), .CLK(CK), .DIN(WX10854) );
  dffs1 \DFF_1548/Q_reg  ( .Q(WX10853), .CLK(CK), .DIN(WX10852) );
  dffs1 \DFF_1547/Q_reg  ( .Q(WX10851), .CLK(CK), .DIN(WX10850) );
  dffs1 \DFF_1546/Q_reg  ( .Q(WX10849), .CLK(CK), .DIN(WX10848) );
  dffs1 \DFF_1545/Q_reg  ( .Q(WX10847), .CLK(CK), .DIN(WX10846) );
  dffs1 \DFF_1544/Q_reg  ( .Q(WX10845), .CLK(CK), .DIN(WX10844) );
  dffs1 \DFF_1543/Q_reg  ( .Q(WX10843), .CLK(CK), .DIN(WX10842) );
  dffs1 \DFF_1542/Q_reg  ( .Q(WX10841), .CLK(CK), .DIN(WX10840) );
  dffs1 \DFF_1541/Q_reg  ( .Q(WX10839), .CLK(CK), .DIN(WX10838) );
  dffs1 \DFF_1540/Q_reg  ( .Q(WX10837), .CLK(CK), .DIN(WX10836) );
  dffs1 \DFF_1539/Q_reg  ( .Q(WX10835), .CLK(CK), .DIN(WX10834) );
  dffs1 \DFF_1538/Q_reg  ( .Q(WX10833), .CLK(CK), .DIN(WX10832) );
  dffs1 \DFF_1537/Q_reg  ( .Q(WX10831), .CLK(CK), .DIN(WX10830) );
  dffs1 \DFF_1536/Q_reg  ( .Q(WX10829), .CLK(CK), .DIN(WX10828) );
  dffs1 \DFF_1535/Q_reg  ( .Q(CRC_OUT_2_31), .CLK(CK), .DIN(WX10377) );
  dffs1 \DFF_1534/Q_reg  ( .Q(CRC_OUT_2_30), .CLK(CK), .DIN(WX10375) );
  dffs1 \DFF_1533/Q_reg  ( .Q(CRC_OUT_2_29), .CLK(CK), .DIN(WX10373) );
  dffs1 \DFF_1532/Q_reg  ( .Q(CRC_OUT_2_28), .CLK(CK), .DIN(WX10371) );
  dffs1 \DFF_1531/Q_reg  ( .Q(CRC_OUT_2_27), .CLK(CK), .DIN(WX10369) );
  dffs1 \DFF_1530/Q_reg  ( .Q(CRC_OUT_2_26), .CLK(CK), .DIN(WX10367) );
  dffs1 \DFF_1529/Q_reg  ( .Q(CRC_OUT_2_25), .CLK(CK), .DIN(WX10365) );
  dffs1 \DFF_1528/Q_reg  ( .Q(CRC_OUT_2_24), .CLK(CK), .DIN(WX10363) );
  dffs1 \DFF_1527/Q_reg  ( .Q(CRC_OUT_2_23), .CLK(CK), .DIN(WX10361) );
  dffs1 \DFF_1526/Q_reg  ( .Q(CRC_OUT_2_22), .CLK(CK), .DIN(WX10359) );
  dffs1 \DFF_1525/Q_reg  ( .Q(CRC_OUT_2_21), .CLK(CK), .DIN(WX10357) );
  dffs1 \DFF_1524/Q_reg  ( .Q(CRC_OUT_2_20), .CLK(CK), .DIN(WX10355) );
  dffs1 \DFF_1523/Q_reg  ( .Q(CRC_OUT_2_19), .CLK(CK), .DIN(WX10353) );
  dffs1 \DFF_1522/Q_reg  ( .Q(CRC_OUT_2_18), .CLK(CK), .DIN(WX10351) );
  dffs1 \DFF_1521/Q_reg  ( .Q(CRC_OUT_2_17), .CLK(CK), .DIN(WX10349) );
  dffs1 \DFF_1520/Q_reg  ( .Q(CRC_OUT_2_16), .CLK(CK), .DIN(WX10347) );
  dffs1 \DFF_1519/Q_reg  ( .Q(CRC_OUT_2_15), .CLK(CK), .DIN(WX10345) );
  dffs1 \DFF_1518/Q_reg  ( .Q(CRC_OUT_2_14), .CLK(CK), .DIN(WX10343) );
  dffs1 \DFF_1517/Q_reg  ( .Q(CRC_OUT_2_13), .CLK(CK), .DIN(WX10341) );
  dffs1 \DFF_1516/Q_reg  ( .Q(CRC_OUT_2_12), .CLK(CK), .DIN(WX10339) );
  dffs1 \DFF_1515/Q_reg  ( .Q(CRC_OUT_2_11), .CLK(CK), .DIN(WX10337) );
  dffs1 \DFF_1514/Q_reg  ( .Q(CRC_OUT_2_10), .CLK(CK), .DIN(WX10335) );
  dffs1 \DFF_1513/Q_reg  ( .Q(CRC_OUT_2_9), .CLK(CK), .DIN(WX10333) );
  dffs1 \DFF_1512/Q_reg  ( .Q(CRC_OUT_2_8), .CLK(CK), .DIN(WX10331) );
  dffs1 \DFF_1511/Q_reg  ( .Q(CRC_OUT_2_7), .CLK(CK), .DIN(WX10329) );
  dffs1 \DFF_1510/Q_reg  ( .Q(CRC_OUT_2_6), .CLK(CK), .DIN(WX10327) );
  dffs1 \DFF_1509/Q_reg  ( .Q(CRC_OUT_2_5), .CLK(CK), .DIN(WX10325) );
  dffs1 \DFF_1508/Q_reg  ( .Q(CRC_OUT_2_4), .CLK(CK), .DIN(WX10323) );
  dffs1 \DFF_1507/Q_reg  ( .Q(CRC_OUT_2_3), .CLK(CK), .DIN(WX10321) );
  dffs1 \DFF_1506/Q_reg  ( .Q(CRC_OUT_2_2), .CLK(CK), .DIN(WX10319) );
  dffs1 \DFF_1505/Q_reg  ( .Q(CRC_OUT_2_1), .CLK(CK), .DIN(WX10317) );
  dffs1 \DFF_1504/Q_reg  ( .Q(CRC_OUT_2_0), .CLK(CK), .DIN(WX10315) );
  dffs1 \DFF_1503/Q_reg  ( .QN(n3205), .Q(WX9950), .CLK(CK), .DIN(WX9949) );
  dffs1 \DFF_1502/Q_reg  ( .QN(n3206), .Q(WX9948), .CLK(CK), .DIN(WX9947) );
  dffs1 \DFF_1501/Q_reg  ( .QN(n3207), .Q(WX9946), .CLK(CK), .DIN(WX9945) );
  dffs1 \DFF_1500/Q_reg  ( .QN(n3208), .Q(WX9944), .CLK(CK), .DIN(WX9943) );
  dffs1 \DFF_1499/Q_reg  ( .QN(n3209), .Q(WX9942), .CLK(CK), .DIN(WX9941) );
  dffs1 \DFF_1498/Q_reg  ( .QN(n3210), .Q(WX9940), .CLK(CK), .DIN(WX9939) );
  dffs1 \DFF_1497/Q_reg  ( .QN(n3211), .Q(WX9938), .CLK(CK), .DIN(WX9937) );
  dffs1 \DFF_1496/Q_reg  ( .QN(n3212), .Q(WX9936), .CLK(CK), .DIN(WX9935) );
  dffs1 \DFF_1495/Q_reg  ( .QN(n3213), .Q(WX9934), .CLK(CK), .DIN(WX9933) );
  dffs1 \DFF_1494/Q_reg  ( .QN(n3214), .Q(WX9932), .CLK(CK), .DIN(WX9931) );
  dffs1 \DFF_1493/Q_reg  ( .QN(n3215), .Q(WX9930), .CLK(CK), .DIN(WX9929) );
  dffs1 \DFF_1492/Q_reg  ( .QN(n3216), .Q(WX9928), .CLK(CK), .DIN(WX9927) );
  dffs1 \DFF_1491/Q_reg  ( .QN(n3217), .Q(WX9926), .CLK(CK), .DIN(WX9925) );
  dffs1 \DFF_1490/Q_reg  ( .QN(n3218), .Q(WX9924), .CLK(CK), .DIN(WX9923) );
  dffs1 \DFF_1489/Q_reg  ( .QN(n3219), .Q(WX9922), .CLK(CK), .DIN(WX9921) );
  dffs1 \DFF_1488/Q_reg  ( .QN(n3220), .Q(WX9920), .CLK(CK), .DIN(WX9919) );
  dffs1 \DFF_1487/Q_reg  ( .Q(WX9918), .CLK(CK), .DIN(WX9917) );
  dffs1 \DFF_1486/Q_reg  ( .Q(WX9916), .CLK(CK), .DIN(WX9915) );
  dffs1 \DFF_1485/Q_reg  ( .Q(WX9914), .CLK(CK), .DIN(WX9913) );
  dffs1 \DFF_1484/Q_reg  ( .Q(WX9912), .CLK(CK), .DIN(WX9911) );
  dffs1 \DFF_1483/Q_reg  ( .Q(WX9910), .CLK(CK), .DIN(WX9909) );
  dffs1 \DFF_1482/Q_reg  ( .Q(WX9908), .CLK(CK), .DIN(WX9907) );
  dffs1 \DFF_1481/Q_reg  ( .Q(WX9906), .CLK(CK), .DIN(WX9905) );
  dffs1 \DFF_1480/Q_reg  ( .Q(WX9904), .CLK(CK), .DIN(WX9903) );
  dffs1 \DFF_1479/Q_reg  ( .Q(WX9902), .CLK(CK), .DIN(WX9901) );
  dffs1 \DFF_1478/Q_reg  ( .Q(WX9900), .CLK(CK), .DIN(WX9899) );
  dffs1 \DFF_1477/Q_reg  ( .Q(WX9898), .CLK(CK), .DIN(WX9897) );
  dffs1 \DFF_1476/Q_reg  ( .Q(WX9896), .CLK(CK), .DIN(WX9895) );
  dffs1 \DFF_1475/Q_reg  ( .Q(WX9894), .CLK(CK), .DIN(WX9893) );
  dffs1 \DFF_1474/Q_reg  ( .Q(WX9892), .CLK(CK), .DIN(WX9891) );
  dffs1 \DFF_1473/Q_reg  ( .Q(WX9890), .CLK(CK), .DIN(WX9889) );
  dffs1 \DFF_1472/Q_reg  ( .Q(WX9888), .CLK(CK), .DIN(WX9887) );
  dffs1 \DFF_1471/Q_reg  ( .Q(WX9886), .CLK(CK), .DIN(WX9885) );
  dffs1 \DFF_1470/Q_reg  ( .Q(WX9884), .CLK(CK), .DIN(WX9883) );
  dffs1 \DFF_1469/Q_reg  ( .Q(WX9882), .CLK(CK), .DIN(WX9881) );
  dffs1 \DFF_1468/Q_reg  ( .Q(WX9880), .CLK(CK), .DIN(WX9879) );
  dffs1 \DFF_1467/Q_reg  ( .Q(WX9878), .CLK(CK), .DIN(WX9877) );
  dffs1 \DFF_1466/Q_reg  ( .Q(WX9876), .CLK(CK), .DIN(WX9875) );
  dffs1 \DFF_1465/Q_reg  ( .Q(WX9874), .CLK(CK), .DIN(WX9873) );
  dffs1 \DFF_1464/Q_reg  ( .Q(WX9872), .CLK(CK), .DIN(WX9871) );
  dffs1 \DFF_1463/Q_reg  ( .Q(WX9870), .CLK(CK), .DIN(WX9869) );
  dffs1 \DFF_1462/Q_reg  ( .Q(WX9868), .CLK(CK), .DIN(WX9867) );
  dffs1 \DFF_1461/Q_reg  ( .Q(WX9866), .CLK(CK), .DIN(WX9865) );
  dffs1 \DFF_1460/Q_reg  ( .Q(WX9864), .CLK(CK), .DIN(WX9863) );
  dffs1 \DFF_1459/Q_reg  ( .Q(WX9862), .CLK(CK), .DIN(WX9861) );
  dffs1 \DFF_1458/Q_reg  ( .Q(WX9860), .CLK(CK), .DIN(WX9859) );
  dffs1 \DFF_1457/Q_reg  ( .Q(WX9858), .CLK(CK), .DIN(WX9857) );
  dffs1 \DFF_1456/Q_reg  ( .Q(WX9856), .CLK(CK), .DIN(WX9855) );
  dffs1 \DFF_1455/Q_reg  ( .Q(WX9854), .CLK(CK), .DIN(WX9853) );
  dffs1 \DFF_1454/Q_reg  ( .Q(WX9852), .CLK(CK), .DIN(WX9851) );
  dffs1 \DFF_1453/Q_reg  ( .Q(WX9850), .CLK(CK), .DIN(WX9849) );
  dffs1 \DFF_1452/Q_reg  ( .Q(WX9848), .CLK(CK), .DIN(WX9847) );
  dffs1 \DFF_1451/Q_reg  ( .Q(WX9846), .CLK(CK), .DIN(WX9845) );
  dffs1 \DFF_1450/Q_reg  ( .Q(WX9844), .CLK(CK), .DIN(WX9843) );
  dffs1 \DFF_1449/Q_reg  ( .Q(WX9842), .CLK(CK), .DIN(WX9841) );
  dffs1 \DFF_1448/Q_reg  ( .Q(WX9840), .CLK(CK), .DIN(WX9839) );
  dffs1 \DFF_1447/Q_reg  ( .Q(WX9838), .CLK(CK), .DIN(WX9837) );
  dffs1 \DFF_1446/Q_reg  ( .Q(WX9836), .CLK(CK), .DIN(WX9835) );
  dffs1 \DFF_1445/Q_reg  ( .Q(WX9834), .CLK(CK), .DIN(WX9833) );
  dffs1 \DFF_1444/Q_reg  ( .Q(WX9832), .CLK(CK), .DIN(WX9831) );
  dffs1 \DFF_1443/Q_reg  ( .Q(WX9830), .CLK(CK), .DIN(WX9829) );
  dffs1 \DFF_1442/Q_reg  ( .Q(WX9828), .CLK(CK), .DIN(WX9827) );
  dffs1 \DFF_1441/Q_reg  ( .Q(WX9826), .CLK(CK), .DIN(WX9825) );
  dffs1 \DFF_1440/Q_reg  ( .Q(WX9824), .CLK(CK), .DIN(WX9823) );
  dffs1 \DFF_1439/Q_reg  ( .Q(WX9822), .CLK(CK), .DIN(WX9821) );
  dffs1 \DFF_1438/Q_reg  ( .Q(WX9820), .CLK(CK), .DIN(WX9819) );
  dffs1 \DFF_1437/Q_reg  ( .Q(WX9818), .CLK(CK), .DIN(WX9817) );
  dffs1 \DFF_1436/Q_reg  ( .Q(WX9816), .CLK(CK), .DIN(WX9815) );
  dffs1 \DFF_1435/Q_reg  ( .Q(WX9814), .CLK(CK), .DIN(WX9813) );
  dffs1 \DFF_1434/Q_reg  ( .Q(WX9812), .CLK(CK), .DIN(WX9811) );
  dffs1 \DFF_1433/Q_reg  ( .Q(WX9810), .CLK(CK), .DIN(WX9809) );
  dffs1 \DFF_1432/Q_reg  ( .Q(WX9808), .CLK(CK), .DIN(WX9807) );
  dffs1 \DFF_1431/Q_reg  ( .Q(WX9806), .CLK(CK), .DIN(WX9805) );
  dffs1 \DFF_1430/Q_reg  ( .Q(WX9804), .CLK(CK), .DIN(WX9803) );
  dffs1 \DFF_1429/Q_reg  ( .Q(WX9802), .CLK(CK), .DIN(WX9801) );
  dffs1 \DFF_1428/Q_reg  ( .Q(WX9800), .CLK(CK), .DIN(WX9799) );
  dffs1 \DFF_1427/Q_reg  ( .Q(WX9798), .CLK(CK), .DIN(WX9797) );
  dffs1 \DFF_1426/Q_reg  ( .Q(WX9796), .CLK(CK), .DIN(WX9795) );
  dffs1 \DFF_1425/Q_reg  ( .Q(WX9794), .CLK(CK), .DIN(WX9793) );
  dffs1 \DFF_1424/Q_reg  ( .Q(WX9792), .CLK(CK), .DIN(WX9791) );
  dffs1 \DFF_1423/Q_reg  ( .QN(n2949), .CLK(CK), .DIN(WX9789) );
  dffs1 \DFF_1422/Q_reg  ( .QN(n2950), .CLK(CK), .DIN(WX9787) );
  dffs1 \DFF_1421/Q_reg  ( .QN(n2951), .CLK(CK), .DIN(WX9785) );
  dffs1 \DFF_1420/Q_reg  ( .QN(n2952), .CLK(CK), .DIN(WX9783) );
  dffs1 \DFF_1419/Q_reg  ( .QN(n2953), .CLK(CK), .DIN(WX9781) );
  dffs1 \DFF_1418/Q_reg  ( .QN(n2954), .CLK(CK), .DIN(WX9779) );
  dffs1 \DFF_1417/Q_reg  ( .QN(n2955), .CLK(CK), .DIN(WX9777) );
  dffs1 \DFF_1416/Q_reg  ( .QN(n2956), .CLK(CK), .DIN(WX9775) );
  dffs1 \DFF_1415/Q_reg  ( .QN(n2957), .CLK(CK), .DIN(WX9773) );
  dffs1 \DFF_1414/Q_reg  ( .QN(n2958), .CLK(CK), .DIN(WX9771) );
  dffs1 \DFF_1413/Q_reg  ( .QN(n2959), .CLK(CK), .DIN(WX9769) );
  dffs1 \DFF_1412/Q_reg  ( .QN(n2960), .CLK(CK), .DIN(WX9767) );
  dffs1 \DFF_1411/Q_reg  ( .QN(n2961), .CLK(CK), .DIN(WX9765) );
  dffs1 \DFF_1410/Q_reg  ( .QN(n2962), .CLK(CK), .DIN(WX9763) );
  dffs1 \DFF_1409/Q_reg  ( .QN(n2963), .CLK(CK), .DIN(WX9761) );
  dffs1 \DFF_1408/Q_reg  ( .QN(n2964), .CLK(CK), .DIN(WX9759) );
  dffs1 \DFF_1407/Q_reg  ( .QN(n3109), .CLK(CK), .DIN(WX9757) );
  dffs1 \DFF_1406/Q_reg  ( .QN(n3110), .CLK(CK), .DIN(WX9755) );
  dffs1 \DFF_1405/Q_reg  ( .QN(n3111), .CLK(CK), .DIN(WX9753) );
  dffs1 \DFF_1404/Q_reg  ( .QN(n3112), .CLK(CK), .DIN(WX9751) );
  dffs1 \DFF_1403/Q_reg  ( .QN(n3113), .CLK(CK), .DIN(WX9749) );
  dffs1 \DFF_1402/Q_reg  ( .QN(n3114), .CLK(CK), .DIN(WX9747) );
  dffs1 \DFF_1401/Q_reg  ( .QN(n3115), .CLK(CK), .DIN(WX9745) );
  dffs1 \DFF_1400/Q_reg  ( .QN(n3116), .CLK(CK), .DIN(WX9743) );
  dffs1 \DFF_1399/Q_reg  ( .QN(n3117), .CLK(CK), .DIN(WX9741) );
  dffs1 \DFF_1398/Q_reg  ( .QN(n3118), .CLK(CK), .DIN(WX9739) );
  dffs1 \DFF_1397/Q_reg  ( .QN(n3119), .CLK(CK), .DIN(WX9737) );
  dffs1 \DFF_1396/Q_reg  ( .QN(n3120), .CLK(CK), .DIN(WX9735) );
  dffs1 \DFF_1395/Q_reg  ( .QN(n3121), .CLK(CK), .DIN(WX9733) );
  dffs1 \DFF_1394/Q_reg  ( .QN(n3122), .CLK(CK), .DIN(WX9731) );
  dffs1 \DFF_1393/Q_reg  ( .QN(n3123), .CLK(CK), .DIN(WX9729) );
  dffs1 \DFF_1392/Q_reg  ( .QN(n3124), .CLK(CK), .DIN(WX9727) );
  dffs1 \DFF_1391/Q_reg  ( .Q(WX9726), .CLK(CK), .DIN(WX9725) );
  dffs1 \DFF_1390/Q_reg  ( .Q(WX9724), .CLK(CK), .DIN(WX9723) );
  dffs1 \DFF_1389/Q_reg  ( .Q(WX9722), .CLK(CK), .DIN(WX9721) );
  dffs1 \DFF_1388/Q_reg  ( .Q(WX9720), .CLK(CK), .DIN(WX9719) );
  dffs1 \DFF_1387/Q_reg  ( .Q(WX9718), .CLK(CK), .DIN(WX9717) );
  dffs1 \DFF_1386/Q_reg  ( .Q(WX9716), .CLK(CK), .DIN(WX9715) );
  dffs1 \DFF_1385/Q_reg  ( .Q(WX9714), .CLK(CK), .DIN(WX9713) );
  dffs1 \DFF_1384/Q_reg  ( .Q(WX9712), .CLK(CK), .DIN(WX9711) );
  dffs1 \DFF_1383/Q_reg  ( .Q(WX9710), .CLK(CK), .DIN(WX9709) );
  dffs1 \DFF_1382/Q_reg  ( .Q(WX9708), .CLK(CK), .DIN(WX9707) );
  dffs1 \DFF_1381/Q_reg  ( .Q(WX9706), .CLK(CK), .DIN(WX9705) );
  dffs1 \DFF_1380/Q_reg  ( .Q(WX9704), .CLK(CK), .DIN(WX9703) );
  dffs1 \DFF_1379/Q_reg  ( .Q(WX9702), .CLK(CK), .DIN(WX9701) );
  dffs1 \DFF_1378/Q_reg  ( .Q(WX9700), .CLK(CK), .DIN(WX9699) );
  dffs1 \DFF_1377/Q_reg  ( .Q(WX9698), .CLK(CK), .DIN(WX9697) );
  dffs1 \DFF_1376/Q_reg  ( .Q(WX9696), .CLK(CK), .DIN(WX9695) );
  dffs1 \DFF_1375/Q_reg  ( .Q(WX9598), .CLK(CK), .DIN(WX9597) );
  dffs1 \DFF_1374/Q_reg  ( .Q(WX9596), .CLK(CK), .DIN(WX9595) );
  dffs1 \DFF_1373/Q_reg  ( .Q(WX9594), .CLK(CK), .DIN(WX9593) );
  dffs1 \DFF_1372/Q_reg  ( .Q(WX9592), .CLK(CK), .DIN(WX9591) );
  dffs1 \DFF_1371/Q_reg  ( .Q(WX9590), .CLK(CK), .DIN(WX9589) );
  dffs1 \DFF_1370/Q_reg  ( .Q(WX9588), .CLK(CK), .DIN(WX9587) );
  dffs1 \DFF_1369/Q_reg  ( .Q(WX9586), .CLK(CK), .DIN(WX9585) );
  dffs1 \DFF_1368/Q_reg  ( .Q(WX9584), .CLK(CK), .DIN(WX9583) );
  dffs1 \DFF_1367/Q_reg  ( .Q(WX9582), .CLK(CK), .DIN(WX9581) );
  dffs1 \DFF_1366/Q_reg  ( .Q(WX9580), .CLK(CK), .DIN(WX9579) );
  dffs1 \DFF_1365/Q_reg  ( .Q(WX9578), .CLK(CK), .DIN(WX9577) );
  dffs1 \DFF_1364/Q_reg  ( .Q(WX9576), .CLK(CK), .DIN(WX9575) );
  dffs1 \DFF_1363/Q_reg  ( .Q(WX9574), .CLK(CK), .DIN(WX9573) );
  dffs1 \DFF_1362/Q_reg  ( .Q(WX9572), .CLK(CK), .DIN(WX9571) );
  dffs1 \DFF_1361/Q_reg  ( .Q(WX9570), .CLK(CK), .DIN(WX9569) );
  dffs1 \DFF_1360/Q_reg  ( .Q(WX9568), .CLK(CK), .DIN(WX9567) );
  dffs1 \DFF_1359/Q_reg  ( .Q(WX9566), .CLK(CK), .DIN(WX9565) );
  dffs1 \DFF_1358/Q_reg  ( .Q(WX9564), .CLK(CK), .DIN(WX9563) );
  dffs1 \DFF_1357/Q_reg  ( .Q(WX9562), .CLK(CK), .DIN(WX9561) );
  dffs1 \DFF_1356/Q_reg  ( .Q(WX9560), .CLK(CK), .DIN(WX9559) );
  dffs1 \DFF_1355/Q_reg  ( .Q(WX9558), .CLK(CK), .DIN(WX9557) );
  dffs1 \DFF_1354/Q_reg  ( .Q(WX9556), .CLK(CK), .DIN(WX9555) );
  dffs1 \DFF_1353/Q_reg  ( .Q(WX9554), .CLK(CK), .DIN(WX9553) );
  dffs1 \DFF_1352/Q_reg  ( .Q(WX9552), .CLK(CK), .DIN(WX9551) );
  dffs1 \DFF_1351/Q_reg  ( .Q(WX9550), .CLK(CK), .DIN(WX9549) );
  dffs1 \DFF_1350/Q_reg  ( .Q(WX9548), .CLK(CK), .DIN(WX9547) );
  dffs1 \DFF_1349/Q_reg  ( .Q(WX9546), .CLK(CK), .DIN(WX9545) );
  dffs1 \DFF_1348/Q_reg  ( .Q(WX9544), .CLK(CK), .DIN(WX9543) );
  dffs1 \DFF_1347/Q_reg  ( .Q(WX9542), .CLK(CK), .DIN(WX9541) );
  dffs1 \DFF_1346/Q_reg  ( .Q(WX9540), .CLK(CK), .DIN(WX9539) );
  dffs1 \DFF_1345/Q_reg  ( .Q(WX9538), .CLK(CK), .DIN(WX9537) );
  dffs1 \DFF_1344/Q_reg  ( .Q(WX9536), .CLK(CK), .DIN(WX9535) );
  dffs1 \DFF_1343/Q_reg  ( .Q(CRC_OUT_3_31), .CLK(CK), .DIN(WX9084) );
  dffs1 \DFF_1342/Q_reg  ( .Q(CRC_OUT_3_30), .CLK(CK), .DIN(WX9082) );
  dffs1 \DFF_1341/Q_reg  ( .Q(CRC_OUT_3_29), .CLK(CK), .DIN(WX9080) );
  dffs1 \DFF_1340/Q_reg  ( .Q(CRC_OUT_3_28), .CLK(CK), .DIN(WX9078) );
  dffs1 \DFF_1339/Q_reg  ( .Q(CRC_OUT_3_27), .CLK(CK), .DIN(WX9076) );
  dffs1 \DFF_1338/Q_reg  ( .Q(CRC_OUT_3_26), .CLK(CK), .DIN(WX9074) );
  dffs1 \DFF_1337/Q_reg  ( .Q(CRC_OUT_3_25), .CLK(CK), .DIN(WX9072) );
  dffs1 \DFF_1336/Q_reg  ( .Q(CRC_OUT_3_24), .CLK(CK), .DIN(WX9070) );
  dffs1 \DFF_1335/Q_reg  ( .Q(CRC_OUT_3_23), .CLK(CK), .DIN(WX9068) );
  dffs1 \DFF_1334/Q_reg  ( .Q(CRC_OUT_3_22), .CLK(CK), .DIN(WX9066) );
  dffs1 \DFF_1333/Q_reg  ( .Q(CRC_OUT_3_21), .CLK(CK), .DIN(WX9064) );
  dffs1 \DFF_1332/Q_reg  ( .Q(CRC_OUT_3_20), .CLK(CK), .DIN(WX9062) );
  dffs1 \DFF_1331/Q_reg  ( .Q(CRC_OUT_3_19), .CLK(CK), .DIN(WX9060) );
  dffs1 \DFF_1330/Q_reg  ( .Q(CRC_OUT_3_18), .CLK(CK), .DIN(WX9058) );
  dffs1 \DFF_1329/Q_reg  ( .Q(CRC_OUT_3_17), .CLK(CK), .DIN(WX9056) );
  dffs1 \DFF_1328/Q_reg  ( .Q(CRC_OUT_3_16), .CLK(CK), .DIN(WX9054) );
  dffs1 \DFF_1327/Q_reg  ( .Q(CRC_OUT_3_15), .CLK(CK), .DIN(WX9052) );
  dffs1 \DFF_1326/Q_reg  ( .Q(CRC_OUT_3_14), .CLK(CK), .DIN(WX9050) );
  dffs1 \DFF_1325/Q_reg  ( .Q(CRC_OUT_3_13), .CLK(CK), .DIN(WX9048) );
  dffs1 \DFF_1324/Q_reg  ( .Q(CRC_OUT_3_12), .CLK(CK), .DIN(WX9046) );
  dffs1 \DFF_1323/Q_reg  ( .Q(CRC_OUT_3_11), .CLK(CK), .DIN(WX9044) );
  dffs1 \DFF_1322/Q_reg  ( .Q(CRC_OUT_3_10), .CLK(CK), .DIN(WX9042) );
  dffs1 \DFF_1321/Q_reg  ( .Q(CRC_OUT_3_9), .CLK(CK), .DIN(WX9040) );
  dffs1 \DFF_1320/Q_reg  ( .Q(CRC_OUT_3_8), .CLK(CK), .DIN(WX9038) );
  dffs1 \DFF_1319/Q_reg  ( .Q(CRC_OUT_3_7), .CLK(CK), .DIN(WX9036) );
  dffs1 \DFF_1318/Q_reg  ( .Q(CRC_OUT_3_6), .CLK(CK), .DIN(WX9034) );
  dffs1 \DFF_1317/Q_reg  ( .Q(CRC_OUT_3_5), .CLK(CK), .DIN(WX9032) );
  dffs1 \DFF_1316/Q_reg  ( .Q(CRC_OUT_3_4), .CLK(CK), .DIN(WX9030) );
  dffs1 \DFF_1315/Q_reg  ( .Q(CRC_OUT_3_3), .CLK(CK), .DIN(WX9028) );
  dffs1 \DFF_1314/Q_reg  ( .Q(CRC_OUT_3_2), .CLK(CK), .DIN(WX9026) );
  dffs1 \DFF_1313/Q_reg  ( .Q(CRC_OUT_3_1), .CLK(CK), .DIN(WX9024) );
  dffs1 \DFF_1312/Q_reg  ( .Q(CRC_OUT_3_0), .CLK(CK), .DIN(WX9022) );
  dffs1 \DFF_1311/Q_reg  ( .QN(n3221), .Q(WX8657), .CLK(CK), .DIN(WX8656) );
  dffs1 \DFF_1310/Q_reg  ( .QN(n3222), .Q(WX8655), .CLK(CK), .DIN(WX8654) );
  dffs1 \DFF_1309/Q_reg  ( .QN(n3223), .Q(WX8653), .CLK(CK), .DIN(WX8652) );
  dffs1 \DFF_1308/Q_reg  ( .QN(n3224), .Q(WX8651), .CLK(CK), .DIN(WX8650) );
  dffs1 \DFF_1307/Q_reg  ( .QN(n3225), .Q(WX8649), .CLK(CK), .DIN(WX8648) );
  dffs1 \DFF_1306/Q_reg  ( .QN(n3226), .Q(WX8647), .CLK(CK), .DIN(WX8646) );
  dffs1 \DFF_1305/Q_reg  ( .QN(n3227), .Q(WX8645), .CLK(CK), .DIN(WX8644) );
  dffs1 \DFF_1304/Q_reg  ( .QN(n3228), .Q(WX8643), .CLK(CK), .DIN(WX8642) );
  dffs1 \DFF_1303/Q_reg  ( .QN(n3229), .Q(WX8641), .CLK(CK), .DIN(WX8640) );
  dffs1 \DFF_1302/Q_reg  ( .QN(n3230), .Q(WX8639), .CLK(CK), .DIN(WX8638) );
  dffs1 \DFF_1301/Q_reg  ( .QN(n3231), .Q(WX8637), .CLK(CK), .DIN(WX8636) );
  dffs1 \DFF_1300/Q_reg  ( .QN(n3232), .Q(WX8635), .CLK(CK), .DIN(WX8634) );
  dffs1 \DFF_1299/Q_reg  ( .QN(n3233), .Q(WX8633), .CLK(CK), .DIN(WX8632) );
  dffs1 \DFF_1298/Q_reg  ( .QN(n3234), .Q(WX8631), .CLK(CK), .DIN(WX8630) );
  dffs1 \DFF_1297/Q_reg  ( .QN(n3235), .Q(WX8629), .CLK(CK), .DIN(WX8628) );
  dffs1 \DFF_1296/Q_reg  ( .QN(n3236), .Q(WX8627), .CLK(CK), .DIN(WX8626) );
  dffs1 \DFF_1295/Q_reg  ( .Q(WX8625), .CLK(CK), .DIN(WX8624) );
  dffs1 \DFF_1294/Q_reg  ( .Q(WX8623), .CLK(CK), .DIN(WX8622) );
  dffs1 \DFF_1293/Q_reg  ( .Q(WX8621), .CLK(CK), .DIN(WX8620) );
  dffs1 \DFF_1292/Q_reg  ( .Q(WX8619), .CLK(CK), .DIN(WX8618) );
  dffs1 \DFF_1291/Q_reg  ( .Q(WX8617), .CLK(CK), .DIN(WX8616) );
  dffs1 \DFF_1290/Q_reg  ( .Q(WX8615), .CLK(CK), .DIN(WX8614) );
  dffs1 \DFF_1289/Q_reg  ( .Q(WX8613), .CLK(CK), .DIN(WX8612) );
  dffs1 \DFF_1288/Q_reg  ( .Q(WX8611), .CLK(CK), .DIN(WX8610) );
  dffs1 \DFF_1287/Q_reg  ( .Q(WX8609), .CLK(CK), .DIN(WX8608) );
  dffs1 \DFF_1286/Q_reg  ( .Q(WX8607), .CLK(CK), .DIN(WX8606) );
  dffs1 \DFF_1285/Q_reg  ( .Q(WX8605), .CLK(CK), .DIN(WX8604) );
  dffs1 \DFF_1284/Q_reg  ( .Q(WX8603), .CLK(CK), .DIN(WX8602) );
  dffs1 \DFF_1283/Q_reg  ( .Q(WX8601), .CLK(CK), .DIN(WX8600) );
  dffs1 \DFF_1282/Q_reg  ( .Q(WX8599), .CLK(CK), .DIN(WX8598) );
  dffs1 \DFF_1281/Q_reg  ( .Q(WX8597), .CLK(CK), .DIN(WX8596) );
  dffs1 \DFF_1280/Q_reg  ( .Q(WX8595), .CLK(CK), .DIN(WX8594) );
  dffs1 \DFF_1279/Q_reg  ( .Q(WX8593), .CLK(CK), .DIN(WX8592) );
  dffs1 \DFF_1278/Q_reg  ( .Q(WX8591), .CLK(CK), .DIN(WX8590) );
  dffs1 \DFF_1277/Q_reg  ( .Q(WX8589), .CLK(CK), .DIN(WX8588) );
  dffs1 \DFF_1276/Q_reg  ( .Q(WX8587), .CLK(CK), .DIN(WX8586) );
  dffs1 \DFF_1275/Q_reg  ( .Q(WX8585), .CLK(CK), .DIN(WX8584) );
  dffs1 \DFF_1274/Q_reg  ( .Q(WX8583), .CLK(CK), .DIN(WX8582) );
  dffs1 \DFF_1273/Q_reg  ( .Q(WX8581), .CLK(CK), .DIN(WX8580) );
  dffs1 \DFF_1272/Q_reg  ( .Q(WX8579), .CLK(CK), .DIN(WX8578) );
  dffs1 \DFF_1271/Q_reg  ( .Q(WX8577), .CLK(CK), .DIN(WX8576) );
  dffs1 \DFF_1270/Q_reg  ( .Q(WX8575), .CLK(CK), .DIN(WX8574) );
  dffs1 \DFF_1269/Q_reg  ( .Q(WX8573), .CLK(CK), .DIN(WX8572) );
  dffs1 \DFF_1268/Q_reg  ( .Q(WX8571), .CLK(CK), .DIN(WX8570) );
  dffs1 \DFF_1267/Q_reg  ( .Q(WX8569), .CLK(CK), .DIN(WX8568) );
  dffs1 \DFF_1266/Q_reg  ( .Q(WX8567), .CLK(CK), .DIN(WX8566) );
  dffs1 \DFF_1265/Q_reg  ( .Q(WX8565), .CLK(CK), .DIN(WX8564) );
  dffs1 \DFF_1264/Q_reg  ( .Q(WX8563), .CLK(CK), .DIN(WX8562) );
  dffs1 \DFF_1263/Q_reg  ( .Q(WX8561), .CLK(CK), .DIN(WX8560) );
  dffs1 \DFF_1262/Q_reg  ( .Q(WX8559), .CLK(CK), .DIN(WX8558) );
  dffs1 \DFF_1261/Q_reg  ( .Q(WX8557), .CLK(CK), .DIN(WX8556) );
  dffs1 \DFF_1260/Q_reg  ( .Q(WX8555), .CLK(CK), .DIN(WX8554) );
  dffs1 \DFF_1259/Q_reg  ( .Q(WX8553), .CLK(CK), .DIN(WX8552) );
  dffs1 \DFF_1258/Q_reg  ( .Q(WX8551), .CLK(CK), .DIN(WX8550) );
  dffs1 \DFF_1257/Q_reg  ( .Q(WX8549), .CLK(CK), .DIN(WX8548) );
  dffs1 \DFF_1256/Q_reg  ( .Q(WX8547), .CLK(CK), .DIN(WX8546) );
  dffs1 \DFF_1255/Q_reg  ( .Q(WX8545), .CLK(CK), .DIN(WX8544) );
  dffs1 \DFF_1254/Q_reg  ( .Q(WX8543), .CLK(CK), .DIN(WX8542) );
  dffs1 \DFF_1253/Q_reg  ( .Q(WX8541), .CLK(CK), .DIN(WX8540) );
  dffs1 \DFF_1252/Q_reg  ( .Q(WX8539), .CLK(CK), .DIN(WX8538) );
  dffs1 \DFF_1251/Q_reg  ( .Q(WX8537), .CLK(CK), .DIN(WX8536) );
  dffs1 \DFF_1250/Q_reg  ( .Q(WX8535), .CLK(CK), .DIN(WX8534) );
  dffs1 \DFF_1249/Q_reg  ( .Q(WX8533), .CLK(CK), .DIN(WX8532) );
  dffs1 \DFF_1248/Q_reg  ( .Q(WX8531), .CLK(CK), .DIN(WX8530) );
  dffs1 \DFF_1247/Q_reg  ( .Q(WX8529), .CLK(CK), .DIN(WX8528) );
  dffs1 \DFF_1246/Q_reg  ( .Q(WX8527), .CLK(CK), .DIN(WX8526) );
  dffs1 \DFF_1245/Q_reg  ( .Q(WX8525), .CLK(CK), .DIN(WX8524) );
  dffs1 \DFF_1244/Q_reg  ( .Q(WX8523), .CLK(CK), .DIN(WX8522) );
  dffs1 \DFF_1243/Q_reg  ( .Q(WX8521), .CLK(CK), .DIN(WX8520) );
  dffs1 \DFF_1242/Q_reg  ( .Q(WX8519), .CLK(CK), .DIN(WX8518) );
  dffs1 \DFF_1241/Q_reg  ( .Q(WX8517), .CLK(CK), .DIN(WX8516) );
  dffs1 \DFF_1240/Q_reg  ( .Q(WX8515), .CLK(CK), .DIN(WX8514) );
  dffs1 \DFF_1239/Q_reg  ( .Q(WX8513), .CLK(CK), .DIN(WX8512) );
  dffs1 \DFF_1238/Q_reg  ( .Q(WX8511), .CLK(CK), .DIN(WX8510) );
  dffs1 \DFF_1237/Q_reg  ( .Q(WX8509), .CLK(CK), .DIN(WX8508) );
  dffs1 \DFF_1236/Q_reg  ( .Q(WX8507), .CLK(CK), .DIN(WX8506) );
  dffs1 \DFF_1235/Q_reg  ( .Q(WX8505), .CLK(CK), .DIN(WX8504) );
  dffs1 \DFF_1234/Q_reg  ( .Q(WX8503), .CLK(CK), .DIN(WX8502) );
  dffs1 \DFF_1233/Q_reg  ( .Q(WX8501), .CLK(CK), .DIN(WX8500) );
  dffs1 \DFF_1232/Q_reg  ( .Q(WX8499), .CLK(CK), .DIN(WX8498) );
  dffs1 \DFF_1231/Q_reg  ( .QN(n2965), .CLK(CK), .DIN(WX8496) );
  dffs1 \DFF_1230/Q_reg  ( .QN(n2966), .CLK(CK), .DIN(WX8494) );
  dffs1 \DFF_1229/Q_reg  ( .QN(n2967), .CLK(CK), .DIN(WX8492) );
  dffs1 \DFF_1228/Q_reg  ( .QN(n2968), .CLK(CK), .DIN(WX8490) );
  dffs1 \DFF_1227/Q_reg  ( .QN(n2969), .CLK(CK), .DIN(WX8488) );
  dffs1 \DFF_1226/Q_reg  ( .QN(n2970), .CLK(CK), .DIN(WX8486) );
  dffs1 \DFF_1225/Q_reg  ( .QN(n2971), .CLK(CK), .DIN(WX8484) );
  dffs1 \DFF_1224/Q_reg  ( .QN(n2972), .CLK(CK), .DIN(WX8482) );
  dffs1 \DFF_1223/Q_reg  ( .QN(n2973), .CLK(CK), .DIN(WX8480) );
  dffs1 \DFF_1222/Q_reg  ( .QN(n2974), .CLK(CK), .DIN(WX8478) );
  dffs1 \DFF_1221/Q_reg  ( .QN(n2975), .CLK(CK), .DIN(WX8476) );
  dffs1 \DFF_1220/Q_reg  ( .QN(n2976), .CLK(CK), .DIN(WX8474) );
  dffs1 \DFF_1219/Q_reg  ( .QN(n2977), .CLK(CK), .DIN(WX8472) );
  dffs1 \DFF_1218/Q_reg  ( .QN(n2978), .CLK(CK), .DIN(WX8470) );
  dffs1 \DFF_1217/Q_reg  ( .QN(n2979), .CLK(CK), .DIN(WX8468) );
  dffs1 \DFF_1216/Q_reg  ( .QN(n2980), .CLK(CK), .DIN(WX8466) );
  dffs1 \DFF_1215/Q_reg  ( .QN(n3125), .CLK(CK), .DIN(WX8464) );
  dffs1 \DFF_1214/Q_reg  ( .QN(n3126), .CLK(CK), .DIN(WX8462) );
  dffs1 \DFF_1213/Q_reg  ( .QN(n3127), .CLK(CK), .DIN(WX8460) );
  dffs1 \DFF_1212/Q_reg  ( .QN(n3128), .CLK(CK), .DIN(WX8458) );
  dffs1 \DFF_1211/Q_reg  ( .QN(n3129), .CLK(CK), .DIN(WX8456) );
  dffs1 \DFF_1210/Q_reg  ( .QN(n3130), .CLK(CK), .DIN(WX8454) );
  dffs1 \DFF_1209/Q_reg  ( .QN(n3131), .CLK(CK), .DIN(WX8452) );
  dffs1 \DFF_1208/Q_reg  ( .QN(n3132), .CLK(CK), .DIN(WX8450) );
  dffs1 \DFF_1207/Q_reg  ( .QN(n3133), .CLK(CK), .DIN(WX8448) );
  dffs1 \DFF_1206/Q_reg  ( .QN(n3134), .CLK(CK), .DIN(WX8446) );
  dffs1 \DFF_1205/Q_reg  ( .QN(n3135), .CLK(CK), .DIN(WX8444) );
  dffs1 \DFF_1204/Q_reg  ( .QN(n3136), .CLK(CK), .DIN(WX8442) );
  dffs1 \DFF_1203/Q_reg  ( .QN(n3137), .CLK(CK), .DIN(WX8440) );
  dffs1 \DFF_1202/Q_reg  ( .QN(n3138), .CLK(CK), .DIN(WX8438) );
  dffs1 \DFF_1201/Q_reg  ( .QN(n3139), .CLK(CK), .DIN(WX8436) );
  dffs1 \DFF_1200/Q_reg  ( .QN(n3140), .CLK(CK), .DIN(WX8434) );
  dffs1 \DFF_1199/Q_reg  ( .Q(WX8433), .CLK(CK), .DIN(WX8432) );
  dffs1 \DFF_1198/Q_reg  ( .Q(WX8431), .CLK(CK), .DIN(WX8430) );
  dffs1 \DFF_1197/Q_reg  ( .Q(WX8429), .CLK(CK), .DIN(WX8428) );
  dffs1 \DFF_1196/Q_reg  ( .Q(WX8427), .CLK(CK), .DIN(WX8426) );
  dffs1 \DFF_1195/Q_reg  ( .Q(WX8425), .CLK(CK), .DIN(WX8424) );
  dffs1 \DFF_1194/Q_reg  ( .Q(WX8423), .CLK(CK), .DIN(WX8422) );
  dffs1 \DFF_1193/Q_reg  ( .Q(WX8421), .CLK(CK), .DIN(WX8420) );
  dffs1 \DFF_1192/Q_reg  ( .Q(WX8419), .CLK(CK), .DIN(WX8418) );
  dffs1 \DFF_1191/Q_reg  ( .Q(WX8417), .CLK(CK), .DIN(WX8416) );
  dffs1 \DFF_1190/Q_reg  ( .Q(WX8415), .CLK(CK), .DIN(WX8414) );
  dffs1 \DFF_1189/Q_reg  ( .Q(WX8413), .CLK(CK), .DIN(WX8412) );
  dffs1 \DFF_1188/Q_reg  ( .Q(WX8411), .CLK(CK), .DIN(WX8410) );
  dffs1 \DFF_1187/Q_reg  ( .Q(WX8409), .CLK(CK), .DIN(WX8408) );
  dffs1 \DFF_1186/Q_reg  ( .Q(WX8407), .CLK(CK), .DIN(WX8406) );
  dffs1 \DFF_1185/Q_reg  ( .Q(WX8405), .CLK(CK), .DIN(WX8404) );
  dffs1 \DFF_1184/Q_reg  ( .Q(WX8403), .CLK(CK), .DIN(WX8402) );
  dffs1 \DFF_1183/Q_reg  ( .Q(WX8305), .CLK(CK), .DIN(WX8304) );
  dffs1 \DFF_1182/Q_reg  ( .Q(WX8303), .CLK(CK), .DIN(WX8302) );
  dffs1 \DFF_1181/Q_reg  ( .Q(WX8301), .CLK(CK), .DIN(WX8300) );
  dffs1 \DFF_1180/Q_reg  ( .Q(WX8299), .CLK(CK), .DIN(WX8298) );
  dffs1 \DFF_1179/Q_reg  ( .Q(WX8297), .CLK(CK), .DIN(WX8296) );
  dffs1 \DFF_1178/Q_reg  ( .Q(WX8295), .CLK(CK), .DIN(WX8294) );
  dffs1 \DFF_1177/Q_reg  ( .Q(WX8293), .CLK(CK), .DIN(WX8292) );
  dffs1 \DFF_1176/Q_reg  ( .Q(WX8291), .CLK(CK), .DIN(WX8290) );
  dffs1 \DFF_1175/Q_reg  ( .Q(WX8289), .CLK(CK), .DIN(WX8288) );
  dffs1 \DFF_1174/Q_reg  ( .Q(WX8287), .CLK(CK), .DIN(WX8286) );
  dffs1 \DFF_1173/Q_reg  ( .Q(WX8285), .CLK(CK), .DIN(WX8284) );
  dffs1 \DFF_1172/Q_reg  ( .Q(WX8283), .CLK(CK), .DIN(WX8282) );
  dffs1 \DFF_1171/Q_reg  ( .Q(WX8281), .CLK(CK), .DIN(WX8280) );
  dffs1 \DFF_1170/Q_reg  ( .Q(WX8279), .CLK(CK), .DIN(WX8278) );
  dffs1 \DFF_1169/Q_reg  ( .Q(WX8277), .CLK(CK), .DIN(WX8276) );
  dffs1 \DFF_1168/Q_reg  ( .Q(WX8275), .CLK(CK), .DIN(WX8274) );
  dffs1 \DFF_1167/Q_reg  ( .Q(WX8273), .CLK(CK), .DIN(WX8272) );
  dffs1 \DFF_1166/Q_reg  ( .Q(WX8271), .CLK(CK), .DIN(WX8270) );
  dffs1 \DFF_1165/Q_reg  ( .Q(WX8269), .CLK(CK), .DIN(WX8268) );
  dffs1 \DFF_1164/Q_reg  ( .Q(WX8267), .CLK(CK), .DIN(WX8266) );
  dffs1 \DFF_1163/Q_reg  ( .Q(WX8265), .CLK(CK), .DIN(WX8264) );
  dffs1 \DFF_1162/Q_reg  ( .Q(WX8263), .CLK(CK), .DIN(WX8262) );
  dffs1 \DFF_1161/Q_reg  ( .Q(WX8261), .CLK(CK), .DIN(WX8260) );
  dffs1 \DFF_1160/Q_reg  ( .Q(WX8259), .CLK(CK), .DIN(WX8258) );
  dffs1 \DFF_1159/Q_reg  ( .Q(WX8257), .CLK(CK), .DIN(WX8256) );
  dffs1 \DFF_1158/Q_reg  ( .Q(WX8255), .CLK(CK), .DIN(WX8254) );
  dffs1 \DFF_1157/Q_reg  ( .Q(WX8253), .CLK(CK), .DIN(WX8252) );
  dffs1 \DFF_1156/Q_reg  ( .Q(WX8251), .CLK(CK), .DIN(WX8250) );
  dffs1 \DFF_1155/Q_reg  ( .Q(WX8249), .CLK(CK), .DIN(WX8248) );
  dffs1 \DFF_1154/Q_reg  ( .Q(WX8247), .CLK(CK), .DIN(WX8246) );
  dffs1 \DFF_1153/Q_reg  ( .Q(WX8245), .CLK(CK), .DIN(WX8244) );
  dffs1 \DFF_1152/Q_reg  ( .Q(WX8243), .CLK(CK), .DIN(WX8242) );
  dffs1 \DFF_1151/Q_reg  ( .Q(CRC_OUT_4_31), .CLK(CK), .DIN(WX7791) );
  dffs1 \DFF_1150/Q_reg  ( .Q(CRC_OUT_4_30), .CLK(CK), .DIN(WX7789) );
  dffs1 \DFF_1149/Q_reg  ( .Q(CRC_OUT_4_29), .CLK(CK), .DIN(WX7787) );
  dffs1 \DFF_1148/Q_reg  ( .Q(CRC_OUT_4_28), .CLK(CK), .DIN(WX7785) );
  dffs1 \DFF_1147/Q_reg  ( .Q(CRC_OUT_4_27), .CLK(CK), .DIN(WX7783) );
  dffs1 \DFF_1146/Q_reg  ( .Q(CRC_OUT_4_26), .CLK(CK), .DIN(WX7781) );
  dffs1 \DFF_1145/Q_reg  ( .Q(CRC_OUT_4_25), .CLK(CK), .DIN(WX7779) );
  dffs1 \DFF_1144/Q_reg  ( .Q(CRC_OUT_4_24), .CLK(CK), .DIN(WX7777) );
  dffs1 \DFF_1143/Q_reg  ( .Q(CRC_OUT_4_23), .CLK(CK), .DIN(WX7775) );
  dffs1 \DFF_1142/Q_reg  ( .Q(CRC_OUT_4_22), .CLK(CK), .DIN(WX7773) );
  dffs1 \DFF_1141/Q_reg  ( .Q(CRC_OUT_4_21), .CLK(CK), .DIN(WX7771) );
  dffs1 \DFF_1140/Q_reg  ( .Q(CRC_OUT_4_20), .CLK(CK), .DIN(WX7769) );
  dffs1 \DFF_1139/Q_reg  ( .Q(CRC_OUT_4_19), .CLK(CK), .DIN(WX7767) );
  dffs1 \DFF_1138/Q_reg  ( .Q(CRC_OUT_4_18), .CLK(CK), .DIN(WX7765) );
  dffs1 \DFF_1137/Q_reg  ( .Q(CRC_OUT_4_17), .CLK(CK), .DIN(WX7763) );
  dffs1 \DFF_1136/Q_reg  ( .Q(CRC_OUT_4_16), .CLK(CK), .DIN(WX7761) );
  dffs1 \DFF_1135/Q_reg  ( .Q(CRC_OUT_4_15), .CLK(CK), .DIN(WX7759) );
  dffs1 \DFF_1134/Q_reg  ( .Q(CRC_OUT_4_14), .CLK(CK), .DIN(WX7757) );
  dffs1 \DFF_1133/Q_reg  ( .Q(CRC_OUT_4_13), .CLK(CK), .DIN(WX7755) );
  dffs1 \DFF_1132/Q_reg  ( .Q(CRC_OUT_4_12), .CLK(CK), .DIN(WX7753) );
  dffs1 \DFF_1131/Q_reg  ( .Q(CRC_OUT_4_11), .CLK(CK), .DIN(WX7751) );
  dffs1 \DFF_1130/Q_reg  ( .Q(CRC_OUT_4_10), .CLK(CK), .DIN(WX7749) );
  dffs1 \DFF_1129/Q_reg  ( .Q(CRC_OUT_4_9), .CLK(CK), .DIN(WX7747) );
  dffs1 \DFF_1128/Q_reg  ( .Q(CRC_OUT_4_8), .CLK(CK), .DIN(WX7745) );
  dffs1 \DFF_1127/Q_reg  ( .Q(CRC_OUT_4_7), .CLK(CK), .DIN(WX7743) );
  dffs1 \DFF_1126/Q_reg  ( .Q(CRC_OUT_4_6), .CLK(CK), .DIN(WX7741) );
  dffs1 \DFF_1125/Q_reg  ( .Q(CRC_OUT_4_5), .CLK(CK), .DIN(WX7739) );
  dffs1 \DFF_1124/Q_reg  ( .Q(CRC_OUT_4_4), .CLK(CK), .DIN(WX7737) );
  dffs1 \DFF_1123/Q_reg  ( .Q(CRC_OUT_4_3), .CLK(CK), .DIN(WX7735) );
  dffs1 \DFF_1122/Q_reg  ( .Q(CRC_OUT_4_2), .CLK(CK), .DIN(WX7733) );
  dffs1 \DFF_1121/Q_reg  ( .Q(CRC_OUT_4_1), .CLK(CK), .DIN(WX7731) );
  dffs1 \DFF_1120/Q_reg  ( .Q(CRC_OUT_4_0), .CLK(CK), .DIN(WX7729) );
  dffs1 \DFF_1119/Q_reg  ( .QN(n3237), .Q(WX7364), .CLK(CK), .DIN(WX7363) );
  dffs1 \DFF_1118/Q_reg  ( .QN(n3238), .Q(WX7362), .CLK(CK), .DIN(WX7361) );
  dffs1 \DFF_1117/Q_reg  ( .QN(n3239), .Q(WX7360), .CLK(CK), .DIN(WX7359) );
  dffs1 \DFF_1116/Q_reg  ( .QN(n3240), .Q(WX7358), .CLK(CK), .DIN(WX7357) );
  dffs1 \DFF_1115/Q_reg  ( .QN(n3241), .Q(WX7356), .CLK(CK), .DIN(WX7355) );
  dffs1 \DFF_1114/Q_reg  ( .QN(n3242), .Q(WX7354), .CLK(CK), .DIN(WX7353) );
  dffs1 \DFF_1113/Q_reg  ( .QN(n3243), .Q(WX7352), .CLK(CK), .DIN(WX7351) );
  dffs1 \DFF_1112/Q_reg  ( .QN(n3244), .Q(WX7350), .CLK(CK), .DIN(WX7349) );
  dffs1 \DFF_1111/Q_reg  ( .QN(n3245), .Q(WX7348), .CLK(CK), .DIN(WX7347) );
  dffs1 \DFF_1110/Q_reg  ( .QN(n3246), .Q(WX7346), .CLK(CK), .DIN(WX7345) );
  dffs1 \DFF_1109/Q_reg  ( .QN(n3247), .Q(WX7344), .CLK(CK), .DIN(WX7343) );
  dffs1 \DFF_1108/Q_reg  ( .QN(n3248), .Q(WX7342), .CLK(CK), .DIN(WX7341) );
  dffs1 \DFF_1107/Q_reg  ( .QN(n3249), .Q(WX7340), .CLK(CK), .DIN(WX7339) );
  dffs1 \DFF_1106/Q_reg  ( .QN(n3250), .Q(WX7338), .CLK(CK), .DIN(WX7337) );
  dffs1 \DFF_1105/Q_reg  ( .QN(n3251), .Q(WX7336), .CLK(CK), .DIN(WX7335) );
  dffs1 \DFF_1104/Q_reg  ( .QN(n3252), .Q(WX7334), .CLK(CK), .DIN(WX7333) );
  dffs1 \DFF_1103/Q_reg  ( .Q(WX7332), .CLK(CK), .DIN(WX7331) );
  dffs1 \DFF_1102/Q_reg  ( .Q(WX7330), .CLK(CK), .DIN(WX7329) );
  dffs1 \DFF_1101/Q_reg  ( .Q(WX7328), .CLK(CK), .DIN(WX7327) );
  dffs1 \DFF_1100/Q_reg  ( .Q(WX7326), .CLK(CK), .DIN(WX7325) );
  dffs1 \DFF_1099/Q_reg  ( .Q(WX7324), .CLK(CK), .DIN(WX7323) );
  dffs1 \DFF_1098/Q_reg  ( .Q(WX7322), .CLK(CK), .DIN(WX7321) );
  dffs1 \DFF_1097/Q_reg  ( .Q(WX7320), .CLK(CK), .DIN(WX7319) );
  dffs1 \DFF_1096/Q_reg  ( .Q(WX7318), .CLK(CK), .DIN(WX7317) );
  dffs1 \DFF_1095/Q_reg  ( .Q(WX7316), .CLK(CK), .DIN(WX7315) );
  dffs1 \DFF_1094/Q_reg  ( .Q(WX7314), .CLK(CK), .DIN(WX7313) );
  dffs1 \DFF_1093/Q_reg  ( .Q(WX7312), .CLK(CK), .DIN(WX7311) );
  dffs1 \DFF_1092/Q_reg  ( .Q(WX7310), .CLK(CK), .DIN(WX7309) );
  dffs1 \DFF_1091/Q_reg  ( .Q(WX7308), .CLK(CK), .DIN(WX7307) );
  dffs1 \DFF_1090/Q_reg  ( .Q(WX7306), .CLK(CK), .DIN(WX7305) );
  dffs1 \DFF_1089/Q_reg  ( .Q(WX7304), .CLK(CK), .DIN(WX7303) );
  dffs1 \DFF_1088/Q_reg  ( .Q(WX7302), .CLK(CK), .DIN(WX7301) );
  dffs1 \DFF_1087/Q_reg  ( .Q(WX7300), .CLK(CK), .DIN(WX7299) );
  dffs1 \DFF_1086/Q_reg  ( .Q(WX7298), .CLK(CK), .DIN(WX7297) );
  dffs1 \DFF_1085/Q_reg  ( .Q(WX7296), .CLK(CK), .DIN(WX7295) );
  dffs1 \DFF_1084/Q_reg  ( .Q(WX7294), .CLK(CK), .DIN(WX7293) );
  dffs1 \DFF_1083/Q_reg  ( .Q(WX7292), .CLK(CK), .DIN(WX7291) );
  dffs1 \DFF_1082/Q_reg  ( .Q(WX7290), .CLK(CK), .DIN(WX7289) );
  dffs1 \DFF_1081/Q_reg  ( .Q(WX7288), .CLK(CK), .DIN(WX7287) );
  dffs1 \DFF_1080/Q_reg  ( .Q(WX7286), .CLK(CK), .DIN(WX7285) );
  dffs1 \DFF_1079/Q_reg  ( .Q(WX7284), .CLK(CK), .DIN(WX7283) );
  dffs1 \DFF_1078/Q_reg  ( .Q(WX7282), .CLK(CK), .DIN(WX7281) );
  dffs1 \DFF_1077/Q_reg  ( .Q(WX7280), .CLK(CK), .DIN(WX7279) );
  dffs1 \DFF_1076/Q_reg  ( .Q(WX7278), .CLK(CK), .DIN(WX7277) );
  dffs1 \DFF_1075/Q_reg  ( .Q(WX7276), .CLK(CK), .DIN(WX7275) );
  dffs1 \DFF_1074/Q_reg  ( .Q(WX7274), .CLK(CK), .DIN(WX7273) );
  dffs1 \DFF_1073/Q_reg  ( .Q(WX7272), .CLK(CK), .DIN(WX7271) );
  dffs1 \DFF_1072/Q_reg  ( .Q(WX7270), .CLK(CK), .DIN(WX7269) );
  dffs1 \DFF_1071/Q_reg  ( .Q(WX7268), .CLK(CK), .DIN(WX7267) );
  dffs1 \DFF_1070/Q_reg  ( .Q(WX7266), .CLK(CK), .DIN(WX7265) );
  dffs1 \DFF_1069/Q_reg  ( .Q(WX7264), .CLK(CK), .DIN(WX7263) );
  dffs1 \DFF_1068/Q_reg  ( .Q(WX7262), .CLK(CK), .DIN(WX7261) );
  dffs1 \DFF_1067/Q_reg  ( .Q(WX7260), .CLK(CK), .DIN(WX7259) );
  dffs1 \DFF_1066/Q_reg  ( .Q(WX7258), .CLK(CK), .DIN(WX7257) );
  dffs1 \DFF_1065/Q_reg  ( .Q(WX7256), .CLK(CK), .DIN(WX7255) );
  dffs1 \DFF_1064/Q_reg  ( .Q(WX7254), .CLK(CK), .DIN(WX7253) );
  dffs1 \DFF_1063/Q_reg  ( .Q(WX7252), .CLK(CK), .DIN(WX7251) );
  dffs1 \DFF_1062/Q_reg  ( .Q(WX7250), .CLK(CK), .DIN(WX7249) );
  dffs1 \DFF_1061/Q_reg  ( .Q(WX7248), .CLK(CK), .DIN(WX7247) );
  dffs1 \DFF_1060/Q_reg  ( .Q(WX7246), .CLK(CK), .DIN(WX7245) );
  dffs1 \DFF_1059/Q_reg  ( .Q(WX7244), .CLK(CK), .DIN(WX7243) );
  dffs1 \DFF_1058/Q_reg  ( .Q(WX7242), .CLK(CK), .DIN(WX7241) );
  dffs1 \DFF_1057/Q_reg  ( .Q(WX7240), .CLK(CK), .DIN(WX7239) );
  dffs1 \DFF_1056/Q_reg  ( .Q(WX7238), .CLK(CK), .DIN(WX7237) );
  dffs1 \DFF_1055/Q_reg  ( .Q(WX7236), .CLK(CK), .DIN(WX7235) );
  dffs1 \DFF_1054/Q_reg  ( .Q(WX7234), .CLK(CK), .DIN(WX7233) );
  dffs1 \DFF_1053/Q_reg  ( .Q(WX7232), .CLK(CK), .DIN(WX7231) );
  dffs1 \DFF_1052/Q_reg  ( .Q(WX7230), .CLK(CK), .DIN(WX7229) );
  dffs1 \DFF_1051/Q_reg  ( .Q(WX7228), .CLK(CK), .DIN(WX7227) );
  dffs1 \DFF_1050/Q_reg  ( .Q(WX7226), .CLK(CK), .DIN(WX7225) );
  dffs1 \DFF_1049/Q_reg  ( .Q(WX7224), .CLK(CK), .DIN(WX7223) );
  dffs1 \DFF_1048/Q_reg  ( .Q(WX7222), .CLK(CK), .DIN(WX7221) );
  dffs1 \DFF_1047/Q_reg  ( .Q(WX7220), .CLK(CK), .DIN(WX7219) );
  dffs1 \DFF_1046/Q_reg  ( .Q(WX7218), .CLK(CK), .DIN(WX7217) );
  dffs1 \DFF_1045/Q_reg  ( .Q(WX7216), .CLK(CK), .DIN(WX7215) );
  dffs1 \DFF_1044/Q_reg  ( .Q(WX7214), .CLK(CK), .DIN(WX7213) );
  dffs1 \DFF_1043/Q_reg  ( .Q(WX7212), .CLK(CK), .DIN(WX7211) );
  dffs1 \DFF_1042/Q_reg  ( .Q(WX7210), .CLK(CK), .DIN(WX7209) );
  dffs1 \DFF_1041/Q_reg  ( .Q(WX7208), .CLK(CK), .DIN(WX7207) );
  dffs1 \DFF_1040/Q_reg  ( .Q(WX7206), .CLK(CK), .DIN(WX7205) );
  dffs1 \DFF_1039/Q_reg  ( .QN(n2981), .CLK(CK), .DIN(WX7203) );
  dffs1 \DFF_1038/Q_reg  ( .QN(n2982), .CLK(CK), .DIN(WX7201) );
  dffs1 \DFF_1037/Q_reg  ( .QN(n2983), .CLK(CK), .DIN(WX7199) );
  dffs1 \DFF_1036/Q_reg  ( .QN(n2984), .CLK(CK), .DIN(WX7197) );
  dffs1 \DFF_1035/Q_reg  ( .QN(n2985), .CLK(CK), .DIN(WX7195) );
  dffs1 \DFF_1034/Q_reg  ( .QN(n2986), .CLK(CK), .DIN(WX7193) );
  dffs1 \DFF_1033/Q_reg  ( .QN(n2987), .CLK(CK), .DIN(WX7191) );
  dffs1 \DFF_1032/Q_reg  ( .QN(n2988), .CLK(CK), .DIN(WX7189) );
  dffs1 \DFF_1031/Q_reg  ( .QN(n2989), .CLK(CK), .DIN(WX7187) );
  dffs1 \DFF_1030/Q_reg  ( .QN(n2990), .CLK(CK), .DIN(WX7185) );
  dffs1 \DFF_1029/Q_reg  ( .QN(n2991), .CLK(CK), .DIN(WX7183) );
  dffs1 \DFF_1028/Q_reg  ( .QN(n2992), .CLK(CK), .DIN(WX7181) );
  dffs1 \DFF_1027/Q_reg  ( .QN(n2993), .CLK(CK), .DIN(WX7179) );
  dffs1 \DFF_1026/Q_reg  ( .QN(n2994), .CLK(CK), .DIN(WX7177) );
  dffs1 \DFF_1025/Q_reg  ( .QN(n2995), .CLK(CK), .DIN(WX7175) );
  dffs1 \DFF_1024/Q_reg  ( .QN(n2996), .CLK(CK), .DIN(WX7173) );
  dffs1 \DFF_1023/Q_reg  ( .QN(n3141), .CLK(CK), .DIN(WX7171) );
  dffs1 \DFF_1022/Q_reg  ( .QN(n3142), .CLK(CK), .DIN(WX7169) );
  dffs1 \DFF_1021/Q_reg  ( .QN(n3143), .CLK(CK), .DIN(WX7167) );
  dffs1 \DFF_1020/Q_reg  ( .QN(n3144), .CLK(CK), .DIN(WX7165) );
  dffs1 \DFF_1019/Q_reg  ( .QN(n3145), .CLK(CK), .DIN(WX7163) );
  dffs1 \DFF_1018/Q_reg  ( .QN(n3146), .CLK(CK), .DIN(WX7161) );
  dffs1 \DFF_1017/Q_reg  ( .QN(n3147), .CLK(CK), .DIN(WX7159) );
  dffs1 \DFF_1016/Q_reg  ( .QN(n3148), .CLK(CK), .DIN(WX7157) );
  dffs1 \DFF_1015/Q_reg  ( .QN(n3149), .CLK(CK), .DIN(WX7155) );
  dffs1 \DFF_1014/Q_reg  ( .QN(n3150), .CLK(CK), .DIN(WX7153) );
  dffs1 \DFF_1013/Q_reg  ( .QN(n3151), .CLK(CK), .DIN(WX7151) );
  dffs1 \DFF_1012/Q_reg  ( .QN(n3152), .CLK(CK), .DIN(WX7149) );
  dffs1 \DFF_1011/Q_reg  ( .QN(n3153), .CLK(CK), .DIN(WX7147) );
  dffs1 \DFF_1010/Q_reg  ( .QN(n3154), .CLK(CK), .DIN(WX7145) );
  dffs1 \DFF_1009/Q_reg  ( .QN(n3155), .CLK(CK), .DIN(WX7143) );
  dffs1 \DFF_1008/Q_reg  ( .QN(n3156), .CLK(CK), .DIN(WX7141) );
  dffs1 \DFF_1007/Q_reg  ( .Q(WX7140), .CLK(CK), .DIN(WX7139) );
  dffs1 \DFF_1006/Q_reg  ( .Q(WX7138), .CLK(CK), .DIN(WX7137) );
  dffs1 \DFF_1005/Q_reg  ( .Q(WX7136), .CLK(CK), .DIN(WX7135) );
  dffs1 \DFF_1004/Q_reg  ( .Q(WX7134), .CLK(CK), .DIN(WX7133) );
  dffs1 \DFF_1003/Q_reg  ( .Q(WX7132), .CLK(CK), .DIN(WX7131) );
  dffs1 \DFF_1002/Q_reg  ( .Q(WX7130), .CLK(CK), .DIN(WX7129) );
  dffs1 \DFF_1001/Q_reg  ( .Q(WX7128), .CLK(CK), .DIN(WX7127) );
  dffs1 \DFF_1000/Q_reg  ( .Q(WX7126), .CLK(CK), .DIN(WX7125) );
  dffs1 \DFF_999/Q_reg  ( .Q(WX7124), .CLK(CK), .DIN(WX7123) );
  dffs1 \DFF_998/Q_reg  ( .Q(WX7122), .CLK(CK), .DIN(WX7121) );
  dffs1 \DFF_997/Q_reg  ( .Q(WX7120), .CLK(CK), .DIN(WX7119) );
  dffs1 \DFF_996/Q_reg  ( .Q(WX7118), .CLK(CK), .DIN(WX7117) );
  dffs1 \DFF_995/Q_reg  ( .Q(WX7116), .CLK(CK), .DIN(WX7115) );
  dffs1 \DFF_994/Q_reg  ( .Q(WX7114), .CLK(CK), .DIN(WX7113) );
  dffs1 \DFF_993/Q_reg  ( .Q(WX7112), .CLK(CK), .DIN(WX7111) );
  dffs1 \DFF_992/Q_reg  ( .Q(WX7110), .CLK(CK), .DIN(WX7109) );
  dffs1 \DFF_991/Q_reg  ( .Q(WX7012), .CLK(CK), .DIN(WX7011) );
  dffs1 \DFF_990/Q_reg  ( .Q(WX7010), .CLK(CK), .DIN(WX7009) );
  dffs1 \DFF_989/Q_reg  ( .Q(WX7008), .CLK(CK), .DIN(WX7007) );
  dffs1 \DFF_988/Q_reg  ( .Q(WX7006), .CLK(CK), .DIN(WX7005) );
  dffs1 \DFF_987/Q_reg  ( .Q(WX7004), .CLK(CK), .DIN(WX7003) );
  dffs1 \DFF_986/Q_reg  ( .Q(WX7002), .CLK(CK), .DIN(WX7001) );
  dffs1 \DFF_985/Q_reg  ( .Q(WX7000), .CLK(CK), .DIN(WX6999) );
  dffs1 \DFF_984/Q_reg  ( .Q(WX6998), .CLK(CK), .DIN(WX6997) );
  dffs1 \DFF_983/Q_reg  ( .Q(WX6996), .CLK(CK), .DIN(WX6995) );
  dffs1 \DFF_982/Q_reg  ( .Q(WX6994), .CLK(CK), .DIN(WX6993) );
  dffs1 \DFF_981/Q_reg  ( .Q(WX6992), .CLK(CK), .DIN(WX6991) );
  dffs1 \DFF_980/Q_reg  ( .Q(WX6990), .CLK(CK), .DIN(WX6989) );
  dffs1 \DFF_979/Q_reg  ( .Q(WX6988), .CLK(CK), .DIN(WX6987) );
  dffs1 \DFF_978/Q_reg  ( .Q(WX6986), .CLK(CK), .DIN(WX6985) );
  dffs1 \DFF_977/Q_reg  ( .Q(WX6984), .CLK(CK), .DIN(WX6983) );
  dffs1 \DFF_976/Q_reg  ( .Q(WX6982), .CLK(CK), .DIN(WX6981) );
  dffs1 \DFF_975/Q_reg  ( .Q(WX6980), .CLK(CK), .DIN(WX6979) );
  dffs1 \DFF_974/Q_reg  ( .Q(WX6978), .CLK(CK), .DIN(WX6977) );
  dffs1 \DFF_973/Q_reg  ( .Q(WX6976), .CLK(CK), .DIN(WX6975) );
  dffs1 \DFF_972/Q_reg  ( .Q(WX6974), .CLK(CK), .DIN(WX6973) );
  dffs1 \DFF_971/Q_reg  ( .Q(WX6972), .CLK(CK), .DIN(WX6971) );
  dffs1 \DFF_970/Q_reg  ( .Q(WX6970), .CLK(CK), .DIN(WX6969) );
  dffs1 \DFF_969/Q_reg  ( .Q(WX6968), .CLK(CK), .DIN(WX6967) );
  dffs1 \DFF_968/Q_reg  ( .Q(WX6966), .CLK(CK), .DIN(WX6965) );
  dffs1 \DFF_967/Q_reg  ( .Q(WX6964), .CLK(CK), .DIN(WX6963) );
  dffs1 \DFF_966/Q_reg  ( .Q(WX6962), .CLK(CK), .DIN(WX6961) );
  dffs1 \DFF_965/Q_reg  ( .Q(WX6960), .CLK(CK), .DIN(WX6959) );
  dffs1 \DFF_964/Q_reg  ( .Q(WX6958), .CLK(CK), .DIN(WX6957) );
  dffs1 \DFF_963/Q_reg  ( .Q(WX6956), .CLK(CK), .DIN(WX6955) );
  dffs1 \DFF_962/Q_reg  ( .Q(WX6954), .CLK(CK), .DIN(WX6953) );
  dffs1 \DFF_961/Q_reg  ( .Q(WX6952), .CLK(CK), .DIN(WX6951) );
  dffs1 \DFF_960/Q_reg  ( .Q(WX6950), .CLK(CK), .DIN(WX6949) );
  dffs1 \DFF_959/Q_reg  ( .Q(CRC_OUT_5_31), .CLK(CK), .DIN(WX6498) );
  dffs1 \DFF_958/Q_reg  ( .Q(CRC_OUT_5_30), .CLK(CK), .DIN(WX6496) );
  dffs1 \DFF_957/Q_reg  ( .Q(CRC_OUT_5_29), .CLK(CK), .DIN(WX6494) );
  dffs1 \DFF_956/Q_reg  ( .Q(CRC_OUT_5_28), .CLK(CK), .DIN(WX6492) );
  dffs1 \DFF_955/Q_reg  ( .Q(CRC_OUT_5_27), .CLK(CK), .DIN(WX6490) );
  dffs1 \DFF_954/Q_reg  ( .Q(CRC_OUT_5_26), .CLK(CK), .DIN(WX6488) );
  dffs1 \DFF_953/Q_reg  ( .Q(CRC_OUT_5_25), .CLK(CK), .DIN(WX6486) );
  dffs1 \DFF_952/Q_reg  ( .Q(CRC_OUT_5_24), .CLK(CK), .DIN(WX6484) );
  dffs1 \DFF_951/Q_reg  ( .Q(CRC_OUT_5_23), .CLK(CK), .DIN(WX6482) );
  dffs1 \DFF_950/Q_reg  ( .Q(CRC_OUT_5_22), .CLK(CK), .DIN(WX6480) );
  dffs1 \DFF_949/Q_reg  ( .Q(CRC_OUT_5_21), .CLK(CK), .DIN(WX6478) );
  dffs1 \DFF_948/Q_reg  ( .Q(CRC_OUT_5_20), .CLK(CK), .DIN(WX6476) );
  dffs1 \DFF_947/Q_reg  ( .Q(CRC_OUT_5_19), .CLK(CK), .DIN(WX6474) );
  dffs1 \DFF_946/Q_reg  ( .Q(CRC_OUT_5_18), .CLK(CK), .DIN(WX6472) );
  dffs1 \DFF_945/Q_reg  ( .Q(CRC_OUT_5_17), .CLK(CK), .DIN(WX6470) );
  dffs1 \DFF_944/Q_reg  ( .Q(CRC_OUT_5_16), .CLK(CK), .DIN(WX6468) );
  dffs1 \DFF_943/Q_reg  ( .Q(CRC_OUT_5_15), .CLK(CK), .DIN(WX6466) );
  dffs1 \DFF_942/Q_reg  ( .Q(CRC_OUT_5_14), .CLK(CK), .DIN(WX6464) );
  dffs1 \DFF_941/Q_reg  ( .Q(CRC_OUT_5_13), .CLK(CK), .DIN(WX6462) );
  dffs1 \DFF_940/Q_reg  ( .Q(CRC_OUT_5_12), .CLK(CK), .DIN(WX6460) );
  dffs1 \DFF_939/Q_reg  ( .Q(CRC_OUT_5_11), .CLK(CK), .DIN(WX6458) );
  dffs1 \DFF_938/Q_reg  ( .Q(CRC_OUT_5_10), .CLK(CK), .DIN(WX6456) );
  dffs1 \DFF_937/Q_reg  ( .Q(CRC_OUT_5_9), .CLK(CK), .DIN(WX6454) );
  dffs1 \DFF_936/Q_reg  ( .Q(CRC_OUT_5_8), .CLK(CK), .DIN(WX6452) );
  dffs1 \DFF_935/Q_reg  ( .Q(CRC_OUT_5_7), .CLK(CK), .DIN(WX6450) );
  dffs1 \DFF_934/Q_reg  ( .Q(CRC_OUT_5_6), .CLK(CK), .DIN(WX6448) );
  dffs1 \DFF_933/Q_reg  ( .Q(CRC_OUT_5_5), .CLK(CK), .DIN(WX6446) );
  dffs1 \DFF_932/Q_reg  ( .Q(CRC_OUT_5_4), .CLK(CK), .DIN(WX6444) );
  dffs1 \DFF_931/Q_reg  ( .Q(CRC_OUT_5_3), .CLK(CK), .DIN(WX6442) );
  dffs1 \DFF_930/Q_reg  ( .Q(CRC_OUT_5_2), .CLK(CK), .DIN(WX6440) );
  dffs1 \DFF_929/Q_reg  ( .Q(CRC_OUT_5_1), .CLK(CK), .DIN(WX6438) );
  dffs1 \DFF_928/Q_reg  ( .Q(CRC_OUT_5_0), .CLK(CK), .DIN(WX6436) );
  dffs1 \DFF_927/Q_reg  ( .QN(n3253), .Q(WX6071), .CLK(CK), .DIN(WX6070) );
  dffs1 \DFF_926/Q_reg  ( .QN(n3254), .Q(WX6069), .CLK(CK), .DIN(WX6068) );
  dffs1 \DFF_925/Q_reg  ( .QN(n3255), .Q(WX6067), .CLK(CK), .DIN(WX6066) );
  dffs1 \DFF_924/Q_reg  ( .QN(n3256), .Q(WX6065), .CLK(CK), .DIN(WX6064) );
  dffs1 \DFF_923/Q_reg  ( .QN(n3257), .Q(WX6063), .CLK(CK), .DIN(WX6062) );
  dffs1 \DFF_922/Q_reg  ( .QN(n3258), .Q(WX6061), .CLK(CK), .DIN(WX6060) );
  dffs1 \DFF_921/Q_reg  ( .QN(n3259), .Q(WX6059), .CLK(CK), .DIN(WX6058) );
  dffs1 \DFF_920/Q_reg  ( .QN(n3260), .Q(WX6057), .CLK(CK), .DIN(WX6056) );
  dffs1 \DFF_919/Q_reg  ( .QN(n3261), .Q(WX6055), .CLK(CK), .DIN(WX6054) );
  dffs1 \DFF_918/Q_reg  ( .QN(n3262), .Q(WX6053), .CLK(CK), .DIN(WX6052) );
  dffs1 \DFF_917/Q_reg  ( .QN(n3263), .Q(WX6051), .CLK(CK), .DIN(WX6050) );
  dffs1 \DFF_916/Q_reg  ( .QN(n3264), .Q(WX6049), .CLK(CK), .DIN(WX6048) );
  dffs1 \DFF_915/Q_reg  ( .QN(n3265), .Q(WX6047), .CLK(CK), .DIN(WX6046) );
  dffs1 \DFF_914/Q_reg  ( .QN(n3266), .Q(WX6045), .CLK(CK), .DIN(WX6044) );
  dffs1 \DFF_913/Q_reg  ( .QN(n3267), .Q(WX6043), .CLK(CK), .DIN(WX6042) );
  dffs1 \DFF_912/Q_reg  ( .QN(n3268), .Q(WX6041), .CLK(CK), .DIN(WX6040) );
  dffs1 \DFF_911/Q_reg  ( .Q(WX6039), .CLK(CK), .DIN(WX6038) );
  dffs1 \DFF_910/Q_reg  ( .Q(WX6037), .CLK(CK), .DIN(WX6036) );
  dffs1 \DFF_909/Q_reg  ( .Q(WX6035), .CLK(CK), .DIN(WX6034) );
  dffs1 \DFF_908/Q_reg  ( .Q(WX6033), .CLK(CK), .DIN(WX6032) );
  dffs1 \DFF_907/Q_reg  ( .Q(WX6031), .CLK(CK), .DIN(WX6030) );
  dffs1 \DFF_906/Q_reg  ( .Q(WX6029), .CLK(CK), .DIN(WX6028) );
  dffs1 \DFF_905/Q_reg  ( .Q(WX6027), .CLK(CK), .DIN(WX6026) );
  dffs1 \DFF_904/Q_reg  ( .Q(WX6025), .CLK(CK), .DIN(WX6024) );
  dffs1 \DFF_903/Q_reg  ( .Q(WX6023), .CLK(CK), .DIN(WX6022) );
  dffs1 \DFF_902/Q_reg  ( .Q(WX6021), .CLK(CK), .DIN(WX6020) );
  dffs1 \DFF_901/Q_reg  ( .Q(WX6019), .CLK(CK), .DIN(WX6018) );
  dffs1 \DFF_900/Q_reg  ( .Q(WX6017), .CLK(CK), .DIN(WX6016) );
  dffs1 \DFF_899/Q_reg  ( .Q(WX6015), .CLK(CK), .DIN(WX6014) );
  dffs1 \DFF_898/Q_reg  ( .Q(WX6013), .CLK(CK), .DIN(WX6012) );
  dffs1 \DFF_897/Q_reg  ( .Q(WX6011), .CLK(CK), .DIN(WX6010) );
  dffs1 \DFF_896/Q_reg  ( .Q(WX6009), .CLK(CK), .DIN(WX6008) );
  dffs1 \DFF_895/Q_reg  ( .Q(WX6007), .CLK(CK), .DIN(WX6006) );
  dffs1 \DFF_894/Q_reg  ( .Q(WX6005), .CLK(CK), .DIN(WX6004) );
  dffs1 \DFF_893/Q_reg  ( .Q(WX6003), .CLK(CK), .DIN(WX6002) );
  dffs1 \DFF_892/Q_reg  ( .Q(WX6001), .CLK(CK), .DIN(WX6000) );
  dffs1 \DFF_891/Q_reg  ( .Q(WX5999), .CLK(CK), .DIN(WX5998) );
  dffs1 \DFF_890/Q_reg  ( .Q(WX5997), .CLK(CK), .DIN(WX5996) );
  dffs1 \DFF_889/Q_reg  ( .Q(WX5995), .CLK(CK), .DIN(WX5994) );
  dffs1 \DFF_888/Q_reg  ( .Q(WX5993), .CLK(CK), .DIN(WX5992) );
  dffs1 \DFF_887/Q_reg  ( .Q(WX5991), .CLK(CK), .DIN(WX5990) );
  dffs1 \DFF_886/Q_reg  ( .Q(WX5989), .CLK(CK), .DIN(WX5988) );
  dffs1 \DFF_885/Q_reg  ( .Q(WX5987), .CLK(CK), .DIN(WX5986) );
  dffs1 \DFF_884/Q_reg  ( .Q(WX5985), .CLK(CK), .DIN(WX5984) );
  dffs1 \DFF_883/Q_reg  ( .Q(WX5983), .CLK(CK), .DIN(WX5982) );
  dffs1 \DFF_882/Q_reg  ( .Q(WX5981), .CLK(CK), .DIN(WX5980) );
  dffs1 \DFF_881/Q_reg  ( .Q(WX5979), .CLK(CK), .DIN(WX5978) );
  dffs1 \DFF_880/Q_reg  ( .Q(WX5977), .CLK(CK), .DIN(WX5976) );
  dffs1 \DFF_879/Q_reg  ( .Q(WX5975), .CLK(CK), .DIN(WX5974) );
  dffs1 \DFF_878/Q_reg  ( .Q(WX5973), .CLK(CK), .DIN(WX5972) );
  dffs1 \DFF_877/Q_reg  ( .Q(WX5971), .CLK(CK), .DIN(WX5970) );
  dffs1 \DFF_876/Q_reg  ( .Q(WX5969), .CLK(CK), .DIN(WX5968) );
  dffs1 \DFF_875/Q_reg  ( .Q(WX5967), .CLK(CK), .DIN(WX5966) );
  dffs1 \DFF_874/Q_reg  ( .Q(WX5965), .CLK(CK), .DIN(WX5964) );
  dffs1 \DFF_873/Q_reg  ( .Q(WX5963), .CLK(CK), .DIN(WX5962) );
  dffs1 \DFF_872/Q_reg  ( .Q(WX5961), .CLK(CK), .DIN(WX5960) );
  dffs1 \DFF_871/Q_reg  ( .Q(WX5959), .CLK(CK), .DIN(WX5958) );
  dffs1 \DFF_870/Q_reg  ( .Q(WX5957), .CLK(CK), .DIN(WX5956) );
  dffs1 \DFF_869/Q_reg  ( .Q(WX5955), .CLK(CK), .DIN(WX5954) );
  dffs1 \DFF_868/Q_reg  ( .Q(WX5953), .CLK(CK), .DIN(WX5952) );
  dffs1 \DFF_867/Q_reg  ( .Q(WX5951), .CLK(CK), .DIN(WX5950) );
  dffs1 \DFF_866/Q_reg  ( .Q(WX5949), .CLK(CK), .DIN(WX5948) );
  dffs1 \DFF_865/Q_reg  ( .Q(WX5947), .CLK(CK), .DIN(WX5946) );
  dffs1 \DFF_864/Q_reg  ( .Q(WX5945), .CLK(CK), .DIN(WX5944) );
  dffs1 \DFF_863/Q_reg  ( .Q(WX5943), .CLK(CK), .DIN(WX5942) );
  dffs1 \DFF_862/Q_reg  ( .Q(WX5941), .CLK(CK), .DIN(WX5940) );
  dffs1 \DFF_861/Q_reg  ( .Q(WX5939), .CLK(CK), .DIN(WX5938) );
  dffs1 \DFF_860/Q_reg  ( .Q(WX5937), .CLK(CK), .DIN(WX5936) );
  dffs1 \DFF_859/Q_reg  ( .Q(WX5935), .CLK(CK), .DIN(WX5934) );
  dffs1 \DFF_858/Q_reg  ( .Q(WX5933), .CLK(CK), .DIN(WX5932) );
  dffs1 \DFF_857/Q_reg  ( .Q(WX5931), .CLK(CK), .DIN(WX5930) );
  dffs1 \DFF_856/Q_reg  ( .Q(WX5929), .CLK(CK), .DIN(WX5928) );
  dffs1 \DFF_855/Q_reg  ( .Q(WX5927), .CLK(CK), .DIN(WX5926) );
  dffs1 \DFF_854/Q_reg  ( .Q(WX5925), .CLK(CK), .DIN(WX5924) );
  dffs1 \DFF_853/Q_reg  ( .Q(WX5923), .CLK(CK), .DIN(WX5922) );
  dffs1 \DFF_852/Q_reg  ( .Q(WX5921), .CLK(CK), .DIN(WX5920) );
  dffs1 \DFF_851/Q_reg  ( .Q(WX5919), .CLK(CK), .DIN(WX5918) );
  dffs1 \DFF_850/Q_reg  ( .Q(WX5917), .CLK(CK), .DIN(WX5916) );
  dffs1 \DFF_849/Q_reg  ( .Q(WX5915), .CLK(CK), .DIN(WX5914) );
  dffs1 \DFF_848/Q_reg  ( .Q(WX5913), .CLK(CK), .DIN(WX5912) );
  dffs1 \DFF_847/Q_reg  ( .QN(n2997), .CLK(CK), .DIN(WX5910) );
  dffs1 \DFF_846/Q_reg  ( .QN(n2998), .CLK(CK), .DIN(WX5908) );
  dffs1 \DFF_845/Q_reg  ( .QN(n2999), .CLK(CK), .DIN(WX5906) );
  dffs1 \DFF_844/Q_reg  ( .QN(n3000), .CLK(CK), .DIN(WX5904) );
  dffs1 \DFF_843/Q_reg  ( .QN(n3001), .CLK(CK), .DIN(WX5902) );
  dffs1 \DFF_842/Q_reg  ( .QN(n3002), .CLK(CK), .DIN(WX5900) );
  dffs1 \DFF_841/Q_reg  ( .QN(n3003), .CLK(CK), .DIN(WX5898) );
  dffs1 \DFF_840/Q_reg  ( .QN(n3004), .CLK(CK), .DIN(WX5896) );
  dffs1 \DFF_839/Q_reg  ( .QN(n3005), .CLK(CK), .DIN(WX5894) );
  dffs1 \DFF_838/Q_reg  ( .QN(n3006), .CLK(CK), .DIN(WX5892) );
  dffs1 \DFF_837/Q_reg  ( .QN(n3007), .CLK(CK), .DIN(WX5890) );
  dffs1 \DFF_836/Q_reg  ( .QN(n3008), .CLK(CK), .DIN(WX5888) );
  dffs1 \DFF_835/Q_reg  ( .QN(n3009), .CLK(CK), .DIN(WX5886) );
  dffs1 \DFF_834/Q_reg  ( .QN(n3010), .CLK(CK), .DIN(WX5884) );
  dffs1 \DFF_833/Q_reg  ( .QN(n3011), .CLK(CK), .DIN(WX5882) );
  dffs1 \DFF_832/Q_reg  ( .QN(n3012), .CLK(CK), .DIN(WX5880) );
  dffs1 \DFF_831/Q_reg  ( .QN(n3157), .CLK(CK), .DIN(WX5878) );
  dffs1 \DFF_830/Q_reg  ( .QN(n3158), .CLK(CK), .DIN(WX5876) );
  dffs1 \DFF_829/Q_reg  ( .QN(n3159), .CLK(CK), .DIN(WX5874) );
  dffs1 \DFF_828/Q_reg  ( .QN(n3160), .CLK(CK), .DIN(WX5872) );
  dffs1 \DFF_827/Q_reg  ( .QN(n3161), .CLK(CK), .DIN(WX5870) );
  dffs1 \DFF_826/Q_reg  ( .QN(n3162), .CLK(CK), .DIN(WX5868) );
  dffs1 \DFF_825/Q_reg  ( .QN(n3163), .CLK(CK), .DIN(WX5866) );
  dffs1 \DFF_824/Q_reg  ( .QN(n3164), .CLK(CK), .DIN(WX5864) );
  dffs1 \DFF_823/Q_reg  ( .QN(n3165), .CLK(CK), .DIN(WX5862) );
  dffs1 \DFF_822/Q_reg  ( .QN(n3166), .CLK(CK), .DIN(WX5860) );
  dffs1 \DFF_821/Q_reg  ( .QN(n3167), .CLK(CK), .DIN(WX5858) );
  dffs1 \DFF_820/Q_reg  ( .QN(n3168), .CLK(CK), .DIN(WX5856) );
  dffs1 \DFF_819/Q_reg  ( .QN(n3169), .CLK(CK), .DIN(WX5854) );
  dffs1 \DFF_818/Q_reg  ( .QN(n3170), .CLK(CK), .DIN(WX5852) );
  dffs1 \DFF_817/Q_reg  ( .QN(n3171), .CLK(CK), .DIN(WX5850) );
  dffs1 \DFF_816/Q_reg  ( .QN(n3172), .CLK(CK), .DIN(WX5848) );
  dffs1 \DFF_815/Q_reg  ( .Q(WX5847), .CLK(CK), .DIN(WX5846) );
  dffs1 \DFF_814/Q_reg  ( .Q(WX5845), .CLK(CK), .DIN(WX5844) );
  dffs1 \DFF_813/Q_reg  ( .Q(WX5843), .CLK(CK), .DIN(WX5842) );
  dffs1 \DFF_812/Q_reg  ( .Q(WX5841), .CLK(CK), .DIN(WX5840) );
  dffs1 \DFF_811/Q_reg  ( .Q(WX5839), .CLK(CK), .DIN(WX5838) );
  dffs1 \DFF_810/Q_reg  ( .Q(WX5837), .CLK(CK), .DIN(WX5836) );
  dffs1 \DFF_809/Q_reg  ( .Q(WX5835), .CLK(CK), .DIN(WX5834) );
  dffs1 \DFF_808/Q_reg  ( .Q(WX5833), .CLK(CK), .DIN(WX5832) );
  dffs1 \DFF_807/Q_reg  ( .Q(WX5831), .CLK(CK), .DIN(WX5830) );
  dffs1 \DFF_806/Q_reg  ( .Q(WX5829), .CLK(CK), .DIN(WX5828) );
  dffs1 \DFF_805/Q_reg  ( .Q(WX5827), .CLK(CK), .DIN(WX5826) );
  dffs1 \DFF_804/Q_reg  ( .Q(WX5825), .CLK(CK), .DIN(WX5824) );
  dffs1 \DFF_803/Q_reg  ( .Q(WX5823), .CLK(CK), .DIN(WX5822) );
  dffs1 \DFF_802/Q_reg  ( .Q(WX5821), .CLK(CK), .DIN(WX5820) );
  dffs1 \DFF_801/Q_reg  ( .Q(WX5819), .CLK(CK), .DIN(WX5818) );
  dffs1 \DFF_800/Q_reg  ( .Q(WX5817), .CLK(CK), .DIN(WX5816) );
  dffs1 \DFF_799/Q_reg  ( .Q(WX5719), .CLK(CK), .DIN(WX5718) );
  dffs1 \DFF_798/Q_reg  ( .Q(WX5717), .CLK(CK), .DIN(WX5716) );
  dffs1 \DFF_797/Q_reg  ( .Q(WX5715), .CLK(CK), .DIN(WX5714) );
  dffs1 \DFF_796/Q_reg  ( .Q(WX5713), .CLK(CK), .DIN(WX5712) );
  dffs1 \DFF_795/Q_reg  ( .Q(WX5711), .CLK(CK), .DIN(WX5710) );
  dffs1 \DFF_794/Q_reg  ( .Q(WX5709), .CLK(CK), .DIN(WX5708) );
  dffs1 \DFF_793/Q_reg  ( .Q(WX5707), .CLK(CK), .DIN(WX5706) );
  dffs1 \DFF_792/Q_reg  ( .Q(WX5705), .CLK(CK), .DIN(WX5704) );
  dffs1 \DFF_791/Q_reg  ( .Q(WX5703), .CLK(CK), .DIN(WX5702) );
  dffs1 \DFF_790/Q_reg  ( .Q(WX5701), .CLK(CK), .DIN(WX5700) );
  dffs1 \DFF_789/Q_reg  ( .Q(WX5699), .CLK(CK), .DIN(WX5698) );
  dffs1 \DFF_788/Q_reg  ( .Q(WX5697), .CLK(CK), .DIN(WX5696) );
  dffs1 \DFF_787/Q_reg  ( .Q(WX5695), .CLK(CK), .DIN(WX5694) );
  dffs1 \DFF_786/Q_reg  ( .Q(WX5693), .CLK(CK), .DIN(WX5692) );
  dffs1 \DFF_785/Q_reg  ( .Q(WX5691), .CLK(CK), .DIN(WX5690) );
  dffs1 \DFF_784/Q_reg  ( .Q(WX5689), .CLK(CK), .DIN(WX5688) );
  dffs1 \DFF_783/Q_reg  ( .Q(WX5687), .CLK(CK), .DIN(WX5686) );
  dffs1 \DFF_782/Q_reg  ( .Q(WX5685), .CLK(CK), .DIN(WX5684) );
  dffs1 \DFF_781/Q_reg  ( .Q(WX5683), .CLK(CK), .DIN(WX5682) );
  dffs1 \DFF_780/Q_reg  ( .Q(WX5681), .CLK(CK), .DIN(WX5680) );
  dffs1 \DFF_779/Q_reg  ( .Q(WX5679), .CLK(CK), .DIN(WX5678) );
  dffs1 \DFF_778/Q_reg  ( .Q(WX5677), .CLK(CK), .DIN(WX5676) );
  dffs1 \DFF_777/Q_reg  ( .Q(WX5675), .CLK(CK), .DIN(WX5674) );
  dffs1 \DFF_776/Q_reg  ( .Q(WX5673), .CLK(CK), .DIN(WX5672) );
  dffs1 \DFF_775/Q_reg  ( .Q(WX5671), .CLK(CK), .DIN(WX5670) );
  dffs1 \DFF_774/Q_reg  ( .Q(WX5669), .CLK(CK), .DIN(WX5668) );
  dffs1 \DFF_773/Q_reg  ( .Q(WX5667), .CLK(CK), .DIN(WX5666) );
  dffs1 \DFF_772/Q_reg  ( .Q(WX5665), .CLK(CK), .DIN(WX5664) );
  dffs1 \DFF_771/Q_reg  ( .Q(WX5663), .CLK(CK), .DIN(WX5662) );
  dffs1 \DFF_770/Q_reg  ( .Q(WX5661), .CLK(CK), .DIN(WX5660) );
  dffs1 \DFF_769/Q_reg  ( .Q(WX5659), .CLK(CK), .DIN(WX5658) );
  dffs1 \DFF_768/Q_reg  ( .Q(WX5657), .CLK(CK), .DIN(WX5656) );
  dffs1 \DFF_767/Q_reg  ( .Q(CRC_OUT_6_31), .CLK(CK), .DIN(WX5205) );
  dffs1 \DFF_766/Q_reg  ( .Q(CRC_OUT_6_30), .CLK(CK), .DIN(WX5203) );
  dffs1 \DFF_765/Q_reg  ( .Q(CRC_OUT_6_29), .CLK(CK), .DIN(WX5201) );
  dffs1 \DFF_764/Q_reg  ( .Q(CRC_OUT_6_28), .CLK(CK), .DIN(WX5199) );
  dffs1 \DFF_763/Q_reg  ( .Q(CRC_OUT_6_27), .CLK(CK), .DIN(WX5197) );
  dffs1 \DFF_762/Q_reg  ( .Q(CRC_OUT_6_26), .CLK(CK), .DIN(WX5195) );
  dffs1 \DFF_761/Q_reg  ( .Q(CRC_OUT_6_25), .CLK(CK), .DIN(WX5193) );
  dffs1 \DFF_760/Q_reg  ( .Q(CRC_OUT_6_24), .CLK(CK), .DIN(WX5191) );
  dffs1 \DFF_759/Q_reg  ( .Q(CRC_OUT_6_23), .CLK(CK), .DIN(WX5189) );
  dffs1 \DFF_758/Q_reg  ( .Q(CRC_OUT_6_22), .CLK(CK), .DIN(WX5187) );
  dffs1 \DFF_757/Q_reg  ( .Q(CRC_OUT_6_21), .CLK(CK), .DIN(WX5185) );
  dffs1 \DFF_756/Q_reg  ( .Q(CRC_OUT_6_20), .CLK(CK), .DIN(WX5183) );
  dffs1 \DFF_755/Q_reg  ( .Q(CRC_OUT_6_19), .CLK(CK), .DIN(WX5181) );
  dffs1 \DFF_754/Q_reg  ( .Q(CRC_OUT_6_18), .CLK(CK), .DIN(WX5179) );
  dffs1 \DFF_753/Q_reg  ( .Q(CRC_OUT_6_17), .CLK(CK), .DIN(WX5177) );
  dffs1 \DFF_752/Q_reg  ( .Q(CRC_OUT_6_16), .CLK(CK), .DIN(WX5175) );
  dffs1 \DFF_751/Q_reg  ( .Q(CRC_OUT_6_15), .CLK(CK), .DIN(WX5173) );
  dffs1 \DFF_750/Q_reg  ( .Q(CRC_OUT_6_14), .CLK(CK), .DIN(WX5171) );
  dffs1 \DFF_749/Q_reg  ( .Q(CRC_OUT_6_13), .CLK(CK), .DIN(WX5169) );
  dffs1 \DFF_748/Q_reg  ( .Q(CRC_OUT_6_12), .CLK(CK), .DIN(WX5167) );
  dffs1 \DFF_747/Q_reg  ( .Q(CRC_OUT_6_11), .CLK(CK), .DIN(WX5165) );
  dffs1 \DFF_746/Q_reg  ( .Q(CRC_OUT_6_10), .CLK(CK), .DIN(WX5163) );
  dffs1 \DFF_745/Q_reg  ( .Q(CRC_OUT_6_9), .CLK(CK), .DIN(WX5161) );
  dffs1 \DFF_744/Q_reg  ( .Q(CRC_OUT_6_8), .CLK(CK), .DIN(WX5159) );
  dffs1 \DFF_743/Q_reg  ( .Q(CRC_OUT_6_7), .CLK(CK), .DIN(WX5157) );
  dffs1 \DFF_742/Q_reg  ( .Q(CRC_OUT_6_6), .CLK(CK), .DIN(WX5155) );
  dffs1 \DFF_741/Q_reg  ( .Q(CRC_OUT_6_5), .CLK(CK), .DIN(WX5153) );
  dffs1 \DFF_740/Q_reg  ( .Q(CRC_OUT_6_4), .CLK(CK), .DIN(WX5151) );
  dffs1 \DFF_739/Q_reg  ( .Q(CRC_OUT_6_3), .CLK(CK), .DIN(WX5149) );
  dffs1 \DFF_738/Q_reg  ( .Q(CRC_OUT_6_2), .CLK(CK), .DIN(WX5147) );
  dffs1 \DFF_737/Q_reg  ( .Q(CRC_OUT_6_1), .CLK(CK), .DIN(WX5145) );
  dffs1 \DFF_736/Q_reg  ( .Q(CRC_OUT_6_0), .CLK(CK), .DIN(WX5143) );
  dffs1 \DFF_735/Q_reg  ( .QN(n3269), .Q(WX4778), .CLK(CK), .DIN(WX4777) );
  dffs1 \DFF_734/Q_reg  ( .QN(n3270), .Q(WX4776), .CLK(CK), .DIN(WX4775) );
  dffs1 \DFF_733/Q_reg  ( .QN(n3271), .Q(WX4774), .CLK(CK), .DIN(WX4773) );
  dffs1 \DFF_732/Q_reg  ( .QN(n3272), .Q(WX4772), .CLK(CK), .DIN(WX4771) );
  dffs1 \DFF_731/Q_reg  ( .QN(n3273), .Q(WX4770), .CLK(CK), .DIN(WX4769) );
  dffs1 \DFF_730/Q_reg  ( .QN(n3274), .Q(WX4768), .CLK(CK), .DIN(WX4767) );
  dffs1 \DFF_729/Q_reg  ( .QN(n3275), .Q(WX4766), .CLK(CK), .DIN(WX4765) );
  dffs1 \DFF_728/Q_reg  ( .QN(n3276), .Q(WX4764), .CLK(CK), .DIN(WX4763) );
  dffs1 \DFF_727/Q_reg  ( .QN(n3277), .Q(WX4762), .CLK(CK), .DIN(WX4761) );
  dffs1 \DFF_726/Q_reg  ( .QN(n3278), .Q(WX4760), .CLK(CK), .DIN(WX4759) );
  dffs1 \DFF_725/Q_reg  ( .QN(n3279), .Q(WX4758), .CLK(CK), .DIN(WX4757) );
  dffs1 \DFF_724/Q_reg  ( .QN(n3280), .Q(WX4756), .CLK(CK), .DIN(WX4755) );
  dffs1 \DFF_723/Q_reg  ( .QN(n3281), .Q(WX4754), .CLK(CK), .DIN(WX4753) );
  dffs1 \DFF_722/Q_reg  ( .QN(n3282), .Q(WX4752), .CLK(CK), .DIN(WX4751) );
  dffs1 \DFF_721/Q_reg  ( .QN(n3283), .Q(WX4750), .CLK(CK), .DIN(WX4749) );
  dffs1 \DFF_720/Q_reg  ( .QN(n3284), .Q(WX4748), .CLK(CK), .DIN(WX4747) );
  dffs1 \DFF_719/Q_reg  ( .Q(WX4746), .CLK(CK), .DIN(WX4745) );
  dffs1 \DFF_718/Q_reg  ( .Q(WX4744), .CLK(CK), .DIN(WX4743) );
  dffs1 \DFF_717/Q_reg  ( .Q(WX4742), .CLK(CK), .DIN(WX4741) );
  dffs1 \DFF_716/Q_reg  ( .Q(WX4740), .CLK(CK), .DIN(WX4739) );
  dffs1 \DFF_715/Q_reg  ( .Q(WX4738), .CLK(CK), .DIN(WX4737) );
  dffs1 \DFF_714/Q_reg  ( .Q(WX4736), .CLK(CK), .DIN(WX4735) );
  dffs1 \DFF_713/Q_reg  ( .Q(WX4734), .CLK(CK), .DIN(WX4733) );
  dffs1 \DFF_712/Q_reg  ( .Q(WX4732), .CLK(CK), .DIN(WX4731) );
  dffs1 \DFF_711/Q_reg  ( .Q(WX4730), .CLK(CK), .DIN(WX4729) );
  dffs1 \DFF_710/Q_reg  ( .Q(WX4728), .CLK(CK), .DIN(WX4727) );
  dffs1 \DFF_709/Q_reg  ( .Q(WX4726), .CLK(CK), .DIN(WX4725) );
  dffs1 \DFF_708/Q_reg  ( .Q(WX4724), .CLK(CK), .DIN(WX4723) );
  dffs1 \DFF_707/Q_reg  ( .Q(WX4722), .CLK(CK), .DIN(WX4721) );
  dffs1 \DFF_706/Q_reg  ( .Q(WX4720), .CLK(CK), .DIN(WX4719) );
  dffs1 \DFF_705/Q_reg  ( .Q(WX4718), .CLK(CK), .DIN(WX4717) );
  dffs1 \DFF_704/Q_reg  ( .Q(WX4716), .CLK(CK), .DIN(WX4715) );
  dffs1 \DFF_703/Q_reg  ( .Q(WX4714), .CLK(CK), .DIN(WX4713) );
  dffs1 \DFF_702/Q_reg  ( .Q(WX4712), .CLK(CK), .DIN(WX4711) );
  dffs1 \DFF_701/Q_reg  ( .Q(WX4710), .CLK(CK), .DIN(WX4709) );
  dffs1 \DFF_700/Q_reg  ( .Q(WX4708), .CLK(CK), .DIN(WX4707) );
  dffs1 \DFF_699/Q_reg  ( .Q(WX4706), .CLK(CK), .DIN(WX4705) );
  dffs1 \DFF_698/Q_reg  ( .Q(WX4704), .CLK(CK), .DIN(WX4703) );
  dffs1 \DFF_697/Q_reg  ( .Q(WX4702), .CLK(CK), .DIN(WX4701) );
  dffs1 \DFF_696/Q_reg  ( .Q(WX4700), .CLK(CK), .DIN(WX4699) );
  dffs1 \DFF_695/Q_reg  ( .Q(WX4698), .CLK(CK), .DIN(WX4697) );
  dffs1 \DFF_694/Q_reg  ( .Q(WX4696), .CLK(CK), .DIN(WX4695) );
  dffs1 \DFF_693/Q_reg  ( .Q(WX4694), .CLK(CK), .DIN(WX4693) );
  dffs1 \DFF_692/Q_reg  ( .Q(WX4692), .CLK(CK), .DIN(WX4691) );
  dffs1 \DFF_691/Q_reg  ( .Q(WX4690), .CLK(CK), .DIN(WX4689) );
  dffs1 \DFF_690/Q_reg  ( .Q(WX4688), .CLK(CK), .DIN(WX4687) );
  dffs1 \DFF_689/Q_reg  ( .Q(WX4686), .CLK(CK), .DIN(WX4685) );
  dffs1 \DFF_688/Q_reg  ( .Q(WX4684), .CLK(CK), .DIN(WX4683) );
  dffs1 \DFF_687/Q_reg  ( .Q(WX4682), .CLK(CK), .DIN(WX4681) );
  dffs1 \DFF_686/Q_reg  ( .Q(WX4680), .CLK(CK), .DIN(WX4679) );
  dffs1 \DFF_685/Q_reg  ( .Q(WX4678), .CLK(CK), .DIN(WX4677) );
  dffs1 \DFF_684/Q_reg  ( .Q(WX4676), .CLK(CK), .DIN(WX4675) );
  dffs1 \DFF_683/Q_reg  ( .Q(WX4674), .CLK(CK), .DIN(WX4673) );
  dffs1 \DFF_682/Q_reg  ( .Q(WX4672), .CLK(CK), .DIN(WX4671) );
  dffs1 \DFF_681/Q_reg  ( .Q(WX4670), .CLK(CK), .DIN(WX4669) );
  dffs1 \DFF_680/Q_reg  ( .Q(WX4668), .CLK(CK), .DIN(WX4667) );
  dffs1 \DFF_679/Q_reg  ( .Q(WX4666), .CLK(CK), .DIN(WX4665) );
  dffs1 \DFF_678/Q_reg  ( .Q(WX4664), .CLK(CK), .DIN(WX4663) );
  dffs1 \DFF_677/Q_reg  ( .Q(WX4662), .CLK(CK), .DIN(WX4661) );
  dffs1 \DFF_676/Q_reg  ( .Q(WX4660), .CLK(CK), .DIN(WX4659) );
  dffs1 \DFF_675/Q_reg  ( .Q(WX4658), .CLK(CK), .DIN(WX4657) );
  dffs1 \DFF_674/Q_reg  ( .Q(WX4656), .CLK(CK), .DIN(WX4655) );
  dffs1 \DFF_673/Q_reg  ( .Q(WX4654), .CLK(CK), .DIN(WX4653) );
  dffs1 \DFF_672/Q_reg  ( .Q(WX4652), .CLK(CK), .DIN(WX4651) );
  dffs1 \DFF_671/Q_reg  ( .Q(WX4650), .CLK(CK), .DIN(WX4649) );
  dffs1 \DFF_670/Q_reg  ( .Q(WX4648), .CLK(CK), .DIN(WX4647) );
  dffs1 \DFF_669/Q_reg  ( .Q(WX4646), .CLK(CK), .DIN(WX4645) );
  dffs1 \DFF_668/Q_reg  ( .Q(WX4644), .CLK(CK), .DIN(WX4643) );
  dffs1 \DFF_667/Q_reg  ( .Q(WX4642), .CLK(CK), .DIN(WX4641) );
  dffs1 \DFF_666/Q_reg  ( .Q(WX4640), .CLK(CK), .DIN(WX4639) );
  dffs1 \DFF_665/Q_reg  ( .Q(WX4638), .CLK(CK), .DIN(WX4637) );
  dffs1 \DFF_664/Q_reg  ( .Q(WX4636), .CLK(CK), .DIN(WX4635) );
  dffs1 \DFF_663/Q_reg  ( .Q(WX4634), .CLK(CK), .DIN(WX4633) );
  dffs1 \DFF_662/Q_reg  ( .Q(WX4632), .CLK(CK), .DIN(WX4631) );
  dffs1 \DFF_661/Q_reg  ( .Q(WX4630), .CLK(CK), .DIN(WX4629) );
  dffs1 \DFF_660/Q_reg  ( .Q(WX4628), .CLK(CK), .DIN(WX4627) );
  dffs1 \DFF_659/Q_reg  ( .Q(WX4626), .CLK(CK), .DIN(WX4625) );
  dffs1 \DFF_658/Q_reg  ( .Q(WX4624), .CLK(CK), .DIN(WX4623) );
  dffs1 \DFF_657/Q_reg  ( .Q(WX4622), .CLK(CK), .DIN(WX4621) );
  dffs1 \DFF_656/Q_reg  ( .Q(WX4620), .CLK(CK), .DIN(WX4619) );
  dffs1 \DFF_655/Q_reg  ( .QN(n3013), .CLK(CK), .DIN(WX4617) );
  dffs1 \DFF_654/Q_reg  ( .QN(n3014), .CLK(CK), .DIN(WX4615) );
  dffs1 \DFF_653/Q_reg  ( .QN(n3015), .CLK(CK), .DIN(WX4613) );
  dffs1 \DFF_652/Q_reg  ( .QN(n3016), .CLK(CK), .DIN(WX4611) );
  dffs1 \DFF_651/Q_reg  ( .QN(n3017), .CLK(CK), .DIN(WX4609) );
  dffs1 \DFF_650/Q_reg  ( .QN(n3018), .CLK(CK), .DIN(WX4607) );
  dffs1 \DFF_649/Q_reg  ( .QN(n3019), .CLK(CK), .DIN(WX4605) );
  dffs1 \DFF_648/Q_reg  ( .QN(n3020), .CLK(CK), .DIN(WX4603) );
  dffs1 \DFF_647/Q_reg  ( .QN(n3021), .CLK(CK), .DIN(WX4601) );
  dffs1 \DFF_646/Q_reg  ( .QN(n3022), .CLK(CK), .DIN(WX4599) );
  dffs1 \DFF_645/Q_reg  ( .QN(n3023), .CLK(CK), .DIN(WX4597) );
  dffs1 \DFF_644/Q_reg  ( .QN(n3024), .CLK(CK), .DIN(WX4595) );
  dffs1 \DFF_643/Q_reg  ( .QN(n3025), .CLK(CK), .DIN(WX4593) );
  dffs1 \DFF_642/Q_reg  ( .QN(n3026), .CLK(CK), .DIN(WX4591) );
  dffs1 \DFF_641/Q_reg  ( .QN(n3027), .CLK(CK), .DIN(WX4589) );
  dffs1 \DFF_640/Q_reg  ( .QN(n3028), .CLK(CK), .DIN(WX4587) );
  dffs1 \DFF_639/Q_reg  ( .QN(n3173), .CLK(CK), .DIN(WX4585) );
  dffs1 \DFF_638/Q_reg  ( .QN(n3174), .CLK(CK), .DIN(WX4583) );
  dffs1 \DFF_637/Q_reg  ( .QN(n3175), .CLK(CK), .DIN(WX4581) );
  dffs1 \DFF_636/Q_reg  ( .QN(n3176), .CLK(CK), .DIN(WX4579) );
  dffs1 \DFF_635/Q_reg  ( .QN(n3177), .CLK(CK), .DIN(WX4577) );
  dffs1 \DFF_634/Q_reg  ( .QN(n3178), .CLK(CK), .DIN(WX4575) );
  dffs1 \DFF_633/Q_reg  ( .QN(n3179), .CLK(CK), .DIN(WX4573) );
  dffs1 \DFF_632/Q_reg  ( .QN(n3180), .CLK(CK), .DIN(WX4571) );
  dffs1 \DFF_631/Q_reg  ( .QN(n3181), .CLK(CK), .DIN(WX4569) );
  dffs1 \DFF_630/Q_reg  ( .QN(n3182), .CLK(CK), .DIN(WX4567) );
  dffs1 \DFF_629/Q_reg  ( .QN(n3183), .CLK(CK), .DIN(WX4565) );
  dffs1 \DFF_628/Q_reg  ( .QN(n3184), .CLK(CK), .DIN(WX4563) );
  dffs1 \DFF_627/Q_reg  ( .QN(n3185), .CLK(CK), .DIN(WX4561) );
  dffs1 \DFF_626/Q_reg  ( .QN(n3186), .CLK(CK), .DIN(WX4559) );
  dffs1 \DFF_625/Q_reg  ( .QN(n3187), .CLK(CK), .DIN(WX4557) );
  dffs1 \DFF_624/Q_reg  ( .QN(n3188), .CLK(CK), .DIN(WX4555) );
  dffs1 \DFF_623/Q_reg  ( .Q(WX4554), .CLK(CK), .DIN(WX4553) );
  dffs1 \DFF_622/Q_reg  ( .Q(WX4552), .CLK(CK), .DIN(WX4551) );
  dffs1 \DFF_621/Q_reg  ( .Q(WX4550), .CLK(CK), .DIN(WX4549) );
  dffs1 \DFF_620/Q_reg  ( .Q(WX4548), .CLK(CK), .DIN(WX4547) );
  dffs1 \DFF_619/Q_reg  ( .Q(WX4546), .CLK(CK), .DIN(WX4545) );
  dffs1 \DFF_618/Q_reg  ( .Q(WX4544), .CLK(CK), .DIN(WX4543) );
  dffs1 \DFF_617/Q_reg  ( .Q(WX4542), .CLK(CK), .DIN(WX4541) );
  dffs1 \DFF_616/Q_reg  ( .Q(WX4540), .CLK(CK), .DIN(WX4539) );
  dffs1 \DFF_615/Q_reg  ( .Q(WX4538), .CLK(CK), .DIN(WX4537) );
  dffs1 \DFF_614/Q_reg  ( .Q(WX4536), .CLK(CK), .DIN(WX4535) );
  dffs1 \DFF_613/Q_reg  ( .Q(WX4534), .CLK(CK), .DIN(WX4533) );
  dffs1 \DFF_612/Q_reg  ( .Q(WX4532), .CLK(CK), .DIN(WX4531) );
  dffs1 \DFF_611/Q_reg  ( .Q(WX4530), .CLK(CK), .DIN(WX4529) );
  dffs1 \DFF_610/Q_reg  ( .Q(WX4528), .CLK(CK), .DIN(WX4527) );
  dffs1 \DFF_609/Q_reg  ( .Q(WX4526), .CLK(CK), .DIN(WX4525) );
  dffs1 \DFF_608/Q_reg  ( .Q(WX4524), .CLK(CK), .DIN(WX4523) );
  dffs1 \DFF_607/Q_reg  ( .Q(WX4426), .CLK(CK), .DIN(WX4425) );
  dffs1 \DFF_606/Q_reg  ( .Q(WX4424), .CLK(CK), .DIN(WX4423) );
  dffs1 \DFF_605/Q_reg  ( .Q(WX4422), .CLK(CK), .DIN(WX4421) );
  dffs1 \DFF_604/Q_reg  ( .Q(WX4420), .CLK(CK), .DIN(WX4419) );
  dffs1 \DFF_603/Q_reg  ( .Q(WX4418), .CLK(CK), .DIN(WX4417) );
  dffs1 \DFF_602/Q_reg  ( .Q(WX4416), .CLK(CK), .DIN(WX4415) );
  dffs1 \DFF_601/Q_reg  ( .Q(WX4414), .CLK(CK), .DIN(WX4413) );
  dffs1 \DFF_600/Q_reg  ( .Q(WX4412), .CLK(CK), .DIN(WX4411) );
  dffs1 \DFF_599/Q_reg  ( .Q(WX4410), .CLK(CK), .DIN(WX4409) );
  dffs1 \DFF_598/Q_reg  ( .Q(WX4408), .CLK(CK), .DIN(WX4407) );
  dffs1 \DFF_597/Q_reg  ( .Q(WX4406), .CLK(CK), .DIN(WX4405) );
  dffs1 \DFF_596/Q_reg  ( .Q(WX4404), .CLK(CK), .DIN(WX4403) );
  dffs1 \DFF_595/Q_reg  ( .Q(WX4402), .CLK(CK), .DIN(WX4401) );
  dffs1 \DFF_594/Q_reg  ( .Q(WX4400), .CLK(CK), .DIN(WX4399) );
  dffs1 \DFF_593/Q_reg  ( .Q(WX4398), .CLK(CK), .DIN(WX4397) );
  dffs1 \DFF_592/Q_reg  ( .Q(WX4396), .CLK(CK), .DIN(WX4395) );
  dffs1 \DFF_591/Q_reg  ( .Q(WX4394), .CLK(CK), .DIN(WX4393) );
  dffs1 \DFF_590/Q_reg  ( .Q(WX4392), .CLK(CK), .DIN(WX4391) );
  dffs1 \DFF_589/Q_reg  ( .Q(WX4390), .CLK(CK), .DIN(WX4389) );
  dffs1 \DFF_588/Q_reg  ( .Q(WX4388), .CLK(CK), .DIN(WX4387) );
  dffs1 \DFF_587/Q_reg  ( .Q(WX4386), .CLK(CK), .DIN(WX4385) );
  dffs1 \DFF_586/Q_reg  ( .Q(WX4384), .CLK(CK), .DIN(WX4383) );
  dffs1 \DFF_585/Q_reg  ( .Q(WX4382), .CLK(CK), .DIN(WX4381) );
  dffs1 \DFF_584/Q_reg  ( .Q(WX4380), .CLK(CK), .DIN(WX4379) );
  dffs1 \DFF_583/Q_reg  ( .Q(WX4378), .CLK(CK), .DIN(WX4377) );
  dffs1 \DFF_582/Q_reg  ( .Q(WX4376), .CLK(CK), .DIN(WX4375) );
  dffs1 \DFF_581/Q_reg  ( .Q(WX4374), .CLK(CK), .DIN(WX4373) );
  dffs1 \DFF_580/Q_reg  ( .Q(WX4372), .CLK(CK), .DIN(WX4371) );
  dffs1 \DFF_579/Q_reg  ( .Q(WX4370), .CLK(CK), .DIN(WX4369) );
  dffs1 \DFF_578/Q_reg  ( .Q(WX4368), .CLK(CK), .DIN(WX4367) );
  dffs1 \DFF_577/Q_reg  ( .Q(WX4366), .CLK(CK), .DIN(WX4365) );
  dffs1 \DFF_576/Q_reg  ( .Q(WX4364), .CLK(CK), .DIN(WX4363) );
  dffs1 \DFF_575/Q_reg  ( .Q(CRC_OUT_7_31), .CLK(CK), .DIN(WX3912) );
  dffs1 \DFF_574/Q_reg  ( .Q(CRC_OUT_7_30), .CLK(CK), .DIN(WX3910) );
  dffs1 \DFF_573/Q_reg  ( .Q(CRC_OUT_7_29), .CLK(CK), .DIN(WX3908) );
  dffs1 \DFF_572/Q_reg  ( .Q(CRC_OUT_7_28), .CLK(CK), .DIN(WX3906) );
  dffs1 \DFF_571/Q_reg  ( .Q(CRC_OUT_7_27), .CLK(CK), .DIN(WX3904) );
  dffs1 \DFF_570/Q_reg  ( .Q(CRC_OUT_7_26), .CLK(CK), .DIN(WX3902) );
  dffs1 \DFF_569/Q_reg  ( .Q(CRC_OUT_7_25), .CLK(CK), .DIN(WX3900) );
  dffs1 \DFF_568/Q_reg  ( .Q(CRC_OUT_7_24), .CLK(CK), .DIN(WX3898) );
  dffs1 \DFF_567/Q_reg  ( .Q(CRC_OUT_7_23), .CLK(CK), .DIN(WX3896) );
  dffs1 \DFF_566/Q_reg  ( .Q(CRC_OUT_7_22), .CLK(CK), .DIN(WX3894) );
  dffs1 \DFF_565/Q_reg  ( .Q(CRC_OUT_7_21), .CLK(CK), .DIN(WX3892) );
  dffs1 \DFF_564/Q_reg  ( .Q(CRC_OUT_7_20), .CLK(CK), .DIN(WX3890) );
  dffs1 \DFF_563/Q_reg  ( .Q(CRC_OUT_7_19), .CLK(CK), .DIN(WX3888) );
  dffs1 \DFF_562/Q_reg  ( .Q(CRC_OUT_7_18), .CLK(CK), .DIN(WX3886) );
  dffs1 \DFF_561/Q_reg  ( .Q(CRC_OUT_7_17), .CLK(CK), .DIN(WX3884) );
  dffs1 \DFF_560/Q_reg  ( .Q(CRC_OUT_7_16), .CLK(CK), .DIN(WX3882) );
  dffs1 \DFF_559/Q_reg  ( .Q(CRC_OUT_7_15), .CLK(CK), .DIN(WX3880) );
  dffs1 \DFF_558/Q_reg  ( .Q(CRC_OUT_7_14), .CLK(CK), .DIN(WX3878) );
  dffs1 \DFF_557/Q_reg  ( .Q(CRC_OUT_7_13), .CLK(CK), .DIN(WX3876) );
  dffs1 \DFF_556/Q_reg  ( .Q(CRC_OUT_7_12), .CLK(CK), .DIN(WX3874) );
  dffs1 \DFF_555/Q_reg  ( .Q(CRC_OUT_7_11), .CLK(CK), .DIN(WX3872) );
  dffs1 \DFF_554/Q_reg  ( .Q(CRC_OUT_7_10), .CLK(CK), .DIN(WX3870) );
  dffs1 \DFF_553/Q_reg  ( .Q(CRC_OUT_7_9), .CLK(CK), .DIN(WX3868) );
  dffs1 \DFF_552/Q_reg  ( .Q(CRC_OUT_7_8), .CLK(CK), .DIN(WX3866) );
  dffs1 \DFF_551/Q_reg  ( .Q(CRC_OUT_7_7), .CLK(CK), .DIN(WX3864) );
  dffs1 \DFF_550/Q_reg  ( .Q(CRC_OUT_7_6), .CLK(CK), .DIN(WX3862) );
  dffs1 \DFF_549/Q_reg  ( .Q(CRC_OUT_7_5), .CLK(CK), .DIN(WX3860) );
  dffs1 \DFF_548/Q_reg  ( .Q(CRC_OUT_7_4), .CLK(CK), .DIN(WX3858) );
  dffs1 \DFF_547/Q_reg  ( .Q(CRC_OUT_7_3), .CLK(CK), .DIN(WX3856) );
  dffs1 \DFF_546/Q_reg  ( .Q(CRC_OUT_7_2), .CLK(CK), .DIN(WX3854) );
  dffs1 \DFF_545/Q_reg  ( .Q(CRC_OUT_7_1), .CLK(CK), .DIN(WX3852) );
  dffs1 \DFF_544/Q_reg  ( .Q(CRC_OUT_7_0), .CLK(CK), .DIN(WX3850) );
  dffs1 \DFF_543/Q_reg  ( .QN(n3285), .Q(WX3485), .CLK(CK), .DIN(WX3484) );
  dffs1 \DFF_542/Q_reg  ( .QN(n3287), .Q(WX3483), .CLK(CK), .DIN(WX3482) );
  dffs1 \DFF_541/Q_reg  ( .QN(n3289), .Q(WX3481), .CLK(CK), .DIN(WX3480) );
  dffs1 \DFF_540/Q_reg  ( .QN(n3291), .Q(WX3479), .CLK(CK), .DIN(WX3478) );
  dffs1 \DFF_539/Q_reg  ( .QN(n3293), .Q(WX3477), .CLK(CK), .DIN(WX3476) );
  dffs1 \DFF_538/Q_reg  ( .QN(n3295), .Q(WX3475), .CLK(CK), .DIN(WX3474) );
  dffs1 \DFF_537/Q_reg  ( .QN(n3297), .Q(WX3473), .CLK(CK), .DIN(WX3472) );
  dffs1 \DFF_536/Q_reg  ( .QN(n3299), .Q(WX3471), .CLK(CK), .DIN(WX3470) );
  dffs1 \DFF_535/Q_reg  ( .QN(n3301), .Q(WX3469), .CLK(CK), .DIN(WX3468) );
  dffs1 \DFF_534/Q_reg  ( .QN(n3303), .Q(WX3467), .CLK(CK), .DIN(WX3466) );
  dffs1 \DFF_533/Q_reg  ( .QN(n3305), .Q(WX3465), .CLK(CK), .DIN(WX3464) );
  dffs1 \DFF_532/Q_reg  ( .QN(n3307), .Q(WX3463), .CLK(CK), .DIN(WX3462) );
  dffs1 \DFF_531/Q_reg  ( .QN(n3309), .Q(WX3461), .CLK(CK), .DIN(WX3460) );
  dffs1 \DFF_530/Q_reg  ( .QN(n3311), .Q(WX3459), .CLK(CK), .DIN(WX3458) );
  dffs1 \DFF_529/Q_reg  ( .QN(n3313), .Q(WX3457), .CLK(CK), .DIN(WX3456) );
  dffs1 \DFF_528/Q_reg  ( .QN(n3315), .Q(WX3455), .CLK(CK), .DIN(WX3454) );
  dffs1 \DFF_527/Q_reg  ( .Q(WX3453), .CLK(CK), .DIN(WX3452) );
  dffs1 \DFF_526/Q_reg  ( .Q(WX3451), .CLK(CK), .DIN(WX3450) );
  dffs1 \DFF_525/Q_reg  ( .Q(WX3449), .CLK(CK), .DIN(WX3448) );
  dffs1 \DFF_524/Q_reg  ( .Q(WX3447), .CLK(CK), .DIN(WX3446) );
  dffs1 \DFF_523/Q_reg  ( .Q(WX3445), .CLK(CK), .DIN(WX3444) );
  dffs1 \DFF_522/Q_reg  ( .Q(WX3443), .CLK(CK), .DIN(WX3442) );
  dffs1 \DFF_521/Q_reg  ( .Q(WX3441), .CLK(CK), .DIN(WX3440) );
  dffs1 \DFF_520/Q_reg  ( .Q(WX3439), .CLK(CK), .DIN(WX3438) );
  dffs1 \DFF_519/Q_reg  ( .Q(WX3437), .CLK(CK), .DIN(WX3436) );
  dffs1 \DFF_518/Q_reg  ( .Q(WX3435), .CLK(CK), .DIN(WX3434) );
  dffs1 \DFF_517/Q_reg  ( .Q(WX3433), .CLK(CK), .DIN(WX3432) );
  dffs1 \DFF_516/Q_reg  ( .Q(WX3431), .CLK(CK), .DIN(WX3430) );
  dffs1 \DFF_515/Q_reg  ( .Q(WX3429), .CLK(CK), .DIN(WX3428) );
  dffs1 \DFF_514/Q_reg  ( .Q(WX3427), .CLK(CK), .DIN(WX3426) );
  dffs1 \DFF_513/Q_reg  ( .Q(WX3425), .CLK(CK), .DIN(WX3424) );
  dffs1 \DFF_512/Q_reg  ( .Q(WX3423), .CLK(CK), .DIN(WX3422) );
  dffs1 \DFF_511/Q_reg  ( .Q(WX3421), .CLK(CK), .DIN(WX3420) );
  dffs1 \DFF_510/Q_reg  ( .Q(WX3419), .CLK(CK), .DIN(WX3418) );
  dffs1 \DFF_509/Q_reg  ( .Q(WX3417), .CLK(CK), .DIN(WX3416) );
  dffs1 \DFF_508/Q_reg  ( .Q(WX3415), .CLK(CK), .DIN(WX3414) );
  dffs1 \DFF_507/Q_reg  ( .Q(WX3413), .CLK(CK), .DIN(WX3412) );
  dffs1 \DFF_506/Q_reg  ( .Q(WX3411), .CLK(CK), .DIN(WX3410) );
  dffs1 \DFF_505/Q_reg  ( .Q(WX3409), .CLK(CK), .DIN(WX3408) );
  dffs1 \DFF_504/Q_reg  ( .Q(WX3407), .CLK(CK), .DIN(WX3406) );
  dffs1 \DFF_503/Q_reg  ( .Q(WX3405), .CLK(CK), .DIN(WX3404) );
  dffs1 \DFF_502/Q_reg  ( .Q(WX3403), .CLK(CK), .DIN(WX3402) );
  dffs1 \DFF_501/Q_reg  ( .Q(WX3401), .CLK(CK), .DIN(WX3400) );
  dffs1 \DFF_500/Q_reg  ( .Q(WX3399), .CLK(CK), .DIN(WX3398) );
  dffs1 \DFF_499/Q_reg  ( .Q(WX3397), .CLK(CK), .DIN(WX3396) );
  dffs1 \DFF_498/Q_reg  ( .Q(WX3395), .CLK(CK), .DIN(WX3394) );
  dffs1 \DFF_497/Q_reg  ( .Q(WX3393), .CLK(CK), .DIN(WX3392) );
  dffs1 \DFF_496/Q_reg  ( .Q(WX3391), .CLK(CK), .DIN(WX3390) );
  dffs1 \DFF_495/Q_reg  ( .Q(WX3389), .CLK(CK), .DIN(WX3388) );
  dffs1 \DFF_494/Q_reg  ( .Q(WX3387), .CLK(CK), .DIN(WX3386) );
  dffs1 \DFF_493/Q_reg  ( .Q(WX3385), .CLK(CK), .DIN(WX3384) );
  dffs1 \DFF_492/Q_reg  ( .Q(WX3383), .CLK(CK), .DIN(WX3382) );
  dffs1 \DFF_491/Q_reg  ( .Q(WX3381), .CLK(CK), .DIN(WX3380) );
  dffs1 \DFF_490/Q_reg  ( .Q(WX3379), .CLK(CK), .DIN(WX3378) );
  dffs1 \DFF_489/Q_reg  ( .Q(WX3377), .CLK(CK), .DIN(WX3376) );
  dffs1 \DFF_488/Q_reg  ( .Q(WX3375), .CLK(CK), .DIN(WX3374) );
  dffs1 \DFF_487/Q_reg  ( .Q(WX3373), .CLK(CK), .DIN(WX3372) );
  dffs1 \DFF_486/Q_reg  ( .Q(WX3371), .CLK(CK), .DIN(WX3370) );
  dffs1 \DFF_485/Q_reg  ( .Q(WX3369), .CLK(CK), .DIN(WX3368) );
  dffs1 \DFF_484/Q_reg  ( .Q(WX3367), .CLK(CK), .DIN(WX3366) );
  dffs1 \DFF_483/Q_reg  ( .Q(WX3365), .CLK(CK), .DIN(WX3364) );
  dffs1 \DFF_482/Q_reg  ( .Q(WX3363), .CLK(CK), .DIN(WX3362) );
  dffs1 \DFF_481/Q_reg  ( .Q(WX3361), .CLK(CK), .DIN(WX3360) );
  dffs1 \DFF_480/Q_reg  ( .Q(WX3359), .CLK(CK), .DIN(WX3358) );
  dffs1 \DFF_479/Q_reg  ( .Q(WX3357), .CLK(CK), .DIN(WX3356) );
  dffs1 \DFF_478/Q_reg  ( .Q(WX3355), .CLK(CK), .DIN(WX3354) );
  dffs1 \DFF_477/Q_reg  ( .Q(WX3353), .CLK(CK), .DIN(WX3352) );
  dffs1 \DFF_476/Q_reg  ( .Q(WX3351), .CLK(CK), .DIN(WX3350) );
  dffs1 \DFF_475/Q_reg  ( .Q(WX3349), .CLK(CK), .DIN(WX3348) );
  dffs1 \DFF_474/Q_reg  ( .Q(WX3347), .CLK(CK), .DIN(WX3346) );
  dffs1 \DFF_473/Q_reg  ( .Q(WX3345), .CLK(CK), .DIN(WX3344) );
  dffs1 \DFF_472/Q_reg  ( .Q(WX3343), .CLK(CK), .DIN(WX3342) );
  dffs1 \DFF_471/Q_reg  ( .Q(WX3341), .CLK(CK), .DIN(WX3340) );
  dffs1 \DFF_470/Q_reg  ( .Q(WX3339), .CLK(CK), .DIN(WX3338) );
  dffs1 \DFF_469/Q_reg  ( .Q(WX3337), .CLK(CK), .DIN(WX3336) );
  dffs1 \DFF_468/Q_reg  ( .Q(WX3335), .CLK(CK), .DIN(WX3334) );
  dffs1 \DFF_467/Q_reg  ( .Q(WX3333), .CLK(CK), .DIN(WX3332) );
  dffs1 \DFF_466/Q_reg  ( .Q(WX3331), .CLK(CK), .DIN(WX3330) );
  dffs1 \DFF_465/Q_reg  ( .Q(WX3329), .CLK(CK), .DIN(WX3328) );
  dffs1 \DFF_464/Q_reg  ( .Q(WX3327), .CLK(CK), .DIN(WX3326) );
  dffs1 \DFF_463/Q_reg  ( .QN(n3045), .CLK(CK), .DIN(WX3324) );
  dffs1 \DFF_462/Q_reg  ( .QN(n3047), .CLK(CK), .DIN(WX3322) );
  dffs1 \DFF_461/Q_reg  ( .QN(n3049), .CLK(CK), .DIN(WX3320) );
  dffs1 \DFF_460/Q_reg  ( .QN(n3051), .CLK(CK), .DIN(WX3318) );
  dffs1 \DFF_459/Q_reg  ( .QN(n3053), .CLK(CK), .DIN(WX3316) );
  dffs1 \DFF_458/Q_reg  ( .QN(n3055), .CLK(CK), .DIN(WX3314) );
  dffs1 \DFF_457/Q_reg  ( .QN(n3057), .CLK(CK), .DIN(WX3312) );
  dffs1 \DFF_456/Q_reg  ( .QN(n3059), .CLK(CK), .DIN(WX3310) );
  dffs1 \DFF_455/Q_reg  ( .QN(n3061), .CLK(CK), .DIN(WX3308) );
  dffs1 \DFF_454/Q_reg  ( .QN(n3063), .CLK(CK), .DIN(WX3306) );
  dffs1 \DFF_453/Q_reg  ( .QN(n3065), .CLK(CK), .DIN(WX3304) );
  dffs1 \DFF_452/Q_reg  ( .QN(n3067), .CLK(CK), .DIN(WX3302) );
  dffs1 \DFF_451/Q_reg  ( .QN(n3069), .CLK(CK), .DIN(WX3300) );
  dffs1 \DFF_450/Q_reg  ( .QN(n3071), .CLK(CK), .DIN(WX3298) );
  dffs1 \DFF_449/Q_reg  ( .QN(n3073), .CLK(CK), .DIN(WX3296) );
  dffs1 \DFF_448/Q_reg  ( .QN(n3075), .CLK(CK), .DIN(WX3294) );
  dffs1 \DFF_447/Q_reg  ( .QN(n3189), .CLK(CK), .DIN(WX3292) );
  dffs1 \DFF_446/Q_reg  ( .QN(n3190), .CLK(CK), .DIN(WX3290) );
  dffs1 \DFF_445/Q_reg  ( .QN(n3191), .CLK(CK), .DIN(WX3288) );
  dffs1 \DFF_444/Q_reg  ( .QN(n3192), .CLK(CK), .DIN(WX3286) );
  dffs1 \DFF_443/Q_reg  ( .QN(n3193), .CLK(CK), .DIN(WX3284) );
  dffs1 \DFF_442/Q_reg  ( .QN(n3194), .CLK(CK), .DIN(WX3282) );
  dffs1 \DFF_441/Q_reg  ( .QN(n3195), .CLK(CK), .DIN(WX3280) );
  dffs1 \DFF_440/Q_reg  ( .QN(n3196), .CLK(CK), .DIN(WX3278) );
  dffs1 \DFF_439/Q_reg  ( .QN(n3197), .CLK(CK), .DIN(WX3276) );
  dffs1 \DFF_438/Q_reg  ( .QN(n3198), .CLK(CK), .DIN(WX3274) );
  dffs1 \DFF_437/Q_reg  ( .QN(n3199), .CLK(CK), .DIN(WX3272) );
  dffs1 \DFF_436/Q_reg  ( .QN(n3200), .CLK(CK), .DIN(WX3270) );
  dffs1 \DFF_435/Q_reg  ( .QN(n3201), .CLK(CK), .DIN(WX3268) );
  dffs1 \DFF_434/Q_reg  ( .QN(n3202), .CLK(CK), .DIN(WX3266) );
  dffs1 \DFF_433/Q_reg  ( .QN(n3203), .CLK(CK), .DIN(WX3264) );
  dffs1 \DFF_432/Q_reg  ( .QN(n3204), .CLK(CK), .DIN(WX3262) );
  dffs1 \DFF_431/Q_reg  ( .Q(WX3261), .CLK(CK), .DIN(WX3260) );
  dffs1 \DFF_430/Q_reg  ( .Q(WX3259), .CLK(CK), .DIN(WX3258) );
  dffs1 \DFF_429/Q_reg  ( .Q(WX3257), .CLK(CK), .DIN(WX3256) );
  dffs1 \DFF_428/Q_reg  ( .Q(WX3255), .CLK(CK), .DIN(WX3254) );
  dffs1 \DFF_427/Q_reg  ( .Q(WX3253), .CLK(CK), .DIN(WX3252) );
  dffs1 \DFF_426/Q_reg  ( .Q(WX3251), .CLK(CK), .DIN(WX3250) );
  dffs1 \DFF_425/Q_reg  ( .Q(WX3249), .CLK(CK), .DIN(WX3248) );
  dffs1 \DFF_424/Q_reg  ( .Q(WX3247), .CLK(CK), .DIN(WX3246) );
  dffs1 \DFF_423/Q_reg  ( .Q(WX3245), .CLK(CK), .DIN(WX3244) );
  dffs1 \DFF_422/Q_reg  ( .Q(WX3243), .CLK(CK), .DIN(WX3242) );
  dffs1 \DFF_421/Q_reg  ( .Q(WX3241), .CLK(CK), .DIN(WX3240) );
  dffs1 \DFF_420/Q_reg  ( .Q(WX3239), .CLK(CK), .DIN(WX3238) );
  dffs1 \DFF_419/Q_reg  ( .Q(WX3237), .CLK(CK), .DIN(WX3236) );
  dffs1 \DFF_418/Q_reg  ( .Q(WX3235), .CLK(CK), .DIN(WX3234) );
  dffs1 \DFF_417/Q_reg  ( .Q(WX3233), .CLK(CK), .DIN(WX3232) );
  dffs1 \DFF_416/Q_reg  ( .Q(WX3231), .CLK(CK), .DIN(WX3230) );
  dffs1 \DFF_415/Q_reg  ( .Q(WX3133), .CLK(CK), .DIN(WX3132) );
  dffs1 \DFF_414/Q_reg  ( .Q(WX3131), .CLK(CK), .DIN(WX3130) );
  dffs1 \DFF_413/Q_reg  ( .Q(WX3129), .CLK(CK), .DIN(WX3128) );
  dffs1 \DFF_412/Q_reg  ( .Q(WX3127), .CLK(CK), .DIN(WX3126) );
  dffs1 \DFF_411/Q_reg  ( .Q(WX3125), .CLK(CK), .DIN(WX3124) );
  dffs1 \DFF_410/Q_reg  ( .Q(WX3123), .CLK(CK), .DIN(WX3122) );
  dffs1 \DFF_409/Q_reg  ( .Q(WX3121), .CLK(CK), .DIN(WX3120) );
  dffs1 \DFF_408/Q_reg  ( .Q(WX3119), .CLK(CK), .DIN(WX3118) );
  dffs1 \DFF_407/Q_reg  ( .Q(WX3117), .CLK(CK), .DIN(WX3116) );
  dffs1 \DFF_406/Q_reg  ( .Q(WX3115), .CLK(CK), .DIN(WX3114) );
  dffs1 \DFF_405/Q_reg  ( .Q(WX3113), .CLK(CK), .DIN(WX3112) );
  dffs1 \DFF_404/Q_reg  ( .Q(WX3111), .CLK(CK), .DIN(WX3110) );
  dffs1 \DFF_403/Q_reg  ( .Q(WX3109), .CLK(CK), .DIN(WX3108) );
  dffs1 \DFF_402/Q_reg  ( .Q(WX3107), .CLK(CK), .DIN(WX3106) );
  dffs1 \DFF_401/Q_reg  ( .Q(WX3105), .CLK(CK), .DIN(WX3104) );
  dffs1 \DFF_400/Q_reg  ( .Q(WX3103), .CLK(CK), .DIN(WX3102) );
  dffs1 \DFF_399/Q_reg  ( .Q(WX3101), .CLK(CK), .DIN(WX3100) );
  dffs1 \DFF_398/Q_reg  ( .Q(WX3099), .CLK(CK), .DIN(WX3098) );
  dffs1 \DFF_397/Q_reg  ( .Q(WX3097), .CLK(CK), .DIN(WX3096) );
  dffs1 \DFF_396/Q_reg  ( .Q(WX3095), .CLK(CK), .DIN(WX3094) );
  dffs1 \DFF_395/Q_reg  ( .Q(WX3093), .CLK(CK), .DIN(WX3092) );
  dffs1 \DFF_394/Q_reg  ( .Q(WX3091), .CLK(CK), .DIN(WX3090) );
  dffs1 \DFF_393/Q_reg  ( .Q(WX3089), .CLK(CK), .DIN(WX3088) );
  dffs1 \DFF_392/Q_reg  ( .Q(WX3087), .CLK(CK), .DIN(WX3086) );
  dffs1 \DFF_391/Q_reg  ( .Q(WX3085), .CLK(CK), .DIN(WX3084) );
  dffs1 \DFF_390/Q_reg  ( .Q(WX3083), .CLK(CK), .DIN(WX3082) );
  dffs1 \DFF_389/Q_reg  ( .Q(WX3081), .CLK(CK), .DIN(WX3080) );
  dffs1 \DFF_388/Q_reg  ( .Q(WX3079), .CLK(CK), .DIN(WX3078) );
  dffs1 \DFF_387/Q_reg  ( .Q(WX3077), .CLK(CK), .DIN(WX3076) );
  dffs1 \DFF_386/Q_reg  ( .Q(WX3075), .CLK(CK), .DIN(WX3074) );
  dffs1 \DFF_385/Q_reg  ( .Q(WX3073), .CLK(CK), .DIN(WX3072) );
  dffs1 \DFF_384/Q_reg  ( .Q(WX3071), .CLK(CK), .DIN(WX3070) );
  dffs1 \DFF_383/Q_reg  ( .Q(CRC_OUT_8_31), .CLK(CK), .DIN(WX2619) );
  dffs1 \DFF_382/Q_reg  ( .Q(CRC_OUT_8_30), .CLK(CK), .DIN(WX2617) );
  dffs1 \DFF_381/Q_reg  ( .Q(CRC_OUT_8_29), .CLK(CK), .DIN(WX2615) );
  dffs1 \DFF_380/Q_reg  ( .Q(CRC_OUT_8_28), .CLK(CK), .DIN(WX2613) );
  dffs1 \DFF_379/Q_reg  ( .Q(CRC_OUT_8_27), .CLK(CK), .DIN(WX2611) );
  dffs1 \DFF_378/Q_reg  ( .Q(CRC_OUT_8_26), .CLK(CK), .DIN(WX2609) );
  dffs1 \DFF_377/Q_reg  ( .Q(CRC_OUT_8_25), .CLK(CK), .DIN(WX2607) );
  dffs1 \DFF_376/Q_reg  ( .Q(CRC_OUT_8_24), .CLK(CK), .DIN(WX2605) );
  dffs1 \DFF_375/Q_reg  ( .Q(CRC_OUT_8_23), .CLK(CK), .DIN(WX2603) );
  dffs1 \DFF_374/Q_reg  ( .Q(CRC_OUT_8_22), .CLK(CK), .DIN(WX2601) );
  dffs1 \DFF_373/Q_reg  ( .Q(CRC_OUT_8_21), .CLK(CK), .DIN(WX2599) );
  dffs1 \DFF_372/Q_reg  ( .Q(CRC_OUT_8_20), .CLK(CK), .DIN(WX2597) );
  dffs1 \DFF_371/Q_reg  ( .Q(CRC_OUT_8_19), .CLK(CK), .DIN(WX2595) );
  dffs1 \DFF_370/Q_reg  ( .Q(CRC_OUT_8_18), .CLK(CK), .DIN(WX2593) );
  dffs1 \DFF_369/Q_reg  ( .Q(CRC_OUT_8_17), .CLK(CK), .DIN(WX2591) );
  dffs1 \DFF_368/Q_reg  ( .Q(CRC_OUT_8_16), .CLK(CK), .DIN(WX2589) );
  dffs1 \DFF_367/Q_reg  ( .Q(CRC_OUT_8_15), .CLK(CK), .DIN(WX2587) );
  dffs1 \DFF_366/Q_reg  ( .Q(CRC_OUT_8_14), .CLK(CK), .DIN(WX2585) );
  dffs1 \DFF_365/Q_reg  ( .Q(CRC_OUT_8_13), .CLK(CK), .DIN(WX2583) );
  dffs1 \DFF_364/Q_reg  ( .Q(CRC_OUT_8_12), .CLK(CK), .DIN(WX2581) );
  dffs1 \DFF_363/Q_reg  ( .Q(CRC_OUT_8_11), .CLK(CK), .DIN(WX2579) );
  dffs1 \DFF_362/Q_reg  ( .Q(CRC_OUT_8_10), .CLK(CK), .DIN(WX2577) );
  dffs1 \DFF_361/Q_reg  ( .Q(CRC_OUT_8_9), .CLK(CK), .DIN(WX2575) );
  dffs1 \DFF_360/Q_reg  ( .Q(CRC_OUT_8_8), .CLK(CK), .DIN(WX2573) );
  dffs1 \DFF_359/Q_reg  ( .Q(CRC_OUT_8_7), .CLK(CK), .DIN(WX2571) );
  dffs1 \DFF_358/Q_reg  ( .Q(CRC_OUT_8_6), .CLK(CK), .DIN(WX2569) );
  dffs1 \DFF_357/Q_reg  ( .Q(CRC_OUT_8_5), .CLK(CK), .DIN(WX2567) );
  dffs1 \DFF_356/Q_reg  ( .Q(CRC_OUT_8_4), .CLK(CK), .DIN(WX2565) );
  dffs1 \DFF_355/Q_reg  ( .Q(CRC_OUT_8_3), .CLK(CK), .DIN(WX2563) );
  dffs1 \DFF_354/Q_reg  ( .Q(CRC_OUT_8_2), .CLK(CK), .DIN(WX2561) );
  dffs1 \DFF_353/Q_reg  ( .Q(CRC_OUT_8_1), .CLK(CK), .DIN(WX2559) );
  dffs1 \DFF_352/Q_reg  ( .Q(CRC_OUT_8_0), .CLK(CK), .DIN(WX2557) );
  dffs1 \DFF_351/Q_reg  ( .QN(n3286), .Q(WX2192), .CLK(CK), .DIN(WX2191) );
  dffs1 \DFF_350/Q_reg  ( .QN(n3288), .Q(WX2190), .CLK(CK), .DIN(WX2189) );
  dffs1 \DFF_349/Q_reg  ( .QN(n3290), .Q(WX2188), .CLK(CK), .DIN(WX2187) );
  dffs1 \DFF_348/Q_reg  ( .QN(n3292), .Q(WX2186), .CLK(CK), .DIN(WX2185) );
  dffs1 \DFF_347/Q_reg  ( .QN(n3294), .Q(WX2184), .CLK(CK), .DIN(WX2183) );
  dffs1 \DFF_346/Q_reg  ( .QN(n3296), .Q(WX2182), .CLK(CK), .DIN(WX2181) );
  dffs1 \DFF_345/Q_reg  ( .QN(n3298), .Q(WX2180), .CLK(CK), .DIN(WX2179) );
  dffs1 \DFF_344/Q_reg  ( .QN(n3300), .Q(WX2178), .CLK(CK), .DIN(WX2177) );
  dffs1 \DFF_343/Q_reg  ( .QN(n3302), .Q(WX2176), .CLK(CK), .DIN(WX2175) );
  dffs1 \DFF_342/Q_reg  ( .QN(n3304), .Q(WX2174), .CLK(CK), .DIN(WX2173) );
  dffs1 \DFF_341/Q_reg  ( .QN(n3306), .Q(WX2172), .CLK(CK), .DIN(WX2171) );
  dffs1 \DFF_340/Q_reg  ( .QN(n3308), .Q(WX2170), .CLK(CK), .DIN(WX2169) );
  dffs1 \DFF_339/Q_reg  ( .QN(n3310), .Q(WX2168), .CLK(CK), .DIN(WX2167) );
  dffs1 \DFF_338/Q_reg  ( .QN(n3312), .Q(WX2166), .CLK(CK), .DIN(WX2165) );
  dffs1 \DFF_337/Q_reg  ( .QN(n3314), .Q(WX2164), .CLK(CK), .DIN(WX2163) );
  dffs1 \DFF_336/Q_reg  ( .QN(n3316), .Q(WX2162), .CLK(CK), .DIN(WX2161) );
  dffs1 \DFF_335/Q_reg  ( .Q(WX2160), .CLK(CK), .DIN(WX2159) );
  dffs1 \DFF_334/Q_reg  ( .Q(WX2158), .CLK(CK), .DIN(WX2157) );
  dffs1 \DFF_333/Q_reg  ( .Q(WX2156), .CLK(CK), .DIN(WX2155) );
  dffs1 \DFF_332/Q_reg  ( .Q(WX2154), .CLK(CK), .DIN(WX2153) );
  dffs1 \DFF_331/Q_reg  ( .Q(WX2152), .CLK(CK), .DIN(WX2151) );
  dffs1 \DFF_330/Q_reg  ( .Q(WX2150), .CLK(CK), .DIN(WX2149) );
  dffs1 \DFF_329/Q_reg  ( .Q(WX2148), .CLK(CK), .DIN(WX2147) );
  dffs1 \DFF_328/Q_reg  ( .Q(WX2146), .CLK(CK), .DIN(WX2145) );
  dffs1 \DFF_327/Q_reg  ( .Q(WX2144), .CLK(CK), .DIN(WX2143) );
  dffs1 \DFF_326/Q_reg  ( .Q(WX2142), .CLK(CK), .DIN(WX2141) );
  dffs1 \DFF_325/Q_reg  ( .Q(WX2140), .CLK(CK), .DIN(WX2139) );
  dffs1 \DFF_324/Q_reg  ( .Q(WX2138), .CLK(CK), .DIN(WX2137) );
  dffs1 \DFF_323/Q_reg  ( .Q(WX2136), .CLK(CK), .DIN(WX2135) );
  dffs1 \DFF_322/Q_reg  ( .Q(WX2134), .CLK(CK), .DIN(WX2133) );
  dffs1 \DFF_321/Q_reg  ( .Q(WX2132), .CLK(CK), .DIN(WX2131) );
  dffs1 \DFF_320/Q_reg  ( .Q(WX2130), .CLK(CK), .DIN(WX2129) );
  dffs1 \DFF_319/Q_reg  ( .Q(WX2128), .CLK(CK), .DIN(WX2127) );
  dffs1 \DFF_318/Q_reg  ( .Q(WX2126), .CLK(CK), .DIN(WX2125) );
  dffs1 \DFF_317/Q_reg  ( .Q(WX2124), .CLK(CK), .DIN(WX2123) );
  dffs1 \DFF_316/Q_reg  ( .Q(WX2122), .CLK(CK), .DIN(WX2121) );
  dffs1 \DFF_315/Q_reg  ( .Q(WX2120), .CLK(CK), .DIN(WX2119) );
  dffs1 \DFF_314/Q_reg  ( .Q(WX2118), .CLK(CK), .DIN(WX2117) );
  dffs1 \DFF_313/Q_reg  ( .Q(WX2116), .CLK(CK), .DIN(WX2115) );
  dffs1 \DFF_312/Q_reg  ( .Q(WX2114), .CLK(CK), .DIN(WX2113) );
  dffs1 \DFF_311/Q_reg  ( .Q(WX2112), .CLK(CK), .DIN(WX2111) );
  dffs1 \DFF_310/Q_reg  ( .Q(WX2110), .CLK(CK), .DIN(WX2109) );
  dffs1 \DFF_309/Q_reg  ( .Q(WX2108), .CLK(CK), .DIN(WX2107) );
  dffs1 \DFF_308/Q_reg  ( .Q(WX2106), .CLK(CK), .DIN(WX2105) );
  dffs1 \DFF_307/Q_reg  ( .Q(WX2104), .CLK(CK), .DIN(WX2103) );
  dffs1 \DFF_306/Q_reg  ( .Q(WX2102), .CLK(CK), .DIN(WX2101) );
  dffs1 \DFF_305/Q_reg  ( .Q(WX2100), .CLK(CK), .DIN(WX2099) );
  dffs1 \DFF_304/Q_reg  ( .Q(WX2098), .CLK(CK), .DIN(WX2097) );
  dffs1 \DFF_303/Q_reg  ( .Q(WX2096), .CLK(CK), .DIN(WX2095) );
  dffs1 \DFF_302/Q_reg  ( .Q(WX2094), .CLK(CK), .DIN(WX2093) );
  dffs1 \DFF_301/Q_reg  ( .Q(WX2092), .CLK(CK), .DIN(WX2091) );
  dffs1 \DFF_300/Q_reg  ( .Q(WX2090), .CLK(CK), .DIN(WX2089) );
  dffs1 \DFF_299/Q_reg  ( .Q(WX2088), .CLK(CK), .DIN(WX2087) );
  dffs1 \DFF_298/Q_reg  ( .Q(WX2086), .CLK(CK), .DIN(WX2085) );
  dffs1 \DFF_297/Q_reg  ( .Q(WX2084), .CLK(CK), .DIN(WX2083) );
  dffs1 \DFF_296/Q_reg  ( .Q(WX2082), .CLK(CK), .DIN(WX2081) );
  dffs1 \DFF_295/Q_reg  ( .Q(WX2080), .CLK(CK), .DIN(WX2079) );
  dffs1 \DFF_294/Q_reg  ( .Q(WX2078), .CLK(CK), .DIN(WX2077) );
  dffs1 \DFF_293/Q_reg  ( .Q(WX2076), .CLK(CK), .DIN(WX2075) );
  dffs1 \DFF_292/Q_reg  ( .Q(WX2074), .CLK(CK), .DIN(WX2073) );
  dffs1 \DFF_291/Q_reg  ( .Q(WX2072), .CLK(CK), .DIN(WX2071) );
  dffs1 \DFF_290/Q_reg  ( .Q(WX2070), .CLK(CK), .DIN(WX2069) );
  dffs1 \DFF_289/Q_reg  ( .Q(WX2068), .CLK(CK), .DIN(WX2067) );
  dffs1 \DFF_288/Q_reg  ( .Q(WX2066), .CLK(CK), .DIN(WX2065) );
  dffs1 \DFF_287/Q_reg  ( .QN(n3029), .CLK(CK), .DIN(WX2063) );
  dffs1 \DFF_286/Q_reg  ( .QN(n3030), .CLK(CK), .DIN(WX2061) );
  dffs1 \DFF_285/Q_reg  ( .QN(n3031), .CLK(CK), .DIN(WX2059) );
  dffs1 \DFF_284/Q_reg  ( .QN(n3032), .CLK(CK), .DIN(WX2057) );
  dffs1 \DFF_283/Q_reg  ( .QN(n3033), .CLK(CK), .DIN(WX2055) );
  dffs1 \DFF_282/Q_reg  ( .QN(n3034), .CLK(CK), .DIN(WX2053) );
  dffs1 \DFF_281/Q_reg  ( .QN(n3035), .CLK(CK), .DIN(WX2051) );
  dffs1 \DFF_280/Q_reg  ( .QN(n3036), .CLK(CK), .DIN(WX2049) );
  dffs1 \DFF_279/Q_reg  ( .QN(n3037), .CLK(CK), .DIN(WX2047) );
  dffs1 \DFF_278/Q_reg  ( .QN(n3038), .CLK(CK), .DIN(WX2045) );
  dffs1 \DFF_277/Q_reg  ( .QN(n3039), .CLK(CK), .DIN(WX2043) );
  dffs1 \DFF_276/Q_reg  ( .QN(n3040), .CLK(CK), .DIN(WX2041) );
  dffs1 \DFF_275/Q_reg  ( .QN(n3041), .CLK(CK), .DIN(WX2039) );
  dffs1 \DFF_274/Q_reg  ( .QN(n3042), .CLK(CK), .DIN(WX2037) );
  dffs1 \DFF_273/Q_reg  ( .QN(n3043), .CLK(CK), .DIN(WX2035) );
  dffs1 \DFF_272/Q_reg  ( .QN(n3044), .CLK(CK), .DIN(WX2033) );
  dffs1 \DFF_271/Q_reg  ( .QN(n3046), .CLK(CK), .DIN(WX2031) );
  dffs1 \DFF_270/Q_reg  ( .QN(n3048), .CLK(CK), .DIN(WX2029) );
  dffs1 \DFF_269/Q_reg  ( .QN(n3050), .CLK(CK), .DIN(WX2027) );
  dffs1 \DFF_268/Q_reg  ( .QN(n3052), .CLK(CK), .DIN(WX2025) );
  dffs1 \DFF_267/Q_reg  ( .QN(n3054), .CLK(CK), .DIN(WX2023) );
  dffs1 \DFF_266/Q_reg  ( .QN(n3056), .CLK(CK), .DIN(WX2021) );
  dffs1 \DFF_265/Q_reg  ( .QN(n3058), .CLK(CK), .DIN(WX2019) );
  dffs1 \DFF_264/Q_reg  ( .QN(n3060), .CLK(CK), .DIN(WX2017) );
  dffs1 \DFF_263/Q_reg  ( .QN(n3062), .CLK(CK), .DIN(WX2015) );
  dffs1 \DFF_262/Q_reg  ( .QN(n3064), .CLK(CK), .DIN(WX2013) );
  dffs1 \DFF_261/Q_reg  ( .QN(n3066), .CLK(CK), .DIN(WX2011) );
  dffs1 \DFF_260/Q_reg  ( .QN(n3068), .CLK(CK), .DIN(WX2009) );
  dffs1 \DFF_259/Q_reg  ( .QN(n3070), .CLK(CK), .DIN(WX2007) );
  dffs1 \DFF_258/Q_reg  ( .QN(n3072), .CLK(CK), .DIN(WX2005) );
  dffs1 \DFF_257/Q_reg  ( .QN(n3074), .CLK(CK), .DIN(WX2003) );
  dffs1 \DFF_256/Q_reg  ( .QN(n3076), .CLK(CK), .DIN(WX2001) );
  dffs1 \DFF_255/Q_reg  ( .Q(WX2000), .CLK(CK), .DIN(WX1999) );
  dffs1 \DFF_254/Q_reg  ( .Q(WX1998), .CLK(CK), .DIN(WX1997) );
  dffs1 \DFF_253/Q_reg  ( .Q(WX1996), .CLK(CK), .DIN(WX1995) );
  dffs1 \DFF_252/Q_reg  ( .Q(WX1994), .CLK(CK), .DIN(WX1993) );
  dffs1 \DFF_251/Q_reg  ( .Q(WX1992), .CLK(CK), .DIN(WX1991) );
  dffs1 \DFF_250/Q_reg  ( .Q(WX1990), .CLK(CK), .DIN(WX1989) );
  dffs1 \DFF_249/Q_reg  ( .Q(WX1988), .CLK(CK), .DIN(WX1987) );
  dffs1 \DFF_248/Q_reg  ( .Q(WX1986), .CLK(CK), .DIN(WX1985) );
  dffs1 \DFF_247/Q_reg  ( .Q(WX1984), .CLK(CK), .DIN(WX1983) );
  dffs1 \DFF_246/Q_reg  ( .Q(WX1982), .CLK(CK), .DIN(WX1981) );
  dffs1 \DFF_245/Q_reg  ( .Q(WX1980), .CLK(CK), .DIN(WX1979) );
  dffs1 \DFF_244/Q_reg  ( .Q(WX1978), .CLK(CK), .DIN(WX1977) );
  dffs1 \DFF_243/Q_reg  ( .Q(WX1976), .CLK(CK), .DIN(WX1975) );
  dffs1 \DFF_242/Q_reg  ( .Q(WX1974), .CLK(CK), .DIN(WX1973) );
  dffs1 \DFF_241/Q_reg  ( .Q(WX1972), .CLK(CK), .DIN(WX1971) );
  dffs1 \DFF_240/Q_reg  ( .Q(WX1970), .CLK(CK), .DIN(WX1969) );
  dffs1 \DFF_239/Q_reg  ( .Q(WX1968), .CLK(CK), .DIN(WX1967) );
  dffs1 \DFF_238/Q_reg  ( .Q(WX1966), .CLK(CK), .DIN(WX1965) );
  dffs1 \DFF_237/Q_reg  ( .Q(WX1964), .CLK(CK), .DIN(WX1963) );
  dffs1 \DFF_236/Q_reg  ( .Q(WX1962), .CLK(CK), .DIN(WX1961) );
  dffs1 \DFF_235/Q_reg  ( .Q(WX1960), .CLK(CK), .DIN(WX1959) );
  dffs1 \DFF_234/Q_reg  ( .Q(WX1958), .CLK(CK), .DIN(WX1957) );
  dffs1 \DFF_233/Q_reg  ( .Q(WX1956), .CLK(CK), .DIN(WX1955) );
  dffs1 \DFF_232/Q_reg  ( .Q(WX1954), .CLK(CK), .DIN(WX1953) );
  dffs1 \DFF_231/Q_reg  ( .Q(WX1952), .CLK(CK), .DIN(WX1951) );
  dffs1 \DFF_230/Q_reg  ( .Q(WX1950), .CLK(CK), .DIN(WX1949) );
  dffs1 \DFF_229/Q_reg  ( .Q(WX1948), .CLK(CK), .DIN(WX1947) );
  dffs1 \DFF_228/Q_reg  ( .Q(WX1946), .CLK(CK), .DIN(WX1945) );
  dffs1 \DFF_227/Q_reg  ( .Q(WX1944), .CLK(CK), .DIN(WX1943) );
  dffs1 \DFF_226/Q_reg  ( .Q(WX1942), .CLK(CK), .DIN(WX1941) );
  dffs1 \DFF_225/Q_reg  ( .Q(WX1940), .CLK(CK), .DIN(WX1939) );
  dffs1 \DFF_224/Q_reg  ( .Q(WX1938), .CLK(CK), .DIN(WX1937) );
  dffs1 \DFF_223/Q_reg  ( .Q(WX1840), .CLK(CK), .DIN(WX1839) );
  dffs1 \DFF_222/Q_reg  ( .Q(WX1838), .CLK(CK), .DIN(WX1837) );
  dffs1 \DFF_221/Q_reg  ( .Q(WX1836), .CLK(CK), .DIN(WX1835) );
  dffs1 \DFF_220/Q_reg  ( .Q(WX1834), .CLK(CK), .DIN(WX1833) );
  dffs1 \DFF_219/Q_reg  ( .Q(WX1832), .CLK(CK), .DIN(WX1831) );
  dffs1 \DFF_218/Q_reg  ( .Q(WX1830), .CLK(CK), .DIN(WX1829) );
  dffs1 \DFF_217/Q_reg  ( .Q(WX1828), .CLK(CK), .DIN(WX1827) );
  dffs1 \DFF_216/Q_reg  ( .Q(WX1826), .CLK(CK), .DIN(WX1825) );
  dffs1 \DFF_215/Q_reg  ( .Q(WX1824), .CLK(CK), .DIN(WX1823) );
  dffs1 \DFF_214/Q_reg  ( .Q(WX1822), .CLK(CK), .DIN(WX1821) );
  dffs1 \DFF_213/Q_reg  ( .Q(WX1820), .CLK(CK), .DIN(WX1819) );
  dffs1 \DFF_212/Q_reg  ( .Q(WX1818), .CLK(CK), .DIN(WX1817) );
  dffs1 \DFF_211/Q_reg  ( .Q(WX1816), .CLK(CK), .DIN(WX1815) );
  dffs1 \DFF_210/Q_reg  ( .Q(WX1814), .CLK(CK), .DIN(WX1813) );
  dffs1 \DFF_209/Q_reg  ( .Q(WX1812), .CLK(CK), .DIN(WX1811) );
  dffs1 \DFF_208/Q_reg  ( .Q(WX1810), .CLK(CK), .DIN(WX1809) );
  dffs1 \DFF_207/Q_reg  ( .Q(WX1808), .CLK(CK), .DIN(WX1807) );
  dffs1 \DFF_206/Q_reg  ( .Q(WX1806), .CLK(CK), .DIN(WX1805) );
  dffs1 \DFF_205/Q_reg  ( .Q(WX1804), .CLK(CK), .DIN(WX1803) );
  dffs1 \DFF_204/Q_reg  ( .Q(WX1802), .CLK(CK), .DIN(WX1801) );
  dffs1 \DFF_203/Q_reg  ( .Q(WX1800), .CLK(CK), .DIN(WX1799) );
  dffs1 \DFF_202/Q_reg  ( .Q(WX1798), .CLK(CK), .DIN(WX1797) );
  dffs1 \DFF_201/Q_reg  ( .Q(WX1796), .CLK(CK), .DIN(WX1795) );
  dffs1 \DFF_200/Q_reg  ( .Q(WX1794), .CLK(CK), .DIN(WX1793) );
  dffs1 \DFF_199/Q_reg  ( .Q(WX1792), .CLK(CK), .DIN(WX1791) );
  dffs1 \DFF_198/Q_reg  ( .Q(WX1790), .CLK(CK), .DIN(WX1789) );
  dffs1 \DFF_197/Q_reg  ( .Q(WX1788), .CLK(CK), .DIN(WX1787) );
  dffs1 \DFF_196/Q_reg  ( .Q(WX1786), .CLK(CK), .DIN(WX1785) );
  dffs1 \DFF_195/Q_reg  ( .Q(WX1784), .CLK(CK), .DIN(WX1783) );
  dffs1 \DFF_194/Q_reg  ( .Q(WX1782), .CLK(CK), .DIN(WX1781) );
  dffs1 \DFF_193/Q_reg  ( .Q(WX1780), .CLK(CK), .DIN(WX1779) );
  dffs1 \DFF_192/Q_reg  ( .Q(WX1778), .CLK(CK), .DIN(WX1777) );
  dffs1 \DFF_191/Q_reg  ( .Q(CRC_OUT_9_31), .CLK(CK), .DIN(WX1326) );
  dffs1 \DFF_190/Q_reg  ( .Q(CRC_OUT_9_30), .CLK(CK), .DIN(WX1324) );
  dffs1 \DFF_189/Q_reg  ( .Q(CRC_OUT_9_29), .CLK(CK), .DIN(WX1322) );
  dffs1 \DFF_188/Q_reg  ( .Q(CRC_OUT_9_28), .CLK(CK), .DIN(WX1320) );
  dffs1 \DFF_187/Q_reg  ( .Q(CRC_OUT_9_27), .CLK(CK), .DIN(WX1318) );
  dffs1 \DFF_186/Q_reg  ( .Q(CRC_OUT_9_26), .CLK(CK), .DIN(WX1316) );
  dffs1 \DFF_185/Q_reg  ( .Q(CRC_OUT_9_25), .CLK(CK), .DIN(WX1314) );
  dffs1 \DFF_184/Q_reg  ( .Q(CRC_OUT_9_24), .CLK(CK), .DIN(WX1312) );
  dffs1 \DFF_183/Q_reg  ( .Q(CRC_OUT_9_23), .CLK(CK), .DIN(WX1310) );
  dffs1 \DFF_182/Q_reg  ( .Q(CRC_OUT_9_22), .CLK(CK), .DIN(WX1308) );
  dffs1 \DFF_181/Q_reg  ( .Q(CRC_OUT_9_21), .CLK(CK), .DIN(WX1306) );
  dffs1 \DFF_180/Q_reg  ( .Q(CRC_OUT_9_20), .CLK(CK), .DIN(WX1304) );
  dffs1 \DFF_179/Q_reg  ( .Q(CRC_OUT_9_19), .CLK(CK), .DIN(WX1302) );
  dffs1 \DFF_178/Q_reg  ( .Q(CRC_OUT_9_18), .CLK(CK), .DIN(WX1300) );
  dffs1 \DFF_177/Q_reg  ( .Q(CRC_OUT_9_17), .CLK(CK), .DIN(WX1298) );
  dffs1 \DFF_176/Q_reg  ( .Q(CRC_OUT_9_16), .CLK(CK), .DIN(WX1296) );
  dffs1 \DFF_175/Q_reg  ( .Q(CRC_OUT_9_15), .CLK(CK), .DIN(WX1294) );
  dffs1 \DFF_174/Q_reg  ( .Q(CRC_OUT_9_14), .CLK(CK), .DIN(WX1292) );
  dffs1 \DFF_173/Q_reg  ( .Q(CRC_OUT_9_13), .CLK(CK), .DIN(WX1290) );
  dffs1 \DFF_172/Q_reg  ( .Q(CRC_OUT_9_12), .CLK(CK), .DIN(WX1288) );
  dffs1 \DFF_171/Q_reg  ( .Q(CRC_OUT_9_11), .CLK(CK), .DIN(WX1286) );
  dffs1 \DFF_170/Q_reg  ( .Q(CRC_OUT_9_10), .CLK(CK), .DIN(WX1284) );
  dffs1 \DFF_169/Q_reg  ( .Q(CRC_OUT_9_9), .CLK(CK), .DIN(WX1282) );
  dffs1 \DFF_168/Q_reg  ( .Q(CRC_OUT_9_8), .CLK(CK), .DIN(WX1280) );
  dffs1 \DFF_167/Q_reg  ( .Q(CRC_OUT_9_7), .CLK(CK), .DIN(WX1278) );
  dffs1 \DFF_166/Q_reg  ( .Q(CRC_OUT_9_6), .CLK(CK), .DIN(WX1276) );
  dffs1 \DFF_165/Q_reg  ( .Q(CRC_OUT_9_5), .CLK(CK), .DIN(WX1274) );
  dffs1 \DFF_164/Q_reg  ( .Q(CRC_OUT_9_4), .CLK(CK), .DIN(WX1272) );
  dffs1 \DFF_163/Q_reg  ( .Q(CRC_OUT_9_3), .CLK(CK), .DIN(WX1270) );
  dffs1 \DFF_162/Q_reg  ( .Q(CRC_OUT_9_2), .CLK(CK), .DIN(WX1268) );
  dffs1 \DFF_161/Q_reg  ( .Q(CRC_OUT_9_1), .CLK(CK), .DIN(WX1266) );
  dffs1 \DFF_160/Q_reg  ( .Q(CRC_OUT_9_0), .CLK(CK), .DIN(WX1264) );
  dffs1 \DFF_159/Q_reg  ( .Q(WX899), .CLK(CK), .DIN(WX898) );
  dffs1 \DFF_158/Q_reg  ( .Q(WX897), .CLK(CK), .DIN(WX896) );
  dffs1 \DFF_157/Q_reg  ( .Q(WX895), .CLK(CK), .DIN(WX894) );
  dffs1 \DFF_156/Q_reg  ( .Q(WX893), .CLK(CK), .DIN(WX892) );
  dffs1 \DFF_155/Q_reg  ( .Q(WX891), .CLK(CK), .DIN(WX890) );
  dffs1 \DFF_154/Q_reg  ( .Q(WX889), .CLK(CK), .DIN(WX888) );
  dffs1 \DFF_153/Q_reg  ( .Q(WX887), .CLK(CK), .DIN(WX886) );
  dffs1 \DFF_152/Q_reg  ( .Q(WX885), .CLK(CK), .DIN(WX884) );
  dffs1 \DFF_151/Q_reg  ( .Q(WX883), .CLK(CK), .DIN(WX882) );
  dffs1 \DFF_150/Q_reg  ( .Q(WX881), .CLK(CK), .DIN(WX880) );
  dffs1 \DFF_149/Q_reg  ( .Q(WX879), .CLK(CK), .DIN(WX878) );
  dffs1 \DFF_148/Q_reg  ( .Q(WX877), .CLK(CK), .DIN(WX876) );
  dffs1 \DFF_147/Q_reg  ( .Q(WX875), .CLK(CK), .DIN(WX874) );
  dffs1 \DFF_146/Q_reg  ( .Q(WX873), .CLK(CK), .DIN(WX872) );
  dffs1 \DFF_145/Q_reg  ( .Q(WX871), .CLK(CK), .DIN(WX870) );
  dffs1 \DFF_144/Q_reg  ( .Q(WX869), .CLK(CK), .DIN(WX868) );
  dffs1 \DFF_143/Q_reg  ( .Q(WX867), .CLK(CK), .DIN(WX866) );
  dffs1 \DFF_142/Q_reg  ( .Q(WX865), .CLK(CK), .DIN(WX864) );
  dffs1 \DFF_141/Q_reg  ( .Q(WX863), .CLK(CK), .DIN(WX862) );
  dffs1 \DFF_140/Q_reg  ( .Q(WX861), .CLK(CK), .DIN(WX860) );
  dffs1 \DFF_139/Q_reg  ( .Q(WX859), .CLK(CK), .DIN(WX858) );
  dffs1 \DFF_138/Q_reg  ( .Q(WX857), .CLK(CK), .DIN(WX856) );
  dffs1 \DFF_137/Q_reg  ( .Q(WX855), .CLK(CK), .DIN(WX854) );
  dffs1 \DFF_136/Q_reg  ( .Q(WX853), .CLK(CK), .DIN(WX852) );
  dffs1 \DFF_135/Q_reg  ( .Q(WX851), .CLK(CK), .DIN(WX850) );
  dffs1 \DFF_134/Q_reg  ( .Q(WX849), .CLK(CK), .DIN(WX848) );
  dffs1 \DFF_133/Q_reg  ( .Q(WX847), .CLK(CK), .DIN(WX846) );
  dffs1 \DFF_132/Q_reg  ( .Q(WX845), .CLK(CK), .DIN(WX844) );
  dffs1 \DFF_131/Q_reg  ( .Q(WX843), .CLK(CK), .DIN(WX842) );
  dffs1 \DFF_130/Q_reg  ( .Q(WX841), .CLK(CK), .DIN(WX840) );
  dffs1 \DFF_129/Q_reg  ( .Q(WX839), .CLK(CK), .DIN(WX838) );
  dffs1 \DFF_128/Q_reg  ( .Q(WX837), .CLK(CK), .DIN(WX836) );
  dffs1 \DFF_127/Q_reg  ( .Q(WX835), .CLK(CK), .DIN(WX834) );
  dffs1 \DFF_126/Q_reg  ( .Q(WX833), .CLK(CK), .DIN(WX832) );
  dffs1 \DFF_125/Q_reg  ( .Q(WX831), .CLK(CK), .DIN(WX830) );
  dffs1 \DFF_124/Q_reg  ( .Q(WX829), .CLK(CK), .DIN(WX828) );
  dffs1 \DFF_123/Q_reg  ( .Q(WX827), .CLK(CK), .DIN(WX826) );
  dffs1 \DFF_122/Q_reg  ( .Q(WX825), .CLK(CK), .DIN(WX824) );
  dffs1 \DFF_121/Q_reg  ( .Q(WX823), .CLK(CK), .DIN(WX822) );
  dffs1 \DFF_120/Q_reg  ( .Q(WX821), .CLK(CK), .DIN(WX820) );
  dffs1 \DFF_119/Q_reg  ( .Q(WX819), .CLK(CK), .DIN(WX818) );
  dffs1 \DFF_118/Q_reg  ( .Q(WX817), .CLK(CK), .DIN(WX816) );
  dffs1 \DFF_117/Q_reg  ( .Q(WX815), .CLK(CK), .DIN(WX814) );
  dffs1 \DFF_116/Q_reg  ( .Q(WX813), .CLK(CK), .DIN(WX812) );
  dffs1 \DFF_115/Q_reg  ( .Q(WX811), .CLK(CK), .DIN(WX810) );
  dffs1 \DFF_114/Q_reg  ( .Q(WX809), .CLK(CK), .DIN(WX808) );
  dffs1 \DFF_113/Q_reg  ( .Q(WX807), .CLK(CK), .DIN(WX806) );
  dffs1 \DFF_112/Q_reg  ( .Q(WX805), .CLK(CK), .DIN(WX804) );
  dffs1 \DFF_111/Q_reg  ( .Q(WX803), .CLK(CK), .DIN(WX802) );
  dffs1 \DFF_110/Q_reg  ( .Q(WX801), .CLK(CK), .DIN(WX800) );
  dffs1 \DFF_109/Q_reg  ( .Q(WX799), .CLK(CK), .DIN(WX798) );
  dffs1 \DFF_108/Q_reg  ( .Q(WX797), .CLK(CK), .DIN(WX796) );
  dffs1 \DFF_107/Q_reg  ( .Q(WX795), .CLK(CK), .DIN(WX794) );
  dffs1 \DFF_106/Q_reg  ( .Q(WX793), .CLK(CK), .DIN(WX792) );
  dffs1 \DFF_105/Q_reg  ( .Q(WX791), .CLK(CK), .DIN(WX790) );
  dffs1 \DFF_104/Q_reg  ( .Q(WX789), .CLK(CK), .DIN(WX788) );
  dffs1 \DFF_103/Q_reg  ( .Q(WX787), .CLK(CK), .DIN(WX786) );
  dffs1 \DFF_102/Q_reg  ( .Q(WX785), .CLK(CK), .DIN(WX784) );
  dffs1 \DFF_101/Q_reg  ( .Q(WX783), .CLK(CK), .DIN(WX782) );
  dffs1 \DFF_100/Q_reg  ( .Q(WX781), .CLK(CK), .DIN(WX780) );
  dffs1 \DFF_99/Q_reg  ( .Q(WX779), .CLK(CK), .DIN(WX778) );
  dffs1 \DFF_98/Q_reg  ( .Q(WX777), .CLK(CK), .DIN(WX776) );
  dffs1 \DFF_97/Q_reg  ( .Q(WX775), .CLK(CK), .DIN(WX774) );
  dffs1 \DFF_96/Q_reg  ( .Q(WX773), .CLK(CK), .DIN(WX772) );
  dffs1 \DFF_95/Q_reg  ( .Q(WX771), .CLK(CK), .DIN(WX770) );
  dffs1 \DFF_94/Q_reg  ( .Q(WX769), .CLK(CK), .DIN(WX768) );
  dffs1 \DFF_93/Q_reg  ( .Q(WX767), .CLK(CK), .DIN(WX766) );
  dffs1 \DFF_92/Q_reg  ( .Q(WX765), .CLK(CK), .DIN(WX764) );
  dffs1 \DFF_91/Q_reg  ( .Q(WX763), .CLK(CK), .DIN(WX762) );
  dffs1 \DFF_90/Q_reg  ( .Q(WX761), .CLK(CK), .DIN(WX760) );
  dffs1 \DFF_89/Q_reg  ( .Q(WX759), .CLK(CK), .DIN(WX758) );
  dffs1 \DFF_88/Q_reg  ( .Q(WX757), .CLK(CK), .DIN(WX756) );
  dffs1 \DFF_87/Q_reg  ( .Q(WX755), .CLK(CK), .DIN(WX754) );
  dffs1 \DFF_86/Q_reg  ( .Q(WX753), .CLK(CK), .DIN(WX752) );
  dffs1 \DFF_85/Q_reg  ( .Q(WX751), .CLK(CK), .DIN(WX750) );
  dffs1 \DFF_84/Q_reg  ( .Q(WX749), .CLK(CK), .DIN(WX748) );
  dffs1 \DFF_83/Q_reg  ( .Q(WX747), .CLK(CK), .DIN(WX746) );
  dffs1 \DFF_82/Q_reg  ( .Q(WX745), .CLK(CK), .DIN(WX744) );
  dffs1 \DFF_81/Q_reg  ( .Q(WX743), .CLK(CK), .DIN(WX742) );
  dffs1 \DFF_80/Q_reg  ( .Q(WX741), .CLK(CK), .DIN(WX740) );
  dffs1 \DFF_79/Q_reg  ( .Q(WX739), .CLK(CK), .DIN(WX738) );
  dffs1 \DFF_78/Q_reg  ( .Q(WX737), .CLK(CK), .DIN(WX736) );
  dffs1 \DFF_77/Q_reg  ( .Q(WX735), .CLK(CK), .DIN(WX734) );
  dffs1 \DFF_76/Q_reg  ( .Q(WX733), .CLK(CK), .DIN(WX732) );
  dffs1 \DFF_75/Q_reg  ( .Q(WX731), .CLK(CK), .DIN(WX730) );
  dffs1 \DFF_74/Q_reg  ( .Q(WX729), .CLK(CK), .DIN(WX728) );
  dffs1 \DFF_73/Q_reg  ( .Q(WX727), .CLK(CK), .DIN(WX726) );
  dffs1 \DFF_72/Q_reg  ( .Q(WX725), .CLK(CK), .DIN(WX724) );
  dffs1 \DFF_71/Q_reg  ( .Q(WX723), .CLK(CK), .DIN(WX722) );
  dffs1 \DFF_70/Q_reg  ( .Q(WX721), .CLK(CK), .DIN(WX720) );
  dffs1 \DFF_69/Q_reg  ( .Q(WX719), .CLK(CK), .DIN(WX718) );
  dffs1 \DFF_68/Q_reg  ( .Q(WX717), .CLK(CK), .DIN(WX716) );
  dffs1 \DFF_67/Q_reg  ( .Q(WX715), .CLK(CK), .DIN(WX714) );
  dffs1 \DFF_66/Q_reg  ( .Q(WX713), .CLK(CK), .DIN(WX712) );
  dffs1 \DFF_65/Q_reg  ( .Q(WX711), .CLK(CK), .DIN(WX710) );
  dffs1 \DFF_64/Q_reg  ( .Q(WX709), .CLK(CK), .DIN(WX708) );
  dffs1 \DFF_63/Q_reg  ( .Q(WX707), .CLK(CK), .DIN(WX706) );
  dffs1 \DFF_62/Q_reg  ( .Q(WX705), .CLK(CK), .DIN(WX704) );
  dffs1 \DFF_61/Q_reg  ( .Q(WX703), .CLK(CK), .DIN(WX702) );
  dffs1 \DFF_60/Q_reg  ( .Q(WX701), .CLK(CK), .DIN(WX700) );
  dffs1 \DFF_59/Q_reg  ( .Q(WX699), .CLK(CK), .DIN(WX698) );
  dffs1 \DFF_58/Q_reg  ( .Q(WX697), .CLK(CK), .DIN(WX696) );
  dffs1 \DFF_57/Q_reg  ( .Q(WX695), .CLK(CK), .DIN(WX694) );
  dffs1 \DFF_56/Q_reg  ( .Q(WX693), .CLK(CK), .DIN(WX692) );
  dffs1 \DFF_55/Q_reg  ( .Q(WX691), .CLK(CK), .DIN(WX690) );
  dffs1 \DFF_54/Q_reg  ( .Q(WX689), .CLK(CK), .DIN(WX688) );
  dffs1 \DFF_53/Q_reg  ( .Q(WX687), .CLK(CK), .DIN(WX686) );
  dffs1 \DFF_52/Q_reg  ( .Q(WX685), .CLK(CK), .DIN(WX684) );
  dffs1 \DFF_51/Q_reg  ( .Q(WX683), .CLK(CK), .DIN(WX682) );
  dffs1 \DFF_50/Q_reg  ( .Q(WX681), .CLK(CK), .DIN(WX680) );
  dffs1 \DFF_49/Q_reg  ( .Q(WX679), .CLK(CK), .DIN(WX678) );
  dffs1 \DFF_48/Q_reg  ( .Q(WX677), .CLK(CK), .DIN(WX676) );
  dffs1 \DFF_47/Q_reg  ( .Q(WX675), .CLK(CK), .DIN(WX674) );
  dffs1 \DFF_46/Q_reg  ( .Q(WX673), .CLK(CK), .DIN(WX672) );
  dffs1 \DFF_45/Q_reg  ( .Q(WX671), .CLK(CK), .DIN(WX670) );
  dffs1 \DFF_44/Q_reg  ( .Q(WX669), .CLK(CK), .DIN(WX668) );
  dffs1 \DFF_43/Q_reg  ( .Q(WX667), .CLK(CK), .DIN(WX666) );
  dffs1 \DFF_42/Q_reg  ( .Q(WX665), .CLK(CK), .DIN(WX664) );
  dffs1 \DFF_41/Q_reg  ( .Q(WX663), .CLK(CK), .DIN(WX662) );
  dffs1 \DFF_40/Q_reg  ( .Q(WX661), .CLK(CK), .DIN(WX660) );
  dffs1 \DFF_39/Q_reg  ( .Q(WX659), .CLK(CK), .DIN(WX658) );
  dffs1 \DFF_38/Q_reg  ( .Q(WX657), .CLK(CK), .DIN(WX656) );
  dffs1 \DFF_37/Q_reg  ( .Q(WX655), .CLK(CK), .DIN(WX654) );
  dffs1 \DFF_36/Q_reg  ( .Q(WX653), .CLK(CK), .DIN(WX652) );
  dffs1 \DFF_35/Q_reg  ( .Q(WX651), .CLK(CK), .DIN(WX650) );
  dffs1 \DFF_34/Q_reg  ( .Q(WX649), .CLK(CK), .DIN(WX648) );
  dffs1 \DFF_33/Q_reg  ( .Q(WX647), .CLK(CK), .DIN(WX646) );
  dffs1 \DFF_32/Q_reg  ( .Q(WX645), .CLK(CK), .DIN(WX644) );
  dffs1 \DFF_31/Q_reg  ( .Q(WX547), .CLK(CK), .DIN(WX546) );
  dffs1 \DFF_30/Q_reg  ( .Q(WX545), .CLK(CK), .DIN(WX544) );
  dffs1 \DFF_29/Q_reg  ( .Q(WX543), .CLK(CK), .DIN(WX542) );
  dffs1 \DFF_28/Q_reg  ( .Q(WX541), .CLK(CK), .DIN(WX540) );
  dffs1 \DFF_27/Q_reg  ( .Q(WX539), .CLK(CK), .DIN(WX538) );
  dffs1 \DFF_26/Q_reg  ( .Q(WX537), .CLK(CK), .DIN(WX536) );
  dffs1 \DFF_25/Q_reg  ( .Q(WX535), .CLK(CK), .DIN(WX534) );
  dffs1 \DFF_24/Q_reg  ( .Q(WX533), .CLK(CK), .DIN(WX532) );
  dffs1 \DFF_23/Q_reg  ( .Q(WX531), .CLK(CK), .DIN(WX530) );
  dffs1 \DFF_22/Q_reg  ( .Q(WX529), .CLK(CK), .DIN(WX528) );
  dffs1 \DFF_21/Q_reg  ( .Q(WX527), .CLK(CK), .DIN(WX526) );
  dffs1 \DFF_20/Q_reg  ( .Q(WX525), .CLK(CK), .DIN(WX524) );
  dffs1 \DFF_19/Q_reg  ( .Q(WX523), .CLK(CK), .DIN(WX522) );
  dffs1 \DFF_18/Q_reg  ( .Q(WX521), .CLK(CK), .DIN(WX520) );
  dffs1 \DFF_17/Q_reg  ( .Q(WX519), .CLK(CK), .DIN(WX518) );
  dffs1 \DFF_16/Q_reg  ( .Q(WX517), .CLK(CK), .DIN(WX516) );
  dffs1 \DFF_15/Q_reg  ( .Q(WX515), .CLK(CK), .DIN(WX514) );
  dffs1 \DFF_14/Q_reg  ( .Q(WX513), .CLK(CK), .DIN(WX512) );
  dffs1 \DFF_13/Q_reg  ( .Q(WX511), .CLK(CK), .DIN(WX510) );
  dffs1 \DFF_12/Q_reg  ( .Q(WX509), .CLK(CK), .DIN(WX508) );
  dffs1 \DFF_11/Q_reg  ( .Q(WX507), .CLK(CK), .DIN(WX506) );
  dffs1 \DFF_10/Q_reg  ( .Q(WX505), .CLK(CK), .DIN(WX504) );
  dffs1 \DFF_9/Q_reg  ( .Q(WX503), .CLK(CK), .DIN(WX502) );
  dffs1 \DFF_8/Q_reg  ( .Q(WX501), .CLK(CK), .DIN(WX500) );
  dffs1 \DFF_7/Q_reg  ( .Q(WX499), .CLK(CK), .DIN(WX498) );
  dffs1 \DFF_6/Q_reg  ( .Q(WX497), .CLK(CK), .DIN(WX496) );
  dffs1 \DFF_5/Q_reg  ( .Q(WX495), .CLK(CK), .DIN(WX494) );
  dffs1 \DFF_4/Q_reg  ( .Q(WX493), .CLK(CK), .DIN(WX492) );
  dffs1 \DFF_3/Q_reg  ( .Q(WX491), .CLK(CK), .DIN(WX490) );
  dffs1 \DFF_2/Q_reg  ( .Q(WX489), .CLK(CK), .DIN(WX488) );
  dffs1 \DFF_1/Q_reg  ( .Q(WX487), .CLK(CK), .DIN(WX486) );
  dffs1 \DFF_0/Q_reg  ( .Q(WX485), .CLK(CK), .DIN(WX484) );
endmodule

