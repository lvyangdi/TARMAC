module c1355 (N1, N8, N15, N22, N29, N36, N43, N50, N57, N64, N71, N78, N85, N92, N99, N106, N113, N120, N127, N134, N141, N148, N155, N162, N169, N176, N183, N190, N197, N204, N211, N218, N225, N226, N227, N228, N229, N230, N231, N232, N233, N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354, N1355);

input N1, N8, N15, N22, N29, N36, N43, N50, N57, N64, N71, N78, N85, N92, N99, N106, N113, N120, N127, N134, N141, N148, N155, N162, N169, N176, N183, N190, N197, N204, N211, N218, N225, N226, N227, N228, N229, N230, N231, N232, N233;

output N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353, N1354, N1355;

wire N242, N245, N248, N251, N254, N257, N260, N263, N266, N269, N272, N275, N278, N281, N284, N287, N290, N293, N296, N299, N302, N305, N308, N311, N314, N317, N320, N323, N326, N329, N332, N335, N338, N341, N344, N347, N350, N353, N356, N359, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N429, N432, N435, N438, N441, N444, N447, N450, N453, N456, N459, N462, N465, N468, N471, N474, N477, N480, N483, N486, N489, N492, N495, N498, N501, N504, N507, N510, N513, N516, N519, N522, N525, N528, N531, N534, N537, N540, N543, N546, N549, N552, N555, N558, N561, N564, N567, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601, N602, N607, N612, N617, N622, N627, N632, N637, N642, N645, N648, N651, N654, N657, N660, N663, N666, N669, N672, N675, N678, N681, N684, N687, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703, N704, N705, N706, N709, N712, N715, N718, N721, N724, N727, N730, N733, N736, N739, N742, N745, N748, N751, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N773, N776, N779, N782, N785, N788, N791, N794, N797, N800, N803, N806, N809, N812, N815, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N847, N860, N873, N886, N899, N912, N925, N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985, N986, N991, N996, N1001, N1006, N1011, N1016, N1021, N1026, N1031, N1036, N1039, N1042, N1045, N1048, N1051, N1054, N1057, N1060, N1063, N1066, N1069, N1072, N1075, N1078, N1081, N1084, N1087, N1090, N1093, N1096, N1099, N1102, N1105, N1108, N1111, N1114, N1117, N1120, N1123, N1126, N1129, N1132, N1135, N1138, N1141, N1144, N1147, N1150, N1153, N1156, N1159, N1162, N1165, N1168, N1171, N1174, N1177, N1180, N1183, N1186, N1189, N1192, N1195, N1198, N1201, N1204, N1207, N1210, N1213, N1216, N1219, N1222, N1225, N1228, N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242, N1243, N1244, N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262, N1263, N1264, N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272, N1273, N1274, N1275, N1276, N1277, N1278, N1279, N1280, N1281, N1282, N1283, N1284, N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292, N1293, N1294, N1295, N1296, N1297, N1298, N1299, N1300, N1301, N1302, N1303, N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313, N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323;

and2s1 U1 (.Q(N242), .DIN1(N225), .DIN2(N233));
and2s1 U2 (.Q(N245), .DIN1(N226), .DIN2(N233));
and2s1 U3 (.Q(N248), .DIN1(N227), .DIN2(N233));
and2s1 U4 (.Q(N251), .DIN1(N228), .DIN2(N233));
and2s1 U5 (.Q(N254), .DIN1(N229), .DIN2(N233));
and2s1 U6 (.Q(N257), .DIN1(N230), .DIN2(N233));
and2s1 U7 (.Q(N260), .DIN1(N231), .DIN2(N233));
and2s1 U8 (.Q(N263), .DIN1(N232), .DIN2(N233));
nnd2s1 U9 (.Q(N266), .DIN1(N1), .DIN2(N8));
nnd2s1 U10 (.Q(N269), .DIN1(N15), .DIN2(N22));
nnd2s1 U11 (.Q(N272), .DIN1(N29), .DIN2(N36));
nnd2s1 U12 (.Q(N275), .DIN1(N43), .DIN2(N50));
nnd2s1 U13 (.Q(N278), .DIN1(N57), .DIN2(N64));
nnd2s1 U14 (.Q(N281), .DIN1(N71), .DIN2(N78));
nnd2s1 U15 (.Q(N284), .DIN1(N85), .DIN2(N92));
nnd2s1 U16 (.Q(N287), .DIN1(N99), .DIN2(N106));
nnd2s1 U17 (.Q(N290), .DIN1(N113), .DIN2(N120));
nnd2s1 U18 (.Q(N293), .DIN1(N127), .DIN2(N134));
nnd2s1 U19 (.Q(N296), .DIN1(N141), .DIN2(N148));
nnd2s1 U20 (.Q(N299), .DIN1(N155), .DIN2(N162));
nnd2s1 U21 (.Q(N302), .DIN1(N169), .DIN2(N176));
nnd2s1 U22 (.Q(N305), .DIN1(N183), .DIN2(N190));
nnd2s1 U23 (.Q(N308), .DIN1(N197), .DIN2(N204));
nnd2s1 U24 (.Q(N311), .DIN1(N211), .DIN2(N218));
nnd2s1 U25 (.Q(N314), .DIN1(N1), .DIN2(N29));
nnd2s1 U26 (.Q(N317), .DIN1(N57), .DIN2(N85));
nnd2s1 U27 (.Q(N320), .DIN1(N8), .DIN2(N36));
nnd2s1 U28 (.Q(N323), .DIN1(N64), .DIN2(N92));
nnd2s1 U29 (.Q(N326), .DIN1(N15), .DIN2(N43));
nnd2s1 U30 (.Q(N329), .DIN1(N71), .DIN2(N99));
nnd2s1 U31 (.Q(N332), .DIN1(N22), .DIN2(N50));
nnd2s1 U32 (.Q(N335), .DIN1(N78), .DIN2(N106));
nnd2s1 U33 (.Q(N338), .DIN1(N113), .DIN2(N141));
nnd2s1 U34 (.Q(N341), .DIN1(N169), .DIN2(N197));
nnd2s1 U35 (.Q(N344), .DIN1(N120), .DIN2(N148));
nnd2s1 U36 (.Q(N347), .DIN1(N176), .DIN2(N204));
nnd2s1 U37 (.Q(N350), .DIN1(N127), .DIN2(N155));
nnd2s1 U38 (.Q(N353), .DIN1(N183), .DIN2(N211));
nnd2s1 U39 (.Q(N356), .DIN1(N134), .DIN2(N162));
nnd2s1 U40 (.Q(N359), .DIN1(N190), .DIN2(N218));
nnd2s1 U41 (.Q(N362), .DIN1(N1), .DIN2(N266));
nnd2s1 U42 (.Q(N363), .DIN1(N8), .DIN2(N266));
nnd2s1 U43 (.Q(N364), .DIN1(N15), .DIN2(N269));
nnd2s1 U44 (.Q(N365), .DIN1(N22), .DIN2(N269));
nnd2s1 U45 (.Q(N366), .DIN1(N29), .DIN2(N272));
nnd2s1 U46 (.Q(N367), .DIN1(N36), .DIN2(N272));
nnd2s1 U47 (.Q(N368), .DIN1(N43), .DIN2(N275));
nnd2s1 U48 (.Q(N369), .DIN1(N50), .DIN2(N275));
nnd2s1 U49 (.Q(N370), .DIN1(N57), .DIN2(N278));
nnd2s1 U50 (.Q(N371), .DIN1(N64), .DIN2(N278));
nnd2s1 U51 (.Q(N372), .DIN1(N71), .DIN2(N281));
nnd2s1 U52 (.Q(N373), .DIN1(N78), .DIN2(N281));
nnd2s1 U53 (.Q(N374), .DIN1(N85), .DIN2(N284));
nnd2s1 U54 (.Q(N375), .DIN1(N92), .DIN2(N284));
nnd2s1 U55 (.Q(N376), .DIN1(N99), .DIN2(N287));
nnd2s1 U56 (.Q(N377), .DIN1(N106), .DIN2(N287));
nnd2s1 U57 (.Q(N378), .DIN1(N113), .DIN2(N290));
nnd2s1 U58 (.Q(N379), .DIN1(N120), .DIN2(N290));
nnd2s1 U59 (.Q(N380), .DIN1(N127), .DIN2(N293));
nnd2s1 U60 (.Q(N381), .DIN1(N134), .DIN2(N293));
nnd2s1 U61 (.Q(N382), .DIN1(N141), .DIN2(N296));
nnd2s1 U62 (.Q(N383), .DIN1(N148), .DIN2(N296));
nnd2s1 U63 (.Q(N384), .DIN1(N155), .DIN2(N299));
nnd2s1 U64 (.Q(N385), .DIN1(N162), .DIN2(N299));
nnd2s1 U65 (.Q(N386), .DIN1(N169), .DIN2(N302));
nnd2s1 U66 (.Q(N387), .DIN1(N176), .DIN2(N302));
nnd2s1 U67 (.Q(N388), .DIN1(N183), .DIN2(N305));
nnd2s1 U68 (.Q(N389), .DIN1(N190), .DIN2(N305));
nnd2s1 U69 (.Q(N390), .DIN1(N197), .DIN2(N308));
nnd2s1 U70 (.Q(N391), .DIN1(N204), .DIN2(N308));
nnd2s1 U71 (.Q(N392), .DIN1(N211), .DIN2(N311));
nnd2s1 U72 (.Q(N393), .DIN1(N218), .DIN2(N311));
nnd2s1 U73 (.Q(N394), .DIN1(N1), .DIN2(N314));
nnd2s1 U74 (.Q(N395), .DIN1(N29), .DIN2(N314));
nnd2s1 U75 (.Q(N396), .DIN1(N57), .DIN2(N317));
nnd2s1 U76 (.Q(N397), .DIN1(N85), .DIN2(N317));
nnd2s1 U77 (.Q(N398), .DIN1(N8), .DIN2(N320));
nnd2s1 U78 (.Q(N399), .DIN1(N36), .DIN2(N320));
nnd2s1 U79 (.Q(N400), .DIN1(N64), .DIN2(N323));
nnd2s1 U80 (.Q(N401), .DIN1(N92), .DIN2(N323));
nnd2s1 U81 (.Q(N402), .DIN1(N15), .DIN2(N326));
nnd2s1 U82 (.Q(N403), .DIN1(N43), .DIN2(N326));
nnd2s1 U83 (.Q(N404), .DIN1(N71), .DIN2(N329));
nnd2s1 U84 (.Q(N405), .DIN1(N99), .DIN2(N329));
nnd2s1 U85 (.Q(N406), .DIN1(N22), .DIN2(N332));
nnd2s1 U86 (.Q(N407), .DIN1(N50), .DIN2(N332));
nnd2s1 U87 (.Q(N408), .DIN1(N78), .DIN2(N335));
nnd2s1 U88 (.Q(N409), .DIN1(N106), .DIN2(N335));
nnd2s1 U89 (.Q(N410), .DIN1(N113), .DIN2(N338));
nnd2s1 U90 (.Q(N411), .DIN1(N141), .DIN2(N338));
nnd2s1 U91 (.Q(N412), .DIN1(N169), .DIN2(N341));
nnd2s1 U92 (.Q(N413), .DIN1(N197), .DIN2(N341));
nnd2s1 U93 (.Q(N414), .DIN1(N120), .DIN2(N344));
nnd2s1 U94 (.Q(N415), .DIN1(N148), .DIN2(N344));
nnd2s1 U95 (.Q(N416), .DIN1(N176), .DIN2(N347));
nnd2s1 U96 (.Q(N417), .DIN1(N204), .DIN2(N347));
nnd2s1 U97 (.Q(N418), .DIN1(N127), .DIN2(N350));
nnd2s1 U98 (.Q(N419), .DIN1(N155), .DIN2(N350));
nnd2s1 U99 (.Q(N420), .DIN1(N183), .DIN2(N353));
nnd2s1 U100 (.Q(N421), .DIN1(N211), .DIN2(N353));
nnd2s1 U101 (.Q(N422), .DIN1(N134), .DIN2(N356));
nnd2s1 U102 (.Q(N423), .DIN1(N162), .DIN2(N356));
nnd2s1 U103 (.Q(N424), .DIN1(N190), .DIN2(N359));
nnd2s1 U104 (.Q(N425), .DIN1(N218), .DIN2(N359));
nnd2s1 U105 (.Q(N426), .DIN1(N362), .DIN2(N363));
nnd2s1 U106 (.Q(N429), .DIN1(N364), .DIN2(N365));
nnd2s1 U107 (.Q(N432), .DIN1(N366), .DIN2(N367));
nnd2s1 U108 (.Q(N435), .DIN1(N368), .DIN2(N369));
nnd2s1 U109 (.Q(N438), .DIN1(N370), .DIN2(N371));
nnd2s1 U110 (.Q(N441), .DIN1(N372), .DIN2(N373));
nnd2s1 U111 (.Q(N444), .DIN1(N374), .DIN2(N375));
nnd2s1 U112 (.Q(N447), .DIN1(N376), .DIN2(N377));
nnd2s1 U113 (.Q(N450), .DIN1(N378), .DIN2(N379));
nnd2s1 U114 (.Q(N453), .DIN1(N380), .DIN2(N381));
nnd2s1 U115 (.Q(N456), .DIN1(N382), .DIN2(N383));
nnd2s1 U116 (.Q(N459), .DIN1(N384), .DIN2(N385));
nnd2s1 U117 (.Q(N462), .DIN1(N386), .DIN2(N387));
nnd2s1 U118 (.Q(N465), .DIN1(N388), .DIN2(N389));
nnd2s1 U119 (.Q(N468), .DIN1(N390), .DIN2(N391));
nnd2s1 U120 (.Q(N471), .DIN1(N392), .DIN2(N393));
nnd2s1 U121 (.Q(N474), .DIN1(N394), .DIN2(N395));
nnd2s1 U122 (.Q(N477), .DIN1(N396), .DIN2(N397));
nnd2s1 U123 (.Q(N480), .DIN1(N398), .DIN2(N399));
nnd2s1 U124 (.Q(N483), .DIN1(N400), .DIN2(N401));
nnd2s1 U125 (.Q(N486), .DIN1(N402), .DIN2(N403));
nnd2s1 U126 (.Q(N489), .DIN1(N404), .DIN2(N405));
nnd2s1 U127 (.Q(N492), .DIN1(N406), .DIN2(N407));
nnd2s1 U128 (.Q(N495), .DIN1(N408), .DIN2(N409));
nnd2s1 U129 (.Q(N498), .DIN1(N410), .DIN2(N411));
nnd2s1 U130 (.Q(N501), .DIN1(N412), .DIN2(N413));
nnd2s1 U131 (.Q(N504), .DIN1(N414), .DIN2(N415));
nnd2s1 U132 (.Q(N507), .DIN1(N416), .DIN2(N417));
nnd2s1 U133 (.Q(N510), .DIN1(N418), .DIN2(N419));
nnd2s1 U134 (.Q(N513), .DIN1(N420), .DIN2(N421));
nnd2s1 U135 (.Q(N516), .DIN1(N422), .DIN2(N423));
nnd2s1 U136 (.Q(N519), .DIN1(N424), .DIN2(N425));
nnd2s1 U137 (.Q(N522), .DIN1(N426), .DIN2(N429));
nnd2s1 U138 (.Q(N525), .DIN1(N432), .DIN2(N435));
nnd2s1 U139 (.Q(N528), .DIN1(N438), .DIN2(N441));
nnd2s1 U140 (.Q(N531), .DIN1(N444), .DIN2(N447));
nnd2s1 U141 (.Q(N534), .DIN1(N450), .DIN2(N453));
nnd2s1 U142 (.Q(N537), .DIN1(N456), .DIN2(N459));
nnd2s1 U143 (.Q(N540), .DIN1(N462), .DIN2(N465));
nnd2s1 U144 (.Q(N543), .DIN1(N468), .DIN2(N471));
nnd2s1 U145 (.Q(N546), .DIN1(N474), .DIN2(N477));
nnd2s1 U146 (.Q(N549), .DIN1(N480), .DIN2(N483));
nnd2s1 U147 (.Q(N552), .DIN1(N486), .DIN2(N489));
nnd2s1 U148 (.Q(N555), .DIN1(N492), .DIN2(N495));
nnd2s1 U149 (.Q(N558), .DIN1(N498), .DIN2(N501));
nnd2s1 U150 (.Q(N561), .DIN1(N504), .DIN2(N507));
nnd2s1 U151 (.Q(N564), .DIN1(N510), .DIN2(N513));
nnd2s1 U152 (.Q(N567), .DIN1(N516), .DIN2(N519));
nnd2s1 U153 (.Q(N570), .DIN1(N426), .DIN2(N522));
nnd2s1 U154 (.Q(N571), .DIN1(N429), .DIN2(N522));
nnd2s1 U155 (.Q(N572), .DIN1(N432), .DIN2(N525));
nnd2s1 U156 (.Q(N573), .DIN1(N435), .DIN2(N525));
nnd2s1 U157 (.Q(N574), .DIN1(N438), .DIN2(N528));
nnd2s1 U158 (.Q(N575), .DIN1(N441), .DIN2(N528));
nnd2s1 U159 (.Q(N576), .DIN1(N444), .DIN2(N531));
nnd2s1 U160 (.Q(N577), .DIN1(N447), .DIN2(N531));
nnd2s1 U161 (.Q(N578), .DIN1(N450), .DIN2(N534));
nnd2s1 U162 (.Q(N579), .DIN1(N453), .DIN2(N534));
nnd2s1 U163 (.Q(N580), .DIN1(N456), .DIN2(N537));
nnd2s1 U164 (.Q(N581), .DIN1(N459), .DIN2(N537));
nnd2s1 U165 (.Q(N582), .DIN1(N462), .DIN2(N540));
nnd2s1 U166 (.Q(N583), .DIN1(N465), .DIN2(N540));
nnd2s1 U167 (.Q(N584), .DIN1(N468), .DIN2(N543));
nnd2s1 U168 (.Q(N585), .DIN1(N471), .DIN2(N543));
nnd2s1 U169 (.Q(N586), .DIN1(N474), .DIN2(N546));
nnd2s1 U170 (.Q(N587), .DIN1(N477), .DIN2(N546));
nnd2s1 U171 (.Q(N588), .DIN1(N480), .DIN2(N549));
nnd2s1 U172 (.Q(N589), .DIN1(N483), .DIN2(N549));
nnd2s1 U173 (.Q(N590), .DIN1(N486), .DIN2(N552));
nnd2s1 U174 (.Q(N591), .DIN1(N489), .DIN2(N552));
nnd2s1 U175 (.Q(N592), .DIN1(N492), .DIN2(N555));
nnd2s1 U176 (.Q(N593), .DIN1(N495), .DIN2(N555));
nnd2s1 U177 (.Q(N594), .DIN1(N498), .DIN2(N558));
nnd2s1 U178 (.Q(N595), .DIN1(N501), .DIN2(N558));
nnd2s1 U179 (.Q(N596), .DIN1(N504), .DIN2(N561));
nnd2s1 U180 (.Q(N597), .DIN1(N507), .DIN2(N561));
nnd2s1 U181 (.Q(N598), .DIN1(N510), .DIN2(N564));
nnd2s1 U182 (.Q(N599), .DIN1(N513), .DIN2(N564));
nnd2s1 U183 (.Q(N600), .DIN1(N516), .DIN2(N567));
nnd2s1 U184 (.Q(N601), .DIN1(N519), .DIN2(N567));
nnd2s1 U185 (.Q(N602), .DIN1(N570), .DIN2(N571));
nnd2s1 U186 (.Q(N607), .DIN1(N572), .DIN2(N573));
nnd2s1 U187 (.Q(N612), .DIN1(N574), .DIN2(N575));
nnd2s1 U188 (.Q(N617), .DIN1(N576), .DIN2(N577));
nnd2s1 U189 (.Q(N622), .DIN1(N578), .DIN2(N579));
nnd2s1 U190 (.Q(N627), .DIN1(N580), .DIN2(N581));
nnd2s1 U191 (.Q(N632), .DIN1(N582), .DIN2(N583));
nnd2s1 U192 (.Q(N637), .DIN1(N584), .DIN2(N585));
nnd2s1 U193 (.Q(N642), .DIN1(N586), .DIN2(N587));
nnd2s1 U194 (.Q(N645), .DIN1(N588), .DIN2(N589));
nnd2s1 U195 (.Q(N648), .DIN1(N590), .DIN2(N591));
nnd2s1 U196 (.Q(N651), .DIN1(N592), .DIN2(N593));
nnd2s1 U197 (.Q(N654), .DIN1(N594), .DIN2(N595));
nnd2s1 U198 (.Q(N657), .DIN1(N596), .DIN2(N597));
nnd2s1 U199 (.Q(N660), .DIN1(N598), .DIN2(N599));
nnd2s1 U200 (.Q(N663), .DIN1(N600), .DIN2(N601));
nnd2s1 U201 (.Q(N666), .DIN1(N602), .DIN2(N607));
nnd2s1 U202 (.Q(N669), .DIN1(N612), .DIN2(N617));
nnd2s1 U203 (.Q(N672), .DIN1(N602), .DIN2(N612));
nnd2s1 U204 (.Q(N675), .DIN1(N607), .DIN2(N617));
nnd2s1 U205 (.Q(N678), .DIN1(N622), .DIN2(N627));
nnd2s1 U206 (.Q(N681), .DIN1(N632), .DIN2(N637));
nnd2s1 U207 (.Q(N684), .DIN1(N622), .DIN2(N632));
nnd2s1 U208 (.Q(N687), .DIN1(N627), .DIN2(N637));
nnd2s1 U209 (.Q(N690), .DIN1(N602), .DIN2(N666));
nnd2s1 U210 (.Q(N691), .DIN1(N607), .DIN2(N666));
nnd2s1 U211 (.Q(N692), .DIN1(N612), .DIN2(N669));
nnd2s1 U212 (.Q(N693), .DIN1(N617), .DIN2(N669));
nnd2s1 U213 (.Q(N694), .DIN1(N602), .DIN2(N672));
nnd2s1 U214 (.Q(N695), .DIN1(N612), .DIN2(N672));
nnd2s1 U215 (.Q(N696), .DIN1(N607), .DIN2(N675));
nnd2s1 U216 (.Q(N697), .DIN1(N617), .DIN2(N675));
nnd2s1 U217 (.Q(N698), .DIN1(N622), .DIN2(N678));
nnd2s1 U218 (.Q(N699), .DIN1(N627), .DIN2(N678));
nnd2s1 U219 (.Q(N700), .DIN1(N632), .DIN2(N681));
nnd2s1 U220 (.Q(N701), .DIN1(N637), .DIN2(N681));
nnd2s1 U221 (.Q(N702), .DIN1(N622), .DIN2(N684));
nnd2s1 U222 (.Q(N703), .DIN1(N632), .DIN2(N684));
nnd2s1 U223 (.Q(N704), .DIN1(N627), .DIN2(N687));
nnd2s1 U224 (.Q(N705), .DIN1(N637), .DIN2(N687));
nnd2s1 U225 (.Q(N706), .DIN1(N690), .DIN2(N691));
nnd2s1 U226 (.Q(N709), .DIN1(N692), .DIN2(N693));
nnd2s1 U227 (.Q(N712), .DIN1(N694), .DIN2(N695));
nnd2s1 U228 (.Q(N715), .DIN1(N696), .DIN2(N697));
nnd2s1 U229 (.Q(N718), .DIN1(N698), .DIN2(N699));
nnd2s1 U230 (.Q(N721), .DIN1(N700), .DIN2(N701));
nnd2s1 U231 (.Q(N724), .DIN1(N702), .DIN2(N703));
nnd2s1 U232 (.Q(N727), .DIN1(N704), .DIN2(N705));
nnd2s1 U233 (.Q(N730), .DIN1(N242), .DIN2(N718));
nnd2s1 U234 (.Q(N733), .DIN1(N245), .DIN2(N721));
nnd2s1 U235 (.Q(N736), .DIN1(N248), .DIN2(N724));
nnd2s1 U236 (.Q(N739), .DIN1(N251), .DIN2(N727));
nnd2s1 U237 (.Q(N742), .DIN1(N254), .DIN2(N706));
nnd2s1 U238 (.Q(N745), .DIN1(N257), .DIN2(N709));
nnd2s1 U239 (.Q(N748), .DIN1(N260), .DIN2(N712));
nnd2s1 U240 (.Q(N751), .DIN1(N263), .DIN2(N715));
nnd2s1 U241 (.Q(N754), .DIN1(N242), .DIN2(N730));
nnd2s1 U242 (.Q(N755), .DIN1(N718), .DIN2(N730));
nnd2s1 U243 (.Q(N756), .DIN1(N245), .DIN2(N733));
nnd2s1 U244 (.Q(N757), .DIN1(N721), .DIN2(N733));
nnd2s1 U245 (.Q(N758), .DIN1(N248), .DIN2(N736));
nnd2s1 U246 (.Q(N759), .DIN1(N724), .DIN2(N736));
nnd2s1 U247 (.Q(N760), .DIN1(N251), .DIN2(N739));
nnd2s1 U248 (.Q(N761), .DIN1(N727), .DIN2(N739));
nnd2s1 U249 (.Q(N762), .DIN1(N254), .DIN2(N742));
nnd2s1 U250 (.Q(N763), .DIN1(N706), .DIN2(N742));
nnd2s1 U251 (.Q(N764), .DIN1(N257), .DIN2(N745));
nnd2s1 U252 (.Q(N765), .DIN1(N709), .DIN2(N745));
nnd2s1 U253 (.Q(N766), .DIN1(N260), .DIN2(N748));
nnd2s1 U254 (.Q(N767), .DIN1(N712), .DIN2(N748));
nnd2s1 U255 (.Q(N768), .DIN1(N263), .DIN2(N751));
nnd2s1 U256 (.Q(N769), .DIN1(N715), .DIN2(N751));
nnd2s1 U257 (.Q(N770), .DIN1(N754), .DIN2(N755));
nnd2s1 U258 (.Q(N773), .DIN1(N756), .DIN2(N757));
nnd2s1 U259 (.Q(N776), .DIN1(N758), .DIN2(N759));
nnd2s1 U260 (.Q(N779), .DIN1(N760), .DIN2(N761));
nnd2s1 U261 (.Q(N782), .DIN1(N762), .DIN2(N763));
nnd2s1 U262 (.Q(N785), .DIN1(N764), .DIN2(N765));
nnd2s1 U263 (.Q(N788), .DIN1(N766), .DIN2(N767));
nnd2s1 U264 (.Q(N791), .DIN1(N768), .DIN2(N769));
nnd2s1 U265 (.Q(N794), .DIN1(N642), .DIN2(N770));
nnd2s1 U266 (.Q(N797), .DIN1(N645), .DIN2(N773));
nnd2s1 U267 (.Q(N800), .DIN1(N648), .DIN2(N776));
nnd2s1 U268 (.Q(N803), .DIN1(N651), .DIN2(N779));
nnd2s1 U269 (.Q(N806), .DIN1(N654), .DIN2(N782));
nnd2s1 U270 (.Q(N809), .DIN1(N657), .DIN2(N785));
nnd2s1 U271 (.Q(N812), .DIN1(N660), .DIN2(N788));
nnd2s1 U272 (.Q(N815), .DIN1(N663), .DIN2(N791));
nnd2s1 U273 (.Q(N818), .DIN1(N642), .DIN2(N794));
nnd2s1 U274 (.Q(N819), .DIN1(N770), .DIN2(N794));
nnd2s1 U275 (.Q(N820), .DIN1(N645), .DIN2(N797));
nnd2s1 U276 (.Q(N821), .DIN1(N773), .DIN2(N797));
nnd2s1 U277 (.Q(N822), .DIN1(N648), .DIN2(N800));
nnd2s1 U278 (.Q(N823), .DIN1(N776), .DIN2(N800));
nnd2s1 U279 (.Q(N824), .DIN1(N651), .DIN2(N803));
nnd2s1 U280 (.Q(N825), .DIN1(N779), .DIN2(N803));
nnd2s1 U281 (.Q(N826), .DIN1(N654), .DIN2(N806));
nnd2s1 U282 (.Q(N827), .DIN1(N782), .DIN2(N806));
nnd2s1 U283 (.Q(N828), .DIN1(N657), .DIN2(N809));
nnd2s1 U284 (.Q(N829), .DIN1(N785), .DIN2(N809));
nnd2s1 U285 (.Q(N830), .DIN1(N660), .DIN2(N812));
nnd2s1 U286 (.Q(N831), .DIN1(N788), .DIN2(N812));
nnd2s1 U287 (.Q(N832), .DIN1(N663), .DIN2(N815));
nnd2s1 U288 (.Q(N833), .DIN1(N791), .DIN2(N815));
nnd2s1 U289 (.Q(N834), .DIN1(N818), .DIN2(N819));
nnd2s1 U290 (.Q(N847), .DIN1(N820), .DIN2(N821));
nnd2s1 U291 (.Q(N860), .DIN1(N822), .DIN2(N823));
nnd2s1 U292 (.Q(N873), .DIN1(N824), .DIN2(N825));
nnd2s1 U293 (.Q(N886), .DIN1(N828), .DIN2(N829));
nnd2s1 U294 (.Q(N899), .DIN1(N832), .DIN2(N833));
nnd2s1 U295 (.Q(N912), .DIN1(N830), .DIN2(N831));
nnd2s1 U296 (.Q(N925), .DIN1(N826), .DIN2(N827));
hi1s1 U297 (.Q(N938), .DIN(N834));
hi1s1 U298 (.Q(N939), .DIN(N847));
hi1s1 U299 (.Q(N940), .DIN(N860));
hi1s1 U300 (.Q(N941), .DIN(N834));
hi1s1 U301 (.Q(N942), .DIN(N847));
hi1s1 U302 (.Q(N943), .DIN(N873));
hi1s1 U303 (.Q(N944), .DIN(N834));
hi1s1 U304 (.Q(N945), .DIN(N860));
hi1s1 U305 (.Q(N946), .DIN(N873));
hi1s1 U306 (.Q(N947), .DIN(N847));
hi1s1 U307 (.Q(N948), .DIN(N860));
hi1s1 U308 (.Q(N949), .DIN(N873));
hi1s1 U309 (.Q(N950), .DIN(N886));
hi1s1 U310 (.Q(N951), .DIN(N899));
hi1s1 U311 (.Q(N952), .DIN(N886));
hi1s1 U312 (.Q(N953), .DIN(N912));
hi1s1 U313 (.Q(N954), .DIN(N925));
hi1s1 U314 (.Q(N955), .DIN(N899));
hi1s1 U315 (.Q(N956), .DIN(N925));
hi1s1 U316 (.Q(N957), .DIN(N912));
hi1s1 U317 (.Q(N958), .DIN(N925));
hi1s1 U318 (.Q(N959), .DIN(N886));
hi1s1 U319 (.Q(N960), .DIN(N912));
hi1s1 U320 (.Q(N961), .DIN(N925));
hi1s1 U321 (.Q(N962), .DIN(N886));
hi1s1 U322 (.Q(N963), .DIN(N899));
hi1s1 U323 (.Q(N964), .DIN(N925));
hi1s1 U324 (.Q(N965), .DIN(N912));
hi1s1 U325 (.Q(N966), .DIN(N899));
hi1s1 U326 (.Q(N967), .DIN(N886));
hi1s1 U327 (.Q(N968), .DIN(N912));
hi1s1 U328 (.Q(N969), .DIN(N899));
hi1s1 U329 (.Q(N970), .DIN(N847));
hi1s1 U330 (.Q(N971), .DIN(N873));
hi1s1 U331 (.Q(N972), .DIN(N847));
hi1s1 U332 (.Q(N973), .DIN(N860));
hi1s1 U333 (.Q(N974), .DIN(N834));
hi1s1 U334 (.Q(N975), .DIN(N873));
hi1s1 U335 (.Q(N976), .DIN(N834));
hi1s1 U336 (.Q(N977), .DIN(N860));
and4s1 U337 (.Q(N978), .DIN1(N938), .DIN2(N939), .DIN3(N940), .DIN4(N873));
and4s1 U338 (.Q(N979), .DIN1(N941), .DIN2(N942), .DIN3(N860), .DIN4(N943));
and4s1 U339 (.Q(N980), .DIN1(N944), .DIN2(N847), .DIN3(N945), .DIN4(N946));
and4s1 U340 (.Q(N981), .DIN1(N834), .DIN2(N947), .DIN3(N948), .DIN4(N949));
and4s1 U341 (.Q(N982), .DIN1(N958), .DIN2(N959), .DIN3(N960), .DIN4(N899));
and4s1 U342 (.Q(N983), .DIN1(N961), .DIN2(N962), .DIN3(N912), .DIN4(N963));
and4s1 U343 (.Q(N984), .DIN1(N964), .DIN2(N886), .DIN3(N965), .DIN4(N966));
and4s1 U344 (.Q(N985), .DIN1(N925), .DIN2(N967), .DIN3(N968), .DIN4(N969));
or4s1 U345 (.Q(N986), .DIN1(N978), .DIN2(N979), .DIN3(N980), .DIN4(N981));
or4s1 U346 (.Q(N991), .DIN1(N982), .DIN2(N983), .DIN3(N984), .DIN4(N985));
and5s1 U347 (.Q(N996), .DIN1(N925), .DIN2(N950), .DIN3(N912), .DIN4(N951), .DIN5(N986));
and5s1 U348 (.Q(N1001), .DIN1(N925), .DIN2(N952), .DIN3(N953), .DIN4(N899), .DIN5(N986));
and5s1 U349 (.Q(N1006), .DIN1(N954), .DIN2(N886), .DIN3(N912), .DIN4(N955), .DIN5(N986));
and5s1 U350 (.Q(N1011), .DIN1(N956), .DIN2(N886), .DIN3(N957), .DIN4(N899), .DIN5(N986));
and5s1 U351 (.Q(N1016), .DIN1(N834), .DIN2(N970), .DIN3(N860), .DIN4(N971), .DIN5(N991));
and5s1 U352 (.Q(N1021), .DIN1(N834), .DIN2(N972), .DIN3(N973), .DIN4(N873), .DIN5(N991));
and5s1 U353 (.Q(N1026), .DIN1(N974), .DIN2(N847), .DIN3(N860), .DIN4(N975), .DIN5(N991));
and5s1 U354 (.Q(N1031), .DIN1(N976), .DIN2(N847), .DIN3(N977), .DIN4(N873), .DIN5(N991));
and2s1 U355 (.Q(N1036), .DIN1(N834), .DIN2(N996));
and2s1 U356 (.Q(N1039), .DIN1(N847), .DIN2(N996));
and2s1 U357 (.Q(N1042), .DIN1(N860), .DIN2(N996));
and2s1 U358 (.Q(N1045), .DIN1(N873), .DIN2(N996));
and2s1 U359 (.Q(N1048), .DIN1(N834), .DIN2(N1001));
and2s1 U360 (.Q(N1051), .DIN1(N847), .DIN2(N1001));
and2s1 U361 (.Q(N1054), .DIN1(N860), .DIN2(N1001));
and2s1 U362 (.Q(N1057), .DIN1(N873), .DIN2(N1001));
and2s1 U363 (.Q(N1060), .DIN1(N834), .DIN2(N1006));
and2s1 U364 (.Q(N1063), .DIN1(N847), .DIN2(N1006));
and2s1 U365 (.Q(N1066), .DIN1(N860), .DIN2(N1006));
and2s1 U366 (.Q(N1069), .DIN1(N873), .DIN2(N1006));
and2s1 U367 (.Q(N1072), .DIN1(N834), .DIN2(N1011));
and2s1 U368 (.Q(N1075), .DIN1(N847), .DIN2(N1011));
and2s1 U369 (.Q(N1078), .DIN1(N860), .DIN2(N1011));
and2s1 U370 (.Q(N1081), .DIN1(N873), .DIN2(N1011));
and2s1 U371 (.Q(N1084), .DIN1(N925), .DIN2(N1016));
and2s1 U372 (.Q(N1087), .DIN1(N886), .DIN2(N1016));
and2s1 U373 (.Q(N1090), .DIN1(N912), .DIN2(N1016));
and2s1 U374 (.Q(N1093), .DIN1(N899), .DIN2(N1016));
and2s1 U375 (.Q(N1096), .DIN1(N925), .DIN2(N1021));
and2s1 U376 (.Q(N1099), .DIN1(N886), .DIN2(N1021));
and2s1 U377 (.Q(N1102), .DIN1(N912), .DIN2(N1021));
and2s1 U378 (.Q(N1105), .DIN1(N899), .DIN2(N1021));
and2s1 U379 (.Q(N1108), .DIN1(N925), .DIN2(N1026));
and2s1 U380 (.Q(N1111), .DIN1(N886), .DIN2(N1026));
and2s1 U381 (.Q(N1114), .DIN1(N912), .DIN2(N1026));
and2s1 U382 (.Q(N1117), .DIN1(N899), .DIN2(N1026));
and2s1 U383 (.Q(N1120), .DIN1(N925), .DIN2(N1031));
and2s1 U384 (.Q(N1123), .DIN1(N886), .DIN2(N1031));
and2s1 U385 (.Q(N1126), .DIN1(N912), .DIN2(N1031));
and2s1 U386 (.Q(N1129), .DIN1(N899), .DIN2(N1031));
nnd2s1 U387 (.Q(N1132), .DIN1(N1), .DIN2(N1036));
nnd2s1 U388 (.Q(N1135), .DIN1(N8), .DIN2(N1039));
nnd2s1 U389 (.Q(N1138), .DIN1(N15), .DIN2(N1042));
nnd2s1 U390 (.Q(N1141), .DIN1(N22), .DIN2(N1045));
nnd2s1 U391 (.Q(N1144), .DIN1(N29), .DIN2(N1048));
nnd2s1 U392 (.Q(N1147), .DIN1(N36), .DIN2(N1051));
nnd2s1 U393 (.Q(N1150), .DIN1(N43), .DIN2(N1054));
nnd2s1 U394 (.Q(N1153), .DIN1(N50), .DIN2(N1057));
nnd2s1 U395 (.Q(N1156), .DIN1(N57), .DIN2(N1060));
nnd2s1 U396 (.Q(N1159), .DIN1(N64), .DIN2(N1063));
nnd2s1 U397 (.Q(N1162), .DIN1(N71), .DIN2(N1066));
nnd2s1 U398 (.Q(N1165), .DIN1(N78), .DIN2(N1069));
nnd2s1 U399 (.Q(N1168), .DIN1(N85), .DIN2(N1072));
nnd2s1 U400 (.Q(N1171), .DIN1(N92), .DIN2(N1075));
nnd2s1 U401 (.Q(N1174), .DIN1(N99), .DIN2(N1078));
nnd2s1 U402 (.Q(N1177), .DIN1(N106), .DIN2(N1081));
nnd2s1 U403 (.Q(N1180), .DIN1(N113), .DIN2(N1084));
nnd2s1 U404 (.Q(N1183), .DIN1(N120), .DIN2(N1087));
nnd2s1 U405 (.Q(N1186), .DIN1(N127), .DIN2(N1090));
nnd2s1 U406 (.Q(N1189), .DIN1(N134), .DIN2(N1093));
nnd2s1 U407 (.Q(N1192), .DIN1(N141), .DIN2(N1096));
nnd2s1 U408 (.Q(N1195), .DIN1(N148), .DIN2(N1099));
nnd2s1 U409 (.Q(N1198), .DIN1(N155), .DIN2(N1102));
nnd2s1 U410 (.Q(N1201), .DIN1(N162), .DIN2(N1105));
nnd2s1 U411 (.Q(N1204), .DIN1(N169), .DIN2(N1108));
nnd2s1 U412 (.Q(N1207), .DIN1(N176), .DIN2(N1111));
nnd2s1 U413 (.Q(N1210), .DIN1(N183), .DIN2(N1114));
nnd2s1 U414 (.Q(N1213), .DIN1(N190), .DIN2(N1117));
nnd2s1 U415 (.Q(N1216), .DIN1(N197), .DIN2(N1120));
nnd2s1 U416 (.Q(N1219), .DIN1(N204), .DIN2(N1123));
nnd2s1 U417 (.Q(N1222), .DIN1(N211), .DIN2(N1126));
nnd2s1 U418 (.Q(N1225), .DIN1(N218), .DIN2(N1129));
nnd2s1 U419 (.Q(N1228), .DIN1(N1), .DIN2(N1132));
nnd2s1 U420 (.Q(N1229), .DIN1(N1036), .DIN2(N1132));
nnd2s1 U421 (.Q(N1230), .DIN1(N8), .DIN2(N1135));
nnd2s1 U422 (.Q(N1231), .DIN1(N1039), .DIN2(N1135));
nnd2s1 U423 (.Q(N1232), .DIN1(N15), .DIN2(N1138));
nnd2s1 U424 (.Q(N1233), .DIN1(N1042), .DIN2(N1138));
nnd2s1 U425 (.Q(N1234), .DIN1(N22), .DIN2(N1141));
nnd2s1 U426 (.Q(N1235), .DIN1(N1045), .DIN2(N1141));
nnd2s1 U427 (.Q(N1236), .DIN1(N29), .DIN2(N1144));
nnd2s1 U428 (.Q(N1237), .DIN1(N1048), .DIN2(N1144));
nnd2s1 U429 (.Q(N1238), .DIN1(N36), .DIN2(N1147));
nnd2s1 U430 (.Q(N1239), .DIN1(N1051), .DIN2(N1147));
nnd2s1 U431 (.Q(N1240), .DIN1(N43), .DIN2(N1150));
nnd2s1 U432 (.Q(N1241), .DIN1(N1054), .DIN2(N1150));
nnd2s1 U433 (.Q(N1242), .DIN1(N50), .DIN2(N1153));
nnd2s1 U434 (.Q(N1243), .DIN1(N1057), .DIN2(N1153));
nnd2s1 U435 (.Q(N1244), .DIN1(N57), .DIN2(N1156));
nnd2s1 U436 (.Q(N1245), .DIN1(N1060), .DIN2(N1156));
nnd2s1 U437 (.Q(N1246), .DIN1(N64), .DIN2(N1159));
nnd2s1 U438 (.Q(N1247), .DIN1(N1063), .DIN2(N1159));
nnd2s1 U439 (.Q(N1248), .DIN1(N71), .DIN2(N1162));
nnd2s1 U440 (.Q(N1249), .DIN1(N1066), .DIN2(N1162));
nnd2s1 U441 (.Q(N1250), .DIN1(N78), .DIN2(N1165));
nnd2s1 U442 (.Q(N1251), .DIN1(N1069), .DIN2(N1165));
nnd2s1 U443 (.Q(N1252), .DIN1(N85), .DIN2(N1168));
nnd2s1 U444 (.Q(N1253), .DIN1(N1072), .DIN2(N1168));
nnd2s1 U445 (.Q(N1254), .DIN1(N92), .DIN2(N1171));
nnd2s1 U446 (.Q(N1255), .DIN1(N1075), .DIN2(N1171));
nnd2s1 U447 (.Q(N1256), .DIN1(N99), .DIN2(N1174));
nnd2s1 U448 (.Q(N1257), .DIN1(N1078), .DIN2(N1174));
nnd2s1 U449 (.Q(N1258), .DIN1(N106), .DIN2(N1177));
nnd2s1 U450 (.Q(N1259), .DIN1(N1081), .DIN2(N1177));
nnd2s1 U451 (.Q(N1260), .DIN1(N113), .DIN2(N1180));
nnd2s1 U452 (.Q(N1261), .DIN1(N1084), .DIN2(N1180));
nnd2s1 U453 (.Q(N1262), .DIN1(N120), .DIN2(N1183));
nnd2s1 U454 (.Q(N1263), .DIN1(N1087), .DIN2(N1183));
nnd2s1 U455 (.Q(N1264), .DIN1(N127), .DIN2(N1186));
nnd2s1 U456 (.Q(N1265), .DIN1(N1090), .DIN2(N1186));
nnd2s1 U457 (.Q(N1266), .DIN1(N134), .DIN2(N1189));
nnd2s1 U458 (.Q(N1267), .DIN1(N1093), .DIN2(N1189));
nnd2s1 U459 (.Q(N1268), .DIN1(N141), .DIN2(N1192));
nnd2s1 U460 (.Q(N1269), .DIN1(N1096), .DIN2(N1192));
nnd2s1 U461 (.Q(N1270), .DIN1(N148), .DIN2(N1195));
nnd2s1 U462 (.Q(N1271), .DIN1(N1099), .DIN2(N1195));
nnd2s1 U463 (.Q(N1272), .DIN1(N155), .DIN2(N1198));
nnd2s1 U464 (.Q(N1273), .DIN1(N1102), .DIN2(N1198));
nnd2s1 U465 (.Q(N1274), .DIN1(N162), .DIN2(N1201));
nnd2s1 U466 (.Q(N1275), .DIN1(N1105), .DIN2(N1201));
nnd2s1 U467 (.Q(N1276), .DIN1(N169), .DIN2(N1204));
nnd2s1 U468 (.Q(N1277), .DIN1(N1108), .DIN2(N1204));
nnd2s1 U469 (.Q(N1278), .DIN1(N176), .DIN2(N1207));
nnd2s1 U470 (.Q(N1279), .DIN1(N1111), .DIN2(N1207));
nnd2s1 U471 (.Q(N1280), .DIN1(N183), .DIN2(N1210));
nnd2s1 U472 (.Q(N1281), .DIN1(N1114), .DIN2(N1210));
nnd2s1 U473 (.Q(N1282), .DIN1(N190), .DIN2(N1213));
nnd2s1 U474 (.Q(N1283), .DIN1(N1117), .DIN2(N1213));
nnd2s1 U475 (.Q(N1284), .DIN1(N197), .DIN2(N1216));
nnd2s1 U476 (.Q(N1285), .DIN1(N1120), .DIN2(N1216));
nnd2s1 U477 (.Q(N1286), .DIN1(N204), .DIN2(N1219));
nnd2s1 U478 (.Q(N1287), .DIN1(N1123), .DIN2(N1219));
nnd2s1 U479 (.Q(N1288), .DIN1(N211), .DIN2(N1222));
nnd2s1 U480 (.Q(N1289), .DIN1(N1126), .DIN2(N1222));
nnd2s1 U481 (.Q(N1290), .DIN1(N218), .DIN2(N1225));
nnd2s1 U482 (.Q(N1291), .DIN1(N1129), .DIN2(N1225));
nnd2s1 U483 (.Q(N1292), .DIN1(N1228), .DIN2(N1229));
nnd2s1 U484 (.Q(N1293), .DIN1(N1230), .DIN2(N1231));
nnd2s1 U485 (.Q(N1294), .DIN1(N1232), .DIN2(N1233));
nnd2s1 U486 (.Q(N1295), .DIN1(N1234), .DIN2(N1235));
nnd2s1 U487 (.Q(N1296), .DIN1(N1236), .DIN2(N1237));
nnd2s1 U488 (.Q(N1297), .DIN1(N1238), .DIN2(N1239));
nnd2s1 U489 (.Q(N1298), .DIN1(N1240), .DIN2(N1241));
nnd2s1 U490 (.Q(N1299), .DIN1(N1242), .DIN2(N1243));
nnd2s1 U491 (.Q(N1300), .DIN1(N1244), .DIN2(N1245));
nnd2s1 U492 (.Q(N1301), .DIN1(N1246), .DIN2(N1247));
nnd2s1 U493 (.Q(N1302), .DIN1(N1248), .DIN2(N1249));
nnd2s1 U494 (.Q(N1303), .DIN1(N1250), .DIN2(N1251));
nnd2s1 U495 (.Q(N1304), .DIN1(N1252), .DIN2(N1253));
nnd2s1 U496 (.Q(N1305), .DIN1(N1254), .DIN2(N1255));
nnd2s1 U497 (.Q(N1306), .DIN1(N1256), .DIN2(N1257));
nnd2s1 U498 (.Q(N1307), .DIN1(N1258), .DIN2(N1259));
nnd2s1 U499 (.Q(N1308), .DIN1(N1260), .DIN2(N1261));
nnd2s1 U500 (.Q(N1309), .DIN1(N1262), .DIN2(N1263));
nnd2s1 U501 (.Q(N1310), .DIN1(N1264), .DIN2(N1265));
nnd2s1 U502 (.Q(N1311), .DIN1(N1266), .DIN2(N1267));
nnd2s1 U503 (.Q(N1312), .DIN1(N1268), .DIN2(N1269));
nnd2s1 U504 (.Q(N1313), .DIN1(N1270), .DIN2(N1271));
nnd2s1 U505 (.Q(N1314), .DIN1(N1272), .DIN2(N1273));
nnd2s1 U506 (.Q(N1315), .DIN1(N1274), .DIN2(N1275));
nnd2s1 U507 (.Q(N1316), .DIN1(N1276), .DIN2(N1277));
nnd2s1 U508 (.Q(N1317), .DIN1(N1278), .DIN2(N1279));
nnd2s1 U509 (.Q(N1318), .DIN1(N1280), .DIN2(N1281));
nnd2s1 U510 (.Q(N1319), .DIN1(N1282), .DIN2(N1283));
nnd2s1 U511 (.Q(N1320), .DIN1(N1284), .DIN2(N1285));
nnd2s1 U512 (.Q(N1321), .DIN1(N1286), .DIN2(N1287));
nnd2s1 U513 (.Q(N1322), .DIN1(N1288), .DIN2(N1289));
nnd2s1 U514 (.Q(N1323), .DIN1(N1290), .DIN2(N1291));
nb1s1 U515 (.Q(N1324), .DIN(N1292));
nb1s1 U516 (.Q(N1325), .DIN(N1293));
nb1s1 U517 (.Q(N1326), .DIN(N1294));
nb1s1 U518 (.Q(N1327), .DIN(N1295));
nb1s1 U519 (.Q(N1328), .DIN(N1296));
nb1s1 U520 (.Q(N1329), .DIN(N1297));
nb1s1 U521 (.Q(N1330), .DIN(N1298));
nb1s1 U522 (.Q(N1331), .DIN(N1299));
nb1s1 U523 (.Q(N1332), .DIN(N1300));
nb1s1 U524 (.Q(N1333), .DIN(N1301));
nb1s1 U525 (.Q(N1334), .DIN(N1302));
nb1s1 U526 (.Q(N1335), .DIN(N1303));
nb1s1 U527 (.Q(N1336), .DIN(N1304));
nb1s1 U528 (.Q(N1337), .DIN(N1305));
nb1s1 U529 (.Q(N1338), .DIN(N1306));
nb1s1 U530 (.Q(N1339), .DIN(N1307));
nb1s1 U531 (.Q(N1340), .DIN(N1308));
nb1s1 U532 (.Q(N1341), .DIN(N1309));
nb1s1 U533 (.Q(N1342), .DIN(N1310));
nb1s1 U534 (.Q(N1343), .DIN(N1311));
nb1s1 U535 (.Q(N1344), .DIN(N1312));
nb1s1 U536 (.Q(N1345), .DIN(N1313));
nb1s1 U537 (.Q(N1346), .DIN(N1314));
nb1s1 U538 (.Q(N1347), .DIN(N1315));
nb1s1 U539 (.Q(N1348), .DIN(N1316));
nb1s1 U540 (.Q(N1349), .DIN(N1317));
nb1s1 U541 (.Q(N1350), .DIN(N1318));
nb1s1 U542 (.Q(N1351), .DIN(N1319));
nb1s1 U543 (.Q(N1352), .DIN(N1320));
nb1s1 U544 (.Q(N1353), .DIN(N1321));
nb1s1 U545 (.Q(N1354), .DIN(N1322));
nb1s1 U546 (.Q(N1355), .DIN(N1323));
endmodule
