module mc ( clk_i, rst_i, wb_data_i, wb_data_o, wb_addr_i, wb_sel_i, 
        wb_we_i, wb_cyc_i, wb_stb_i, wb_ack_o, wb_err_o, susp_req_i, 
        resume_req_i, suspended_o, poc_o, mc_clk_i, mc_br_pad_i, mc_bg_pad_o, 
        mc_ack_pad_i, mc_addr_pad_o, mc_data_pad_i, mc_data_pad_o, mc_dp_pad_i, 
        mc_dp_pad_o, mc_doe_pad_doe_o, mc_dqm_pad_o, mc_oe_pad_o_, 
        mc_we_pad_o_, mc_cas_pad_o_, mc_ras_pad_o_, mc_cke_pad_o_, 
        mc_cs_pad_o_, mc_sts_pad_i, mc_rp_pad_o_, mc_vpen_pad_o, 
        mc_adsc_pad_o_, mc_adv_pad_o_, mc_zz_pad_o, mc_coe_pad_coe_o );
  input [31:0] wb_data_i;
  output [31:0] wb_data_o;
  input [31:0] wb_addr_i;
  input [3:0] wb_sel_i;
  output [31:0] poc_o;
  output [23:0] mc_addr_pad_o;
  input [31:0] mc_data_pad_i;
  output [31:0] mc_data_pad_o;
  input [3:0] mc_dp_pad_i;
  output [3:0] mc_dp_pad_o;
  output [3:0] mc_dqm_pad_o;
  output [7:0] mc_cs_pad_o_;
  input clk_i, rst_i, wb_we_i, wb_cyc_i, wb_stb_i, susp_req_i, resume_req_i,
         mc_clk_i, mc_br_pad_i, mc_ack_pad_i, mc_sts_pad_i;
  output wb_ack_o, wb_err_o, suspended_o, mc_bg_pad_o, mc_doe_pad_doe_o,
         mc_oe_pad_o_, mc_we_pad_o_, mc_cas_pad_o_, mc_ras_pad_o_,
         mc_cke_pad_o_, mc_rp_pad_o_, mc_vpen_pad_o, mc_adsc_pad_o_,
         mc_adv_pad_o_, mc_zz_pad_o, mc_coe_pad_coe_o;
  wire   \u5_temp_cs[1] , u5_cs_le, u0_csc_10, u0_csc_9, u0_sp_csc_10,
         u0_sp_csc_9, u5_init_ack, u5_lmr_ack, u0_init_req, N872, N873, N874,
         N875, N876, N877, N878, N879, N880, N881, N882, N883, N884,
         \u1_u0_out_r[12] , u5_susp_sel_r, u5_mem_ack_r, u5_dv, N1549,
         u4_rfr_req, rfr_ack, u5_cmd_asserted2, u5_cke_r, u5_wb_wait_r,
         u5_wb_cycle, u5_cnt, u5_resume_req_r, u5_suspended_d, u5_tmr2_done,
         u5_tmr_done, u5_ap_en, u5_wb_write_go_r, u5_wb_stb_first, u7_mc_br_r,
         n4530, n4531, n4532, n4533, n4535, n4536, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4611, n4612,
         n4616, n4618, n4625, n4629, n4770, n4771, n4814, n4820, n4975, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n5504, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9180, n9182, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9677, n9678, n9679, n9680, n9682, n9683, n9684, n9685, n9686, n9688,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9764, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n15470, n15471, n15472,
         n15473, n15474, n15475, n15477, n15478, n15479, n15481, n15482,
         n15483, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15521, n15523,
         n19404, n19405, n19406, n19407, n19409, n19410, n19411, n19412,
         n19413, n9689, u5_rsts, u5_rfr_ack_d, n9924, n9923, n9922, n9860,
         n9765, n9763, n9681, n9676, n9675, n9532, n9196, n9183, n9181, n9179,
         n5503, n5499, n5496, n5495, n5492, n5491, n5487, n5484, n5483, n5477,
         n5476, n5471, n5470, n5465, n5464, n5458, n5453, n5452, n5448, n5446,
         n5445, n5441, n5439, n5438, n5434, n5432, n5431, n5428, n5427, n5424,
         n5423, n5420, n5419, n5416, n5415, n5412, n5411, n5408, n5407, n5404,
         n5403, n5400, n5399, n5396, n5395, n5392, n5391, n5388, n5387, n5384,
         n5383, n5380, n5379, n5376, n5375, n5372, n5371, n5368, n5367, n5364,
         n5363, n5360, n5359, n5356, n5355, n5352, n5351, n5348, n5347, n5344,
         n5343, n5340, n5339, n5336, n5335, n5332, n5331, n5328, n5327, n5324,
         n5323, n5320, n5319, n5316, n5315, n5312, n5311, n5308, n5307, n5304,
         n5303, n5300, n5299, n5296, n5295, n5292, n5291, n5288, n5287, n5284,
         n5283, n5280, n5279, n5276, n5275, n5272, n5271, n5268, n5267, n5264,
         n5263, n5260, n5259, n5256, n5255, n5252, n5251, n5248, n5247, n5244,
         n5243, n5240, n5239, n5236, n5235, n5232, n5231, n5228, n5227, n5224,
         n5223, n5220, n5219, n5216, n5215, n5212, n5211, n5208, n5207, n5204,
         n5203, n5200, n5199, n5196, n5195, n5192, n5191, n5188, n5187, n5184,
         n5183, n5180, n5179, n5176, n5175, n4529, n19408, n19403, n19402,
         n19401, n15531, n15530, n15529, n15528, n15527, n15526, n15525,
         n31021, n31022, n31023, n31024, n31025, n31026, n31027, n31028,
         n31029, n31030, n31031, n31032, n31033, n31034, n31035, n31036,
         n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044,
         n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052,
         n31053, n31054, n31055, n31056, n31057, n31058, n31059, n31060,
         n31061, n31062, n31063, n31064, n31065, n31066, n31067, n31068,
         n31069, n31070, n31071, n31072, n31073, n31074, n31075, n31076,
         n31077, n31078, n31079, n31080, n31081, n31082, n31083, n31084,
         n31085, n31086, n31087, n31088, n31089, n31090, n31091, n31092,
         n31093, n31094, n31095, n31096, n31097, n31098, n31099, n31100,
         n31101, n31102, n31103, n31104, n31105, n31106, n31107, n31108,
         n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116,
         n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124,
         n31125, n31126, n31127, n31128, n31129, n31130, n31131, n31132,
         n31133, n31134, n31135, n31136, n31137, n31138, n31139, n31140,
         n31141, n31142, n31143, n31144, n31145, n31146, n31147, n31148,
         n31149, n31150, n31151, n31152, n31153, n31154, n31155, n31156,
         n31157, n31158, n31159, n31160, n31161, n31162, n31163, n31164,
         n31165, n31166, n31167, n31168, n31169, n31170, n31171, n31172,
         n31173, n31174, n31175, n31176, n31177, n31178, n31179, n31180,
         n31181, n31182, n31183, n31184, n31185, n31186, n31187, n31188,
         n31189, n31190, n31191, n31192, n31193, n31194, n31195, n31196,
         n31197, n31198, n31199, n31200, n31201, n31202, n31203, n31204,
         n31205, n31206, n31207, n31208, n31209, n31210, n31211, n31212,
         n31213, n31214, n31215, n31216, n31217, n31218, n31219, n31220,
         n31221, n31222, n31223, n31224, n31225, n31226, n31227, n31228,
         n31229, n31230, n31231, n31232, n31233, n31234, n31235, n31236,
         n31237, n31238, n31239, n31240, n31241, n31242, n31243, n31244,
         n31245, n31246, n31247, n31248, n31249, n31250, n31251, n31252,
         n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260,
         n31261, n31262, n31263, n31264, n31265, n31266, n31267, n31268,
         n31269, n31270, n31271, n31272, n31273, n31274, n31275, n31276,
         n31277, n31278, n31279, n31280, n31281, n31282, n31283, n31284,
         n31285, n31286, n31287, n31288, n31289, n31290, n31291, n31292,
         n31293, n31294, n31295, n31296, n31297, n31298, n31299, n31300,
         n31301, n31302, n31303, n31304, n31305, n31306, n31307, n31308,
         n31309, n31310, n31311, n31312, n31313, n31314, n31315, n31316,
         n31317, n31318, n31319, n31320, n31321, n31322, n31323, n31324,
         n31325, n31326, n31327, n31328, n31329, n31330, n31331, n31332,
         n31333, n31334, n31335, n31336, n31337, n31338, n31339, n31340,
         n31341, n31342, n31343, n31344, n31345, n31346, n31347, n31348,
         n31349, n31350, n31351, n31352, n31353, n31354, n31355, n31356,
         n31357, n31358, n31359, n31360, n31361, n31362, n31363, n31364,
         n31365, n31366, n31367, n31368, n31369, n31370, n31371, n31372,
         n31373, n31374, n31375, n31376, n31377, n31378, n31379, n31380,
         n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388,
         n31389, n31390, n31391, n31392, n31393, n31394, n31395, n31396,
         n31397, n31398, n31399, n31400, n31401, n31402, n31403, n31404,
         n31405, n31406, n31407, n31408, n31409, n31410, n31411, n31412,
         n31413, n31414, n31415, n31416, n31417, n31418, n31419, n31420,
         n31421, n31422, n31423, n31424, n31425, n31426, n31427, n31428,
         n31429, n31430, n31431, n31432, n31433, n31434, n31435, n31436,
         n31437, n31438, n31439, n31440, n31441, n31442, n31443, n31444,
         n31445, n31446, n31447, n31448, n31449, n31450, n31451, n31452,
         n31453, n31454, n31455, n31456, n31457, n31458, n31459, n31460,
         n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468,
         n31469, n31470, n31471, n31472, n31473, n31474, n31475, n31476,
         n31477, n31478, n31479, n31480, n31481, n31482, n31483, n31484,
         n31485, n31486, n31487, n31488, n31489, n31490, n31491, n31492,
         n31493, n31494, n31495, n31496, n31497, n31498, n31499, n31500,
         n31501, n31502, n31503, n31504, n31505, n31506, n31507, n31508,
         n31509, n31510, n31511, n31512, n31513, n31514, n31515, n31516,
         n31517, n31518, n31519, n31520, n31521, n31522, n31523, n31524,
         n31525, n31526, n31527, n31528, n31529, n31530, n31531, n31532,
         n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540,
         n31541, n31542, n31543, n31544, n31545, n31546, n31547, n31548,
         n31549, n31550, n31551, n31552, n31553, n31554, n31555, n31556,
         n31557, n31558, n31559, n31560, n31561, n31562, n31563, n31564,
         n31565, n31566, n31567, n31568, n31569, n31570, n31571, n31572,
         n31573, n31574, n31575, n31576, n31577, n31578, n31579, n31580,
         n31581, n31582, n31583, n31584, n31585, n31586, n31587, n31588,
         n31589, n31590, n31591, n31592, n31593, n31594, n31595, n31596,
         n31597, n31598, n31599, n31600, n31601, n31602, n31603, n31604,
         n31605, n31606, n31607, n31608, n31609, n31610, n31611, n31612,
         n31613, n31614, n31615, n31616, n31617, n31618, n31619, n31620,
         n31621, n31622, n31623, n31624, n31625, n31626, n31627, n31628,
         n31629, n31630, n31631, n31632, n31633, n31634, n31635, n31636,
         n31637, n31638, n31639, n31640, n31641, n31642, n31643, n31644,
         n31645, n31646, n31647, n31648, n31649, n31650, n31651, n31652,
         n31653, n31654, n31655, n31656, n31657, n31658, n31659, n31660,
         n31661, n31662, n31663, n31664, n31665, n31666, n31667, n31668,
         n31669, n31670, n31671, n31672, n31673, n31674, n31675, n31676,
         n31677, n31678, n31679, n31680, n31681, n31682, n31683, n31684,
         n31685, n31686, n31687, n31688, n31689, n31690, n31691, n31692,
         n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700,
         n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708,
         n31709, n31710, n31711, n31712, n31713, n31714, n31715, n31716,
         n31717, n31718, n31719, n31720, n31721, n31722, n31723, n31724,
         n31725, n31726, n31727, n31728, n31729, n31730, n31731, n31732,
         n31733, n31734, n31735, n31736, n31737, n31738, n31739, n31740,
         n31741, n31742, n31743, n31744, n31745, n31746, n31747, n31748,
         n31749, n31750, n31751, n31752, n31753, n31754, n31755, n31756,
         n31757, n31758, n31759, n31760, n31761, n31762, n31763, n31764,
         n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772,
         n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780,
         n31781, n31782, n31783, n31784, n31785, n31786, n31787, n31788,
         n31789, n31790, n31791, n31792, n31793, n31794, n31795, n31796,
         n31797, n31798, n31799, n31800, n31801, n31802, n31803, n31804,
         n31805, n31806, n31807, n31808, n31809, n31810, n31811, n31812,
         n31813, n31814, n31815, n31816, n31817, n31818, n31819, n31820,
         n31821, n31822, n31823, n31824, n31825, n31826, n31827, n31828,
         n31829, n31830, n31831, n31832, n31833, n31834, n31835, n31836,
         n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844,
         n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852,
         n31853, n31854, n31855, n31856, n31857, n31858, n31859, n31860,
         n31861, n31862, n31863, n31864, n31865, n31866, n31867, n31868,
         n31869, n31870, n31871, n31872, n31873, n31874, n31875, n31876,
         n31877, n31878, n31879, n31880, n31881, n31882, n31883, n31884,
         n31885, n31886, n31887, n31888, n31889, n31890, n31891, n31892,
         n31893, n31894, n31895, n31896, n31897, n31898, n31899, n31900,
         n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908,
         n31909, n31910, n31911, n31912, n31913, n31914, n31915, n31916,
         n31917, n31918, n31919, n31920, n31921, n31922, n31923, n31924,
         n31925, n31926, n31927, n31928, n31929, n31930, n31931, n31932,
         n31933, n31934, n31935, n31936, n31937, n31938, n31939, n31940,
         n31941, n31942, n31943, n31944, n31945, n31946, n31947, n31948,
         n31949, n31950, n31951, n31952, n31953, n31954, n31955, n31956,
         n31957, n31958, n31959, n31960, n31961, n31962, n31963, n31964,
         n31965, n31966, n31967, n31968, n31969, n31970, n31971, n31972,
         n31973, n31974, n31975, n31976, n31977, n31978, n31979, n31980,
         n31981, n31982, n31983, n31984, n31985, n31986, n31987, n31988,
         n31989, n31990, n31991, n31992, n31993, n31994, n31995, n31996,
         n31997, n31998, n31999, n32000, n32001, n32002, n32003, n32004,
         n32005, n32006, n32007, n32008, n32009, n32010, n32011, n32012,
         n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020,
         n32021, n32022, n32023, n32024, n32025, n32026, n32027, n32028,
         n32029, n32030, n32031, n32032, n32033, n32034, n32035, n32036,
         n32037, n32038, n32039, n32040, n32041, n32042, n32043, n32044,
         n32045, n32046, n32047, n32048, n32049, n32050, n32051, n32052,
         n32053, n32054, n32055, n32056, n32057, n32058, n32059, n32060,
         n32061, n32062, n32063, n32064, n32065, n32066, n32067, n32068,
         n32069, n32070, n32071, n32072, n32073, n32074, n32075, n32076,
         n32077, n32078, n32079, n32080, n32081, n32082, n32083, n32084,
         n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092,
         n32093, n32094, n32095, n32096, n32097, n32098, n32099, n32100,
         n32101, n32102, n32103, n32104, n32105, n32106, n32107, n32108,
         n32109, n32110, n32111, n32112, n32113, n32114, n32115, n32116,
         n32117, n32118, n32119, n32120, n32121, n32122, n32123, n32124,
         n32125, n32126, n32127, n32128, n32129, n32130, n32131, n32132,
         n32133, n32134, n32135, n32136, n32137, n32138, n32139, n32140,
         n32141, n32142, n32143, n32144, n32145, n32146, n32147, n32148,
         n32149, n32150, n32151, n32152, n32153, n32154, n32155, n32156,
         n32157, n32158, n32159, n32160, n32161, n32162, n32163, n32164,
         n32165, n32166, n32167, n32168, n32169, n32170, n32171, n32172,
         n32173, n32174, n32175, n32176, n32177, n32178, n32179, n32180,
         n32181, n32182, n32183, n32184, n32185, n32186, n32187, n32188,
         n32189, n32190, n32191, n32192, n32193, n32194, n32195, n32196,
         n32197, n32198, n32199, n32200, n32201, n32202, n32203, n32204,
         n32205, n32206, n32207, n32208, n32209, n32210, n32211, n32212,
         n32213, n32214, n32215, n32216, n32217, n32218, n32219, n32220,
         n32221, n32222, n32223, n32224, n32225, n32226, n32227, n32228,
         n32229, n32230, n32231, n32232, n32233, n32234, n32235, n32236,
         n32237, n32238, n32239, n32240, n32241, n32242, n32243, n32244,
         n32245, n32246, n32247, n32248, n32249, n32250, n32251, n32252,
         n32253, n32254, n32255, n32256, n32257, n32258, n32259, n32260,
         n32261, n32262, n32263, n32264, n32265, n32266, n32267, n32268,
         n32269, n32270, n32271, n32272, n32273, n32274, n32275, n32276,
         n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284,
         n32285, n32286, n32287, n32288, n32289, n32290, n32291, n32292,
         n32293, n32294, n32295, n32296, n32297, n32298, n32299, n32300,
         n32301, n32302, n32303, n32304, n32305, n32306, n32307, n32308,
         n32309, n32310, n32311, n32312, n32313, n32314, n32315, n32316,
         n32317, n32318, n32319, n32320, n32321, n32322, n32323, n32324,
         n32325, n32326, n32327, n32328, n32329, n32330, n32331, n32332,
         n32333, n32334, n32335, n32336, n32337, n32338, n32339, n32340,
         n32341, n32342, n32343, n32344, n32345, n32346, n32347, n32348,
         n32349, n32350, n32351, n32352, n32353, n32354, n32355, n32356,
         n32357, n32358, n32359, n32360, n32361, n32362, n32363, n32364,
         n32365, n32366, n32367, n32368, n32369, n32370, n32371, n32372,
         n32373, n32374, n32375, n32376, n32377, n32378, n32379, n32380,
         n32381, n32382, n32383, n32384, n32385, n32386, n32387, n32388,
         n32389, n32390, n32391, n32392, n32393, n32394, n32395, n32396,
         n32397, n32398, n32399, n32400, n32401, n32402, n32403, n32404,
         n32405, n32406, n32407, n32408, n32409, n32410, n32411, n32412,
         n32413, n32414, n32415, n32416, n32417, n32418, n32419, n32420,
         n32421, n32422, n32423, n32424, n32425, n32426, n32427, n32428,
         n32429, n32430, n32431, n32432, n32433, n32434, n32435, n32436,
         n32437, n32438, n32439, n32440, n32441, n32442, n32443, n32444,
         n32445, n32446, n32447, n32448, n32449, n32450, n32451, n32452,
         n32453, n32454, n32455, n32456, n32457, n32458, n32459, n32460,
         n32461, n32462, n32463, n32464, n32465, n32466, n32467, n32468,
         n32469, n32470, n32471, n32472, n32473, n32474, n32475, n32476,
         n32477, n32478, n32479, n32480, n32481, n32482, n32483, n32484,
         n32485, n32486, n32487, n32488, n32489, n32490, n32491, n32492,
         n32493, n32494, n32495, n32496, n32497, n32498, n32499, n32500,
         n32501, n32502, n32503, n32504, n32505, n32506, n32507, n32508,
         n32509, n32510, n32511, n32512, n32513, n32514, n32515, n32516,
         n32517, n32518, n32519, n32520, n32521, n32522, n32523, n32524,
         n32525, n32526, n32527, n32528, n32529, n32530, n32531, n32532,
         n32533, n32534, n32535, n32536, n32537, n32538, n32539, n32540,
         n32541, n32542, n32543, n32544, n32545, n32546, n32547, n32548,
         n32549, n32550, n32551, n32552, n32553, n32554, n32555, n32556,
         n32557, n32558, n32559, n32560, n32561, n32562, n32563, n32564,
         n32565, n32566, n32567, n32568, n32569, n32570, n32571, n32572,
         n32573, n32574, n32575, n32576, n32577, n32578, n32579, n32580,
         n32581, n32582, n32583, n32584, n32585, n32586, n32587, n32588,
         n32589, n32590, n32591, n32592, n32593, n32594, n32595, n32596,
         n32597, n32598, n32599, n32600, n32601, n32602, n32603, n32604,
         n32605, n32606, n32607, n32608, n32609, n32610, n32611, n32612,
         n32613, n32614, n32615, n32616, n32617, n32618, n32619, n32620,
         n32621, n32622, n32623, n32624, n32625, n32626, n32627, n32628,
         n32629, n32630, n32631, n32632, n32633, n32634, n32635, n32636,
         n32637, n32638, n32639, n32640, n32641, n32642, n32643, n32644,
         n32645, n32646, n32647, n32648, n32649, n32650, n32651, n32652,
         n32653, n32654, n32655, n32656, n32657, n32658, n32659, n32660,
         n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668,
         n32669, n32670, n32671, n32672, n32673, n32674, n32675, n32676,
         n32677, n32678, n32679, n32680, n32681, n32682, n32683, n32684,
         n32685, n32686, n32687, n32688, n32689, n32690, n32691, n32692,
         n32693, n32694, n32695, n32696, n32697, n32698, n32699, n32700,
         n32701, n32702, n32703, n32704, n32705, n32706, n32707, n32708,
         n32709, n32710, n32711, n32712, n32713, n32714, n32715, n32716,
         n32717, n32718, n32719, n32720, n32721, n32722, n32723, n32724,
         n32725, n32726, n32727, n32728, n32729, n32730, n32731, n32732,
         n32733, n32734, n32735, n32736, n32737, n32738, n32739, n32740,
         n32741, n32742, n32743, n32744, n32745, n32746, n32747, n32748,
         n32749, n32750, n32751, n32752, n32753, n32754, n32755, n32756,
         n32757, n32758, n32759, n32760, n32761, n32762, n32763, n32764,
         n32765, n32766, n32767, n32768, n32769, n32770, n32771, n32772,
         n32773, n32774, n32775, n32776, n32777, n32778, n32779, n32780,
         n32781, n32782, n32783, n32784, n32785, n32786, n32787, n32788,
         n32789, n32790, n32791, n32792, n32793, n32794, n32795, n32796,
         n32797, n32798, n32799, n32800, n32801, n32802, n32803, n32804,
         n32805, n32806, n32807, n32808, n32809, n32810, n32811, n32812,
         n32813, n32814, n32815, n32816, n32817, n32818, n32819, n32820,
         n32821, n32822, n32823, n32824, n32825, n32826, n32827, n32828,
         n32829, n32830, n32831, n32832, n32833, n32834, n32835, n32836,
         n32837, n32838, n32839, n32840, n32841, n32842, n32843, n32844,
         n32845, n32846, n32847, n32848, n32849, n32850, n32851, n32852,
         n32853, n32854, n32855, n32856, n32857, n32858, n32859, n32860,
         n32861, n32862, n32863, n32864, n32865, n32866, n32867, n32868,
         n32869, n32870, n32871, n32872, n32873, n32874, n32875, n32876,
         n32877, n32878, n32879, n32880, n32881, n32882, n32883, n32884,
         n32885, n32886, n32887, n32888, n32889, n32890, n32891, n32892,
         n32893, n32894, n32895, n32896, n32897, n32898, n32899, n32900,
         n32901, n32902, n32903, n32904, n32905, n32906, n32907, n32908,
         n32909, n32910, n32911, n32912, n32913, n32914, n32915, n32916,
         n32917, n32918, n32919, n32920, n32921, n32922, n32923, n32924,
         n32925, n32926, n32927, n32928, n32929, n32930, n32931, n32932,
         n32933, n32934, n32935, n32936, n32937, n32938, n32939, n32940,
         n32941, n32942, n32943, n32944, n32945, n32946, n32947, n32948,
         n32949, n32950, n32951, n32952, n32953, n32954, n32955, n32956,
         n32957, n32958, n32959, n32960, n32961, n32962, n32963, n32964,
         n32965, n32966, n32967, n32968, n32969, n32970, n32971, n32972,
         n32973, n32974, n32975, n32976, n32977, n32978, n32979, n32980,
         n32981, n32982, n32983, n32984, n32985, n32986, n32987, n32988,
         n32989, n32990, n32991, n32992, n32993, n32994, n32995, n32996,
         n32997, n32998, n32999, n33000, n33001, n33002, n33003, n33004,
         n33005, n33006, n33007, n33008, n33009, n33010, n33011, n33012,
         n33013, n33014, n33015, n33016, n33017, n33018, n33019, n33020,
         n33021, n33022, n33023, n33024, n33025, n33026, n33027, n33028,
         n33029, n33030, n33031, n33032, n33033, n33034, n33035, n33036,
         n33037, n33038, n33039, n33040, n33041, n33042, n33043, n33044,
         n33045, n33046, n33047, n33048, n33049, n33050, n33051, n33052,
         n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060,
         n33061, n33062, n33063, n33064, n33065, n33066, n33067, n33068,
         n33069, n33070, n33071, n33072, n33073, n33074, n33075, n33076,
         n33077, n33078, n33079, n33080, n33081, n33082, n33083, n33084,
         n33085, n33086, n33087, n33088, n33089, n33090, n33091, n33092,
         n33093, n33094, n33095, n33096, n33097, n33098, n33099, n33100,
         n33101, n33102, n33103, n33104, n33105, n33106, n33107, n33108,
         n33109, n33110, n33111, n33112, n33113, n33114, n33115, n33116,
         n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33124,
         n33125, n33126, n33127, n33128, n33129, n33130, n33131, n33132,
         n33133, n33134, n33135, n33136, n33137, n33138, n33139, n33140,
         n33141, n33142, n33143, n33144, n33145, n33146, n33147, n33148,
         n33149, n33150, n33151, n33152, n33153, n33154, n33155, n33156,
         n33157, n33158, n33159, n33160, n33161, n33162, n33163, n33164,
         n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172,
         n33173, n33174, n33175, n33176, n33177, n33178, n33179, n33180,
         n33181, n33182, n33183, n33184, n33185, n33186, n33187, n33188,
         n33189, n33190, n33191, n33192, n33193, n33194, n33195, n33196,
         n33197, n33198, n33199, n33200, n33201, n33202, n33203, n33204,
         n33205, n33206, n33207, n33208, n33209, n33210, n33211, n33212,
         n33213, n33214, n33215, n33216, n33217, n33218, n33219, n33220,
         n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228,
         n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236,
         n33237, n33238, n33239, n33240, n33241, n33242, n33243, n33244,
         n33245, n33246, n33247, n33248, n33249, n33250, n33251, n33252,
         n33253, n33254, n33255, n33256, n33257, n33258, n33259, n33260,
         n33261, n33262, n33263, n33264, n33265, n33266, n33267, n33268,
         n33269, n33270, n33271, n33272, n33273, n33274, n33275, n33276,
         n33277, n33278, n33279, n33280, n33281, n33282, n33283, n33284,
         n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292,
         n33293, n33294, n33295, n33296, n33297, n33298, n33299, n33300,
         n33301, n33302, n33303, n33304, n33305, n33306, n33307, n33308,
         n33309, n33310, n33311, n33312, n33313, n33314, n33315, n33316,
         n33317, n33318, n33319, n33320, n33321, n33322, n33323, n33324,
         n33325, n33326, n33327, n33328, n33329, n33330, n33331, n33332,
         n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33340,
         n33341, n33342, n33343, n33344, n33345, n33346, n33347, n33348,
         n33349, n33350, n33351, n33352, n33353, n33354, n33355, n33356,
         n33357, n33358, n33359, n33360, n33361, n33362, n33363, n33364,
         n33365, n33366, n33367, n33368, n33369, n33370, n33371, n33372,
         n33373, n33374, n33375, n33376, n33377, n33378, n33379, n33380,
         n33381, n33382, n33383, n33384, n33385, n33386, n33387, n33388,
         n33389, n33390, n33391, n33392, n33393, n33394, n33395, n33396,
         n33397, n33398, n33399, n33400, n33401, n33402, n33403, n33404,
         n33405, n33406, n33407, n33408, n33409, n33410, n33411, n33412,
         n33413, n33414, n33415, n33416, n33417, n33418, n33419, n33420,
         n33421, n33422, n33423, n33424, n33425, n33426, n33427, n33428,
         n33429, n33430, n33431, n33432, n33433, n33434, n33435, n33436,
         n33437, n33438, n33439, n33440, n33441, n33442, n33443, n33444,
         n33445, n33446, n33447, n33448, n33449, n33450, n33451, n33452,
         n33453, n33454, n33455, n33456, n33457, n33458, n33459, n33460,
         n33461, n33462, n33463, n33464, n33465, n33466, n33467, n33468,
         n33469, n33470, n33471, n33472, n33473, n33474, n33475, n33476,
         n33477, n33478, n33479, n33480, n33481, n33482, n33483, n33484,
         n33485, n33486, n33487, n33488, n33489, n33490, n33491, n33492,
         n33493, n33494, n33495, n33496, n33497, n33498, n33499, n33500,
         n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508,
         n33509, n33510, n33511, n33512, n33513, n33514, n33515, n33516,
         n33517, n33518, n33519, n33520, n33521, n33522, n33523, n33524,
         n33525, n33526, n33527, n33528, n33529, n33530, n33531, n33532,
         n33533, n33534, n33535, n33536, n33537, n33538, n33539, n33540,
         n33541, n33542, n33543, n33544, n33545, n33546, n33547, n33548,
         n33549, n33550, n33551, n33552, n33553, n33554, n33555, n33556,
         n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564,
         n33565, n33566, n33567, n33568, n33569, n33570, n33571, n33572,
         n33573, n33574, n33575, n33576, n33577, n33578, n33579, n33580,
         n33581, n33582, n33583, n33584, n33585, n33586, n33587, n33588,
         n33589, n33590, n33591, n33592, n33593, n33594, n33595, n33596,
         n33597, n33598, n33599, n33600, n33601, n33602, n33603, n33604,
         n33605, n33606, n33607, n33608, n33609, n33610, n33611, n33612,
         n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620,
         n33621, n33622, n33623, n33624, n33625, n33626, n33627, n33628,
         n33629, n33630, n33631, n33632, n33633, n33634, n33635, n33636,
         n33637, n33638, n33639, n33640, n33641, n33642, n33643, n33644,
         n33645, n33646, n33647, n33648, n33649, n33650, n33651, n33652,
         n33653, n33654, n33655, n33656, n33657, n33658, n33659, n33660,
         n33661, n33662, n33663, n33664, n33665, n33666, n33667, n33668,
         n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676,
         n33677, n33678, n33679, n33680, n33681, n33682, n33683, n33684,
         n33685, n33686, n33687, n33688, n33689, n33690, n33691, n33692,
         n33693, n33694, n33695, n33696, n33697, n33698, n33699, n33700,
         n33701, n33702, n33703, n33704, n33705, n33706, n33707, n33708,
         n33709, n33710, n33711, n33712, n33713, n33714, n33715, n33716,
         n33717, n33718, n33719, n33720, n33721, n33722, n33723, n33724,
         n33725, n33726, n33727, n33728, n33729, n33730, n33731, n33732,
         n33733, n33734, n33735, n33736, n33737, n33738, n33739, n33740,
         n33741, n33742, n33743, n33744, n33745, n33746, n33747, n33748,
         n33749, n33750, n33751, n33752, n33753, n33754, n33755, n33756,
         n33757, n33758, n33759, n33760, n33761, n33762, n33763, n33764,
         n33765, n33766, n33767, n33768, n33769, n33770, n33771, n33772,
         n33773, n33774, n33775, n33776, n33777, n33778, n33779, n33780,
         n33781, n33782, n33783, n33784, n33785, n33786, n33787, n33788,
         n33789, n33790, n33791, n33792, n33793, n33794, n33795, n33796,
         n33797, n33798, n33799, n33800, n33801, n33802, n33803, n33804,
         n33805, n33806, n33807, n33808, n33809, n33810, n33811, n33812,
         n33813, n33814, n33815, n33816, n33817, n33818, n33819, n33820,
         n33821, n33822, n33823, n33824, n33825, n33826, n33827, n33828,
         n33829, n33830, n33831, n33832, n33833, n33834, n33835, n33836,
         n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844,
         n33845, n33846, n33847, n33848, n33849, n33850, n33851, n33852,
         n33853, n33854, n33855, n33856, n33857, n33858, n33859, n33860,
         n33861, n33862, n33863, n33864, n33865, n33866, n33867, n33868,
         n33869, n33870, n33871, n33872, n33873, n33874, n33875, n33876,
         n33877, n33878, n33879, n33880, n33881, n33882, n33883, n33884,
         n33885, n33886, n33887, n33888, n33889, n33890, n33891, n33892,
         n33893, n33894, n33895, n33896, n33897, n33898, n33899, n33900,
         n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908,
         n33909, n33910, n33911, n33912, n33913, n33914, n33915, n33916,
         n33917, n33918, n33919, n33920, n33921, n33922, n33923, n33924,
         n33925, n33926, n33927, n33928, n33929, n33930, n33931, n33932,
         n33933, n33934, n33935, n33936, n33937, n33938, n33939, n33940,
         n33941, n33942, n33943, n33944, n33945, n33946, n33947, n33948,
         n33949, n33950, n33951, n33952, n33953, n33954, n33955, n33956,
         n33957, n33958, n33959, n33960, n33961, n33962, n33963, n33964,
         n33965, n33966, n33967, n33968, n33969, n33970, n33971, n33972,
         n33973, n33974, n33975, n33976, n33977, n33978, n33979, n33980,
         n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988,
         n33989, n33990, n33991, n33992, n33993, n33994, n33995, n33996,
         n33997, n33998, n33999, n34000, n34001, n34002, n34003, n34004,
         n34005, n34006, n34007, n34008, n34009, n34010, n34011, n34012,
         n34013, n34014, n34015, n34016, n34017, n34018, n34019, n34020,
         n34021, n34022, n34023, n34024, n34025, n34026, n34027, n34028,
         n34029, n34030, n34031, n34032, n34033, n34034, n34035, n34036,
         n34037, n34038, n34039, n34040, n34041, n34042, n34043, n34044,
         n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052,
         n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060,
         n34061, n34062, n34063, n34064, n34065, n34066, n34067, n34068,
         n34069, n34070, n34071, n34072, n34073, n34074, n34075, n34076,
         n34077, n34078, n34079, n34080, n34081, n34082, n34083, n34084,
         n34085, n34086, n34087, n34088, n34089, n34090, n34091, n34092,
         n34093, n34094, n34095, n34096, n34097, n34098, n34099, n34100,
         n34101, n34102, n34103, n34104, n34105, n34106, n34107, n34108,
         n34109, n34110, n34111, n34112, n34113, n34114, n34115, n34116,
         n34117, n34118, n34119, n34120, n34121, n34122, n34123, n34124,
         n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132,
         n34133, n34134, n34135, n34136, n34137, n34138, n34139, n34140,
         n34141, n34142, n34143, n34144, n34145, n34146, n34147, n34148,
         n34149, n34150, n34151, n34152, n34153, n34154, n34155, n34156,
         n34157, n34158, n34159, n34160, n34161, n34162, n34163, n34164,
         n34165, n34166, n34167, n34168, n34169, n34170, n34171, n34172,
         n34173, n34174, n34175, n34176, n34177, n34178, n34179, n34180,
         n34181, n34182, n34183, n34184, n34185, n34186, n34187, n34188,
         n34189, n34190, n34191, n34192, n34193, n34194, n34195, n34196,
         n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34204,
         n34205, n34206, n34207, n34208, n34209, n34210, n34211, n34212,
         n34213, n34214, n34215, n34216, n34217, n34218, n34219, n34220,
         n34221, n34222, n34223, n34224, n34225, n34226, n34227, n34228,
         n34229, n34230, n34231, n34232, n34233, n34234, n34235, n34236,
         n34237, n34238, n34239, n34240, n34241, n34242, n34243, n34244,
         n34245, n34246, n34247, n34248, n34249, n34250, n34251, n34252,
         n34253, n34254, n34255, n34256, n34257, n34258, n34259, n34260,
         n34261, n34262, n34263, n34264, n34265, n34266, n34267, n34268,
         n34269, n34270, n34271, n34272, n34273, n34274, n34275, n34276,
         n34277, n34278, n34279, n34280, n34281, n34282, n34283, n34284,
         n34285, n34286, n34287, n34288, n34289, n34290, n34291, n34292,
         n34293, n34294, n34295, n34296, n34297, n34298, n34299, n34300,
         n34301, n34302, n34303, n34304, n34305, n34306, n34307, n34308,
         n34309, n34310, n34311, n34312, n34313, n34314, n34315, n34316,
         n34317, n34318, n34319, n34320, n34321, n34322, n34323, n34324,
         n34325, n34326, n34327, n34328, n34329, n34330, n34331, n34332,
         n34333, n34334, n34335, n34336, n34337, n34338, n34339, n34340,
         n34341, n34342, n34343, n34344, n34345, n34346, n34347, n34348,
         n34349, n34350, n34351, n34352, n34353, n34354, n34355, n34356,
         n34357, n34358, n34359, n34360, n34361, n34362, n34363, n34364,
         n34365, n34366, n34367, n34368, n34369, n34370, n34371, n34372,
         n34373, n34374, n34375, n34376, n34377, n34378, n34379, n34380,
         n34381, n34382, n34383, n34384, n34385, n34386, n34387, n34388,
         n34389, n34390, n34391, n34392, n34393, n34394, n34395, n34396,
         n34397, n34398, n34399, n34400, n34401, n34402, n34403, n34404,
         n34405, n34406, n34407, n34408, n34409, n34410, n34411, n34412,
         n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420,
         n34421, n34422, n34423, n34424, n34425, n34426, n34427, n34428,
         n34429, n34430, n34431, n34432, n34433, n34434, n34435, n34436,
         n34437, n34438, n34439, n34440, n34441, n34442, n34443, n34444,
         n34445, n34446, n34447, n34448, n34449, n34450, n34451, n34452,
         n34453, n34454, n34455, n34456, n34457, n34458, n34459, n34460,
         n34461, n34462, n34463, n34464, n34465, n34466, n34467, n34468,
         n34469, n34470, n34471, n34472, n34473, n34474, n34475, n34476,
         n34477, n34478, n34479, n34480, n34481, n34482, n34483, n34484,
         n34485, n34486, n34487, n34488, n34489, n34490, n34491, n34492,
         n34493, n34494, n34495, n34496, n34497, n34498, n34499, n34500,
         n34501, n34502, n34503, n34504, n34505, n34506, n34507, n34508,
         n34509, n34510, n34511, n34512, n34513, n34514, n34515, n34516,
         n34517, n34518, n34519, n34520, n34521, n34522, n34523, n34524,
         n34525, n34526, n34527, n34528, n34529, n34530, n34531, n34532,
         n34533, n34534, n34535, n34536, n34537, n34538, n34539, n34540,
         n34541, n34542, n34543, n34544, n34545, n34546, n34547, n34548,
         n34549, n34550, n34551, n34552, n34553, n34554, n34555, n34556,
         n34557, n34558, n34559, n34560, n34561, n34562, n34563, n34564,
         n34565, n34566, n34567, n34568, n34569, n34570, n34571, n34572,
         n34573, n34574, n34575, n34576, n34577, n34578, n34579, n34580,
         n34581, n34582, n34583, n34584, n34585, n34586, n34587, n34588,
         n34589, n34590, n34591, n34592, n34593, n34594, n34595, n34596,
         n34597, n34598, n34599, n34600, n34601, n34602, n34603, n34604,
         n34605, n34606, n34607, n34608, n34609, n34610, n34611, n34612,
         n34613, n34614, n34615, n34616, n34617, n34618, n34619, n34620,
         n34621, n34622, n34623, n34624, n34625, n34626, n34627, n34628,
         n34629, n34630, n34631, n34632, n34633, n34634, n34635, n34636,
         n34637, n34638, n34639, n34640, n34641, n34642, n34643, n34644,
         n34645, n34646, n34647, n34648, n34649, n34650, n34651, n34652,
         n34653, n34654, n34655, n34656, n34657, n34658, n34659, n34660,
         n34661, n34662, n34663, n34664, n34665, n34666, n34667, n34668,
         n34669, n34670, n34671, n34672, n34673, n34674, n34675, n34676,
         n34677, n34678, n34679, n34680, n34681, n34682, n34683, n34684,
         n34685, n34686, n34687, n34688, n34689, n34690, n34691, n34692,
         n34693, n34694, n34695, n34696, n34697, n34698, n34699, n34700,
         n34701, n34702, n34703, n34704, n34705, n34706, n34707, n34708,
         n34709, n34710, n34711, n34712, n34713, n34714, n34715, n34716,
         n34717, n34718, n34719, n34720, n34721, n34722, n34723, n34724,
         n34725, n34726, n34727, n34728, n34729, n34730, n34731, n34732,
         n34733, n34734, n34735, n34736, n34737, n34738, n34739, n34740,
         n34741, n34742, n34743, n34744, n34745, n34746, n34747, n34748,
         n34749, n34750, n34751, n34752, n34753, n34754, n34755, n34756,
         n34757, n34758, n34759, n34760, n34761, n34762, n34763, n34764,
         n34765, n34766, n34767, n34768, n34769, n34770, n34771, n34772,
         n34773, n34774, n34775, n34776, n34777, n34778, n34779, n34780,
         n34781, n34782, n34783, n34784, n34785, n34786, n34787, n34788,
         n34789, n34790, n34791, n34792, n34793, n34794, n34795, n34796,
         n34797, n34798, n34799, n34800, n34801, n34802, n34803, n34804,
         n34805, n34806, n34807, n34808, n34809, n34810, n34811, n34812,
         n34813, n34814, n34815, n34816, n34817, n34818, n34819, n34820,
         n34821, n34822, n34823, n34824, n34825, n34826, n34827, n34828,
         n34829, n34830, n34831, n34832, n34833, n34834, n34835, n34836,
         n34837, n34838, n34839, n34840, n34841, n34842, n34843, n34844,
         n34845, n34846, n34847, n34848, n34849, n34850, n34851, n34852,
         n34853, n34854, n34855, n34856, n34857, n34858, n34859, n34860,
         n34861, n34862, n34863, n34864, n34865, n34866, n34867, n34868,
         n34869, n34870, n34871, n34872, n34873, n34874, n34875, n34876,
         n34877, n34878, n34879, n34880, n34881, n34882, n34883, n34884,
         n34885, n34886, n34887, n34888, n34889, n34890, n34891, n34892,
         n34893, n34894, n34895, n34896, n34897, n34898, n34899, n34900,
         n34901, n34902, n34903, n34904, n34905, n34906, n34907, n34908,
         n34909, n34910, n34911, n34912, n34913, n34914, n34915, n34916,
         n34917, n34918, n34919, n34920, n34921, n34922, n34923, n34924,
         n34925, n34926, n34927, n34928, n34929, n34930, n34931, n34932,
         n34933, n34934, n34935, n34936, n34937, n34938, n34939, n34940,
         n34941, n34942, n34943, n34944, n34945, n34946, n34947, n34948,
         n34949, n34950, n34951, n34952, n34953, n34954, n34955, n34956,
         n34957, n34958, n34959, n34960, n34961, n34962, n34963, n34964,
         n34965, n34966, n34967, n34968, n34969, n34970, n34971, n34972,
         n34973, n34974, n34975, n34976, n34977, n34978, n34979, n34980,
         n34981, n34982, n34983, n34984, n34985, n34986, n34987, n34988,
         n34989, n34990, n34991, n34992, n34993, n34994, n34995, n34996,
         n34997, n34998, n34999, n35000, n35001, n35002, n35003, n35004,
         n35005, n35006, n35007, n35008, n35009, n35010, n35011, n35012,
         n35013, n35014, n35015, n35016, n35017, n35018, n35019, n35020,
         n35021, n35022, n35023, n35024, n35025, n35026, n35027, n35028,
         n35029, n35030, n35031, n35032, n35033, n35034, n35035, n35036,
         n35037, n35038, n35039, n35040, n35041, n35042, n35043, n35044,
         n35045, n35046, n35047, n35048, n35049, n35050, n35051, n35052,
         n35053, n35054, n35055, n35056, n35057, n35058, n35059, n35060,
         n35061, n35062, n35063, n35064, n35065, n35066, n35067, n35068,
         n35069, n35070, n35071, n35072, n35073, n35074, n35075, n35076,
         n35077, n35078, n35079, n35080, n35081, n35082, n35083, n35084,
         n35085, n35086, n35087, n35088, n35089, n35090, n35091, n35092,
         n35093, n35094, n35095, n35096, n35097, n35098, n35099, n35100,
         n35101, n35102, n35103, n35104, n35105, n35106, n35107, n35108,
         n35109, n35110, n35111, n35112, n35113, n35114, n35115, n35116,
         n35117, n35118, n35119, n35120, n35121, n35122, n35123, n35124,
         n35125, n35126, n35127, n35128, n35129, n35130, n35131, n35132,
         n35133, n35134, n35135, n35136, n35137, n35138, n35139, n35140,
         n35141, n35142, n35143, n35144, n35145, n35146, n35147, n35148,
         n35149, n35150, n35151, n35152, n35153, n35154, n35155, n35156,
         n35157, n35158, n35159, n35160, n35161, n35162, n35163, n35164,
         n35165, n35166, n35167, n35168, n35169, n35170, n35171, n35172,
         n35173, n35174, n35175, n35176, n35177, n35178, n35179, n35180,
         n35181, n35182, n35183, n35184, n35185, n35186, n35187, n35188,
         n35189, n35190, n35191, n35192, n35193, n35194, n35195, n35196,
         n35197, n35198, n35199, n35200, n35201, n35202, n35203, n35204,
         n35205, n35206, n35207, n35208, n35209, n35210, n35211, n35212,
         n35213, n35214, n35215, n35216, n35217, n35218, n35219, n35220,
         n35221, n35222, n35223, n35224, n35225, n35226, n35227, n35228,
         n35229, n35230, n35231, n35232, n35233, n35234, n35235, n35236,
         n35237, n35238, n35239, n35240, n35241, n35242, n35243, n35244,
         n35245, n35246, n35247, n35248, n35249, n35250, n35251, n35252,
         n35253, n35254, n35255, n35256, n35257, n35258, n35259, n35260,
         n35261, n35262, n35263, n35264, n35265, n35266, n35267, n35268,
         n35269, n35270, n35271, n35272, n35273, n35274, n35275, n35276,
         n35277, n35278, n35279, n35280, n35281, n35282, n35283, n35284,
         n35285, n35286, n35287, n35288, n35289, n35290, n35291, n35292,
         n35293, n35294, n35295, n35296, n35297, n35298, n35299, n35300,
         n35301, n35302, n35303, n35304, n35305, n35306, n35307, n35308,
         n35309, n35310, n35311, n35312, n35313, n35314, n35315, n35316,
         n35317, n35318, n35319, n35320, n35321, n35322, n35323, n35324,
         n35325, n35326, n35327, n35328, n35329, n35330, n35331, n35332,
         n35333, n35334, n35335, n35336, n35337, n35338, n35339, n35340,
         n35341, n35342, n35343, n35344, n35345, n35346, n35347, n35348,
         n35349, n35350, n35351, n35352, n35353, n35354, n35355, n35356,
         n35357, n35358, n35359, n35360, n35361, n35362, n35363, n35364,
         n35365, n35366, n35367, n35368, n35369, n35370, n35371, n35372,
         n35373, n35374, n35375, n35376, n35377, n35378, n35379, n35380,
         n35381, n35382, n35383, n35384, n35385, n35386, n35387, n35388,
         n35389, n35390, n35391, n35392, n35393, n35394, n35395, n35396,
         n35397, n35398, n35399, n35400, n35401, n35402, n35403, n35404,
         n35405, n35406, n35407, n35408, n35409, n35410, n35411, n35412,
         n35413, n35414, n35415, n35416, n35417, n35418, n35419, n35420,
         n35421, n35422, n35423, n35424, n35425, n35426, n35427, n35428,
         n35429, n35430, n35431, n35432, n35433, n35434, n35435, n35436,
         n35437, n35438, n35439, n35440, n35441, n35442, n35443, n35444,
         n35445, n35446, n35447, n35448, n35449, n35450, n35451, n35452,
         n35453, n35454, n35455, n35456, n35457, n35458, n35459, n35460,
         n35461, n35462, n35463, n35464, n35465, n35466, n35467, n35468,
         n35469, n35470, n35471, n35472, n35473, n35474, n35475, n35476,
         n35477, n35478, n35479, n35480, n35481, n35482, n35483, n35484,
         n35485, n35486, n35487, n35488, n35489, n35490, n35491, n35492,
         n35493, n35494, n35495, n35496, n35497, n35498, n35499, n35500,
         n35501, n35502, n35503, n35504, n35505, n35506, n35507, n35508,
         n35509, n35510, n35511, n35512, n35513, n35514, n35515, n35516,
         n35517, n35518, n35519, n35520, n35521, n35522, n35523, n35524,
         n35525, n35526, n35527, n35528, n35529, n35530, n35531, n35532,
         n35533, n35534, n35535, n35536, n35537, n35538, n35539, n35540,
         n35541, n35542, n35543, n35544, n35545, n35546, n35547, n35548,
         n35549, n35550, n35551, n35552, n35553, n35554, n35555, n35556,
         n35557, n35558, n35559, n35560, n35561, n35562, n35563, n35564,
         n35565, n35566, n35567, n35568, n35569, n35570, n35571, n35572,
         n35573, n35574, n35575, n35576, n35577, n35578, n35579, n35580,
         n35581, n35582, n35583, n35584, n35585, n35586, n35587, n35588,
         n35589, n35590, n35591, n35592, n35593, n35594, n35595, n35596,
         n35597, n35598, n35599, n35600, n35601, n35602, n35603, n35604,
         n35605, n35606, n35607, n35608, n35609, n35610, n35611, n35612,
         n35613, n35614, n35615, n35616, n35617, n35618, n35619, n35620,
         n35621, n35622, n35623, n35624, n35625, n35626, n35627, n35628,
         n35629, n35630, n35631, n35632, n35633, n35634, n35635, n35636,
         n35637, n35638, n35639, n35640, n35641, n35642, n35643, n35644,
         n35645, n35646, n35647, n35648, n35649, n35650, n35651, n35652,
         n35653, n35654, n35655, n35656, n35657, n35658, n35659, n35660,
         n35661, n35662, n35663, n35664, n35665, n35666, n35667, n35668,
         n35669, n35670, n35671, n35672, n35673, n35674, n35675, n35676,
         n35677, n35678, n35679, n35680, n35681, n35682, n35683, n35684,
         n35685, n35686, n35687, n35688, n35689, n35690, n35691, n35692,
         n35693, n35694, n35695, n35696, n35697, n35698, n35699, n35700,
         n35701, n35702, n35703, n35704, n35705, n35706, n35707, n35708,
         n35709, n35710, n35711, n35712, n35713, n35714, n35715, n35716,
         n35717, n35718, n35719, n35720, n35721, n35722, n35723, n35724,
         n35725, n35726, n35727, n35728, n35729, n35730, n35731, n35732,
         n35733, n35734, n35735, n35736, n35737, n35738, n35739, n35740,
         n35741, n35742, n35743, n35744, n35745, n35746, n35747, n35748,
         n35749, n35750, n35751, n35752, n35753, n35754, n35755, n35756,
         n35757, n35758, n35759, n35760, n35761, n35762, n35763, n35764,
         n35765, n35766, n35767, n35768, n35769, n35770, n35771, n35772,
         n35773, n35774, n35775, n35776, n35777, n35778, n35779, n35780,
         n35781, n35782, n35783, n35784, n35785, n35786, n35787, n35788,
         n35789, n35790, n35791, n35792, n35793, n35794, n35795, n35796,
         n35797, n35798, n35799, n35800, n35801, n35802, n35803, n35804,
         n35805, n35806, n35807, n35808, n35809, n35810, n35811, n35812,
         n35813, n35814, n35815, n35816, n35817, n35818, n35819, n35820,
         n35821, n35822, n35823, n35824, n35825, n35826, n35827, n35828,
         n35829, n35830, n35831, n35832, n35833, n35834, n35835, n35836,
         n35837, n35838, n35839, n35840, n35841, n35842, n35843, n35844,
         n35845, n35846, n35847, n35848, n35849, n35850, n35851, n35852,
         n35853, n35854, n35855, n35856, n35857, n35858, n35859, n35860,
         n35861, n35862, n35863, n35864, n35865, n35866, n35867, n35868,
         n35869, n35870, n35871, n35872, n35873, n35874, n35875, n35876,
         n35877, n35878, n35879, n35880, n35881, n35882, n35883, n35884,
         n35885, n35886, n35887, n35888, n35889, n35890, n35891, n35892,
         n35893, n35894, n35895, n35896, n35897, n35898, n35899, n35900,
         n35901, n35902, n35903, n35904, n35905, n35906, n35907, n35908,
         n35909, n35910, n35911, n35912, n35913, n35914, n35915, n35916,
         n35917, n35918, n35919, n35920, n35921, n35922, n35923, n35924,
         n35925, n35926, n35927, n35928, n35929, n35930, n35931, n35932,
         n35933, n35934, n35935, n35936, n35937, n35938, n35939, n35940,
         n35941, n35942, n35943, n35944, n35945, n35946, n35947, n35948,
         n35949, n35950, n35951, n35952, n35953, n35954, n35955, n35956,
         n35957, n35958, n35959, n35960, n35961, n35962, n35963, n35964,
         n35965, n35966, n35967, n35968, n35969, n35970, n35971, n35972,
         n35973, n35974, n35975, n35976, n35977, n35978, n35979, n35980,
         n35981, n35982, n35983, n35984, n35985, n35986, n35987, n35988,
         n35989, n35990, n35991, n35992, n35993, n35994, n35995, n35996,
         n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004,
         n36005, n36006, n36007, n36008, n36009, n36010, n36011, n36012,
         n36013, n36014, n36015, n36016, n36017, n36018, n36019, n36020,
         n36021, n36022, n36023, n36024, n36025, n36026, n36027, n36028,
         n36029, n36030, n36031, n36032, n36033, n36034, n36035, n36036,
         n36037, n36038, n36039, n36040, n36041, n36042, n36043, n36044,
         n36045, n36046, n36047, n36048, n36049, n36050, n36051, n36052,
         n36053, n36054, n36055, n36056, n36057, n36058, n36059, n36060,
         n36061, n36062, n36063, n36064, n36065, n36066, n36067, n36068,
         n36069, n36070, n36071, n36072, n36073, n36074, n36075, n36076,
         n36077, n36078, n36079, n36080, n36081, n36082, n36083, n36084,
         n36085, n36086, n36087, n36088, n36089, n36090, n36091, n36092,
         n36093, n36094, n36095, n36096, n36097, n36098, n36099, n36100,
         n36101, n36102, n36103, n36104, n36105, n36106, n36107, n36108,
         n36109, n36110, n36111, n36112, n36113, n36114, n36115, n36116,
         n36117, n36118, n36119, n36120, n36121, n36122, n36123, n36124,
         n36125, n36126, n36127, n36128, n36129, n36130, n36131, n36132,
         n36133, n36134, n36135, n36136, n36137, n36138, n36139, n36140,
         n36141, n36142, n36143, n36144, n36145, n36146, n36147, n36148,
         n36149, n36150, n36151, n36152, n36153, n36154, n36155, n36156,
         n36157, n36158, n36159, n36160, n36161, n36162, n36163, n36164,
         n36165, n36166, n36167, n36168, n36169, n36170, n36171, n36172,
         n36173, n36174, n36175, n36176, n36177, n36178, n36179, n36180,
         n36181, n36182, n36183, n36184, n36185, n36186, n36187, n36188,
         n36189, n36190, n36191, n36192, n36193, n36194, n36195, n36196,
         n36197, n36198, n36199, n36200, n36201, n36202, n36203, n36204,
         n36205, n36206, n36207, n36208, n36209, n36210, n36211, n36212,
         n36213, n36214, n36215, n36216, n36217, n36218, n36219, n36220,
         n36221, n36222, n36223, n36224, n36225, n36226, n36227, n36228,
         n36229, n36230, n36231, n36232, n36233, n36234, n36235, n36236,
         n36237, n36238, n36239, n36240, n36241, n36242, n36243, n36244,
         n36245, n36246, n36247, n36248, n36249, n36250, n36251, n36252,
         n36253, n36254, n36255, n36256, n36257, n36258, n36259, n36260,
         n36261, n36262, n36263, n36264, n36265, n36266, n36267, n36268,
         n36269, n36270, n36271, n36272, n36273, n36274, n36275, n36276,
         n36277, n36278, n36279, n36280, n36281, n36282, n36283, n36284,
         n36285, n36286, n36287, n36288, n36289, n36290, n36291, n36292,
         n36293, n36294, n36295, n36296, n36297, n36298, n36299, n36300,
         n36301, n36302, n36303, n36304, n36305, n36306, n36307, n36308,
         n36309, n36310, n36311, n36312, n36313, n36314, n36315, n36316,
         n36317, n36318, n36319, n36320, n36321, n36322, n36323, n36324,
         n36325, n36326, n36327, n36328, n36329, n36330, n36331, n36332,
         n36333, n36334, n36335, n36336, n36337, n36338, n36339, n36340,
         n36341, n36342, n36343, n36344, n36345, n36346, n36347, n36348,
         n36349, n36350, n36351, n36352, n36353, n36354, n36355, n36356,
         n36357, n36358, n36359, n36360, n36361, n36362, n36363, n36364,
         n36365, n36366, n36367, n36368, n36369, n36370, n36371, n36372,
         n36373, n36374, n36375, n36376, n36377, n36378, n36379, n36380,
         n36381, n36382, n36383, n36384, n36385, n36386, n36387, n36388,
         n36389, n36390, n36391, n36392, n36393, n36394, n36395, n36396,
         n36397, n36398, n36399, n36400, n36401, n36402, n36403, n36404,
         n36405, n36406, n36407, n36408, n36409, n36410, n36411, n36412,
         n36413, n36414, n36415, n36416, n36417, n36418, n36419, n36420,
         n36421, n36422, n36423, n36424, n36425, n36426, n36427, n36428,
         n36429, n36430, n36431, n36432, n36433, n36434, n36435, n36436,
         n36437, n36438, n36439, n36440, n36441, n36442, n36443, n36444,
         n36445, n36446, n36447, n36448, n36449, n36450, n36451, n36452,
         n36453, n36454, n36455, n36456, n36457, n36458, n36459, n36460,
         n36461, n36462, n36463, n36464, n36465, n36466, n36467, n36468,
         n36469, n36470, n36471, n36472, n36473, n36474, n36475, n36476,
         n36477, n36478, n36479, n36480, n36481, n36482, n36483, n36484,
         n36485, n36486, n36487, n36488, n36489, n36490, n36491, n36492,
         n36493, n36494, n36495, n36496, n36497, n36498, n36499, n36500,
         n36501, n36502, n36503, n36504, n36505, n36506, n36507, n36508,
         n36509, n36510, n36511, n36512, n36513, n36514, n36515, n36516,
         n36517, n36518, n36519, n36520, n36521, n36522, n36523, n36524,
         n36525, n36526, n36527, n36528, n36529, n36530, n36531, n36532,
         n36533, n36534, n36535, n36536, n36537, n36538, n36539, n36540,
         n36541, n36542, n36543, n36544, n36545, n36546, n36547, n36548,
         n36549, n36550, n36551, n36552, n36553, n36554, n36555, n36556,
         n36557, n36558, n36559, n36560, n36561, n36562, n36563, n36564,
         n36565, n36566, n36567, n36568, n36569, n36570, n36571, n36572,
         n36573, n36574, n36575, n36576, n36577, n36578, n36579, n36580,
         n36581, n36582, n36583, n36584, n36585, n36586, n36587, n36588,
         n36589, n36590, n36591, n36592, n36593, n36594, n36595, n36596,
         n36597, n36598, n36599, n36600, n36601, n36602, n36603, n36604,
         n36605, n36606, n36607, n36608, n36609, n36610, n36611, n36612,
         n36613, n36614, n36615, n36616, n36617, n36618, n36619, n36620,
         n36621, n36622, n36623, n36624, n36625, n36626, n36627, n36628,
         n36629, n36630, n36631, n36632, n36633, n36634, n36635, n36636,
         n36637, n36638, n36639, n36640, n36641, n36642, n36643, n36644,
         n36645, n36646, n36647, n36648, n36649, n36650, n36651, n36652,
         n36653, n36654, n36655, n36656, n36657, n36658, n36659, n36660,
         n36661, n36662, n36663, n36664, n36665, n36666, n36667, n36668,
         n36669, n36670, n36671, n36672, n36673, n36674, n36675, n36676,
         n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684,
         n36685, n36686, n36687, n36688, n36689, n36690, n36691, n36692,
         n36693, n36694, n36695, n36696, n36697, n36698, n36699, n36700,
         n36701, n36702, n36703, n36704, n36705, n36706, n36707, n36708,
         n36709, n36710, n36711, n36712;
  wire   [10:2] u0_csr_r;
  wire   [7:0] u0_csr_r2;
  wire   [10:0] u0_csc_mask_r;
  wire   [6:2] u0_wb_addr_r;
  wire   [7:0] u0_csr_tj_val;
  wire   [7:0] u0_cs;
  wire   [7:1] u0_csc;
  wire   [27:0] u0_tms;
  wire   [7:0] u0_spec_req_cs;
  wire   [7:1] u0_sp_csc;
  wire   [27:0] u0_sp_tms;
  wire   [31:0] u0_csc0;
  wire   [31:0] u0_csc1;
  wire   [22:0] u1_u0_inc_in;
  wire   [3:0] u5_ack_cnt;
  wire   [3:0] u3_u0_rd_adr;
  wire   [7:0] u4_ps_cnt;
  wire   [7:0] u4_rfr_cnt;
  wire   [8:0] u5_timer2;
  wire   [7:0] u5_timer;
  wire   [1:0] u5_ir_cnt;
  wire   [10:0] u5_burst_cnt;
  wire   [65:0] u5_state;

  dffs1  \u5_burst_val_reg[10]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9017) );
  dffs1  \u1_page_size_reg[10]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n15531) );
  dffs1  \u5_burst_val_reg[9]  ( .DIN1(1'b0), .CLK(1'b0), .Q(n9018) );
  dffs1  \u1_page_size_reg[9]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n15530) );
  dffs1  \u5_burst_val_reg[8]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9019) );
  dffs1  \u1_page_size_reg[8]  ( .DIN1(1'b0), .CLK(1'b0), .Q(n15529) );
  dffs1  \u5_burst_val_reg[7]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9020) );
  dffs1  \u1_page_size_reg[7]  ( .DIN1(1'b0), .CLK(1'b0), 
                .Q(n15528) );
  dffs1  \u5_burst_val_reg[6]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9021) );
  dffs1  \u1_page_size_reg[6]  ( .DIN1(1'b0), .CLK(1'b0), 
                .Q(n15527) );
  dffs1  \u5_burst_val_reg[5]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9022) );
  dffs1  \u1_page_size_reg[5]  ( .DIN1(1'b0), .CLK(1'b0), 
                .Q(n15526) );
  dffs1  \u5_burst_val_reg[4]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9023) );
  dffs1  \u1_page_size_reg[4]  ( .DIN1(1'b0), .CLK(1'b0), 
                .Q(n15525) );
  dffs1  \u5_burst_val_reg[3]  ( .DIN1(1'b0), .CLK(1'b0), .Q(n9024) );
  dffs1  \u1_page_size_reg[3]  ( .DIN1(1'b0), .CLK(1'b0), 
                .QN(n4529) );
  dffs1  \u5_burst_val_reg[2]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9025) );
  dffs1  \u1_page_size_reg[2]  ( .DIN1(1'b0), .CLK(1'b0), 
                .Q(n5448) );
  dffs1  \u5_burst_val_reg[1]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9026) );
  dffs1  \u1_page_size_reg[1]  ( .DIN1(1'b0), .CLK(1'b0), 
                .Q(n5441) );
  dffs1  \u5_burst_val_reg[0]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9027) );
  dffs1  \u1_page_size_reg[0]  ( .DIN1(1'b0), .CLK(1'b0), 
                .Q(n5434) );
  dffs1  \u3_u0_dout_reg[31]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9028) );
  dffs1  \u3_u0_dout_reg[30]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9029) );
  dffs1  \u3_u0_dout_reg[29]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9030) );
  dffs1  \u3_u0_dout_reg[28]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9031) );
  dffs1  \u3_u0_dout_reg[27]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9032) );
  dffs1  \u3_u0_dout_reg[26]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9033) );
  dffs1  \u3_u0_dout_reg[25]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9034) );
  dffs1  \u3_u0_dout_reg[24]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9035) );
  dffs1  \u3_u0_dout_reg[23]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9036) );
  dffs1  \u3_u0_dout_reg[22]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9037) );
  dffs1  \u3_u0_dout_reg[21]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9038) );
  dffs1  \u3_u0_dout_reg[20]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9039) );
  dffs1  \u3_u0_dout_reg[19]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9040) );
  dffs1  \u3_u0_dout_reg[18]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9041) );
  dffs1  \u3_u0_dout_reg[17]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9042) );
  dffs1  \u3_u0_dout_reg[16]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9043) );
  dffs1  \u3_u0_dout_reg[15]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9044) );
  dffs1  \u3_u0_dout_reg[14]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9045) );
  dffs1  \u3_u0_dout_reg[13]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9046) );
  dffs1  \u3_u0_dout_reg[12]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9047) );
  dffs1  \u3_u0_dout_reg[11]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9048) );
  dffs1  \u3_u0_dout_reg[10]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9049) );
  dffs1  \u3_u0_dout_reg[9]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9050) );
  dffs1  \u3_u0_dout_reg[8]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9051) );
  dffs1  \u3_u0_dout_reg[7]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9052) );
  dffs1  \u3_u0_dout_reg[6]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9053) );
  dffs1  \u3_u0_dout_reg[5]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9054) );
  dffs1  \u3_u0_dout_reg[4]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9055) );
  dffs1  \u3_u0_dout_reg[3]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9056) );
  dffs1  \u3_u0_dout_reg[2]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9057) );
  dffs1  \u3_u0_dout_reg[1]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9058) );
  dffs1  \u3_u0_dout_reg[0]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9059) );
  dffs1  \u0_rf_dout_reg[4]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9060) );
  dffs1  \u0_rf_dout_reg[0]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9061) );
  dffs1  \u0_rf_dout_reg[5]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9062) );
  dffs1  \u0_rf_dout_reg[1]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9063) );
  dffs1  \u0_rf_dout_reg[2]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9064) );
  dffs1  \u0_rf_dout_reg[3]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9065) );
  dffs1  \u0_rf_dout_reg[6]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9066) );
  dffs1  \u0_rf_dout_reg[7]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9067) );
  dffs1  \u0_rf_dout_reg[8]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9068) );
  dffs1  \u0_rf_dout_reg[9]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9069) );
  dffs1  \u0_rf_dout_reg[10]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9070) );
  dffs1  \u0_rf_dout_reg[11]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9071) );
  dffs1  \u0_rf_dout_reg[12]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9072) );
  dffs1  \u0_rf_dout_reg[13]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9073) );
  dffs1  \u0_rf_dout_reg[14]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9074) );
  dffs1  \u0_rf_dout_reg[15]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9075) );
  dffs1  \u0_rf_dout_reg[16]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9076) );
  dffs1  \u0_rf_dout_reg[17]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9077) );
  dffs1  \u0_rf_dout_reg[18]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9078) );
  dffs1  \u0_rf_dout_reg[19]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9079) );
  dffs1  \u0_rf_dout_reg[20]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9080) );
  dffs1  \u0_rf_dout_reg[21]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9081) );
  dffs1  \u0_rf_dout_reg[22]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9082) );
  dffs1  \u0_rf_dout_reg[23]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9083) );
  dffs1  \u0_rf_dout_reg[24]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9084) );
  dffs1  \u0_rf_dout_reg[25]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9085) );
  dffs1  \u0_rf_dout_reg[26]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9086) );
  dffs1  \u0_rf_dout_reg[27]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9087) );
  dffs1  \u0_rf_dout_reg[28]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9088) );
  dffs1  \u0_rf_dout_reg[29]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9089) );
  dffs1  \u0_rf_dout_reg[30]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9090) );
  dffs1  \u0_rf_dout_reg[31]  ( .DIN1(1'b0), .CLK(1'b0),         .Q(n9091) );
  dffs1  u7_mc_adv__reg ( .DIN1(n9092), .CLK(mc_clk_i),         .Q(mc_adv_pad_o_) );
  dffs1  u7_mc_adsc__reg ( .DIN1(n19410), .CLK(mc_clk_i),         .Q(mc_adsc_pad_o_) );
  dffs1  u7_mc_cs_7_reg ( .DIN1(n9094), .CLK(mc_clk_i),         .Q(mc_cs_pad_o_[7]) );
  dffs1  u7_mc_cs_6_reg ( .DIN1(n9095), .CLK(mc_clk_i),         .Q(mc_cs_pad_o_[6]) );
  dffs1  u7_mc_cs_5_reg ( .DIN1(n9096), .CLK(mc_clk_i),         .Q(mc_cs_pad_o_[5]) );
  dffs1  u7_mc_cs_4_reg ( .DIN1(n9097), .CLK(mc_clk_i),         .Q(mc_cs_pad_o_[4]) );
  dffs1  u7_mc_cs_3_reg ( .DIN1(n9098), .CLK(mc_clk_i),         .Q(mc_cs_pad_o_[3]) );
  dffs1  u7_mc_cs_2_reg ( .DIN1(n9099), .CLK(mc_clk_i),         .Q(mc_cs_pad_o_[2]) );
  dffs1  u7_mc_cs_1_reg ( .DIN1(n9100), .CLK(mc_clk_i),         .Q(mc_cs_pad_o_[1]) );
  dffs1  u7_mc_cs_0_reg ( .DIN1(n9101), .CLK(mc_clk_i),         .Q(mc_cs_pad_o_[0]) );
  dffs1  u7_mc_ras__reg ( .DIN1(n9102), .CLK(mc_clk_i),         .Q(mc_ras_pad_o_) );
  dffs1  u7_mc_cas__reg ( .DIN1(\u5_temp_cs[1] ), .CLK(mc_clk_i), 
        .Q(mc_cas_pad_o_) );
  dffs1  u7_mc_we__reg ( .DIN1(n9103), .CLK(mc_clk_i),         .Q(mc_we_pad_o_) );
  dffs1  u7_mc_oe__reg ( .DIN1(n9104), .CLK(mc_clk_i),         .Q(mc_oe_pad_o_) );
  dffs1  \u7_mc_dqm_reg[0]  ( .DIN1(n9105), .CLK(mc_clk_i),         .Q(mc_dqm_pad_o[0]) );
  dffs1  \u7_mc_dqm_reg[1]  ( .DIN1(n9106), .CLK(mc_clk_i),         .Q(mc_dqm_pad_o[1]) );
  dffs1  \u7_mc_dqm_reg[2]  ( .DIN1(n9107), .CLK(mc_clk_i),         .Q(mc_dqm_pad_o[2]) );
  dffs1  \u7_mc_dqm_reg[3]  ( .DIN1(n9108), .CLK(mc_clk_i),         .Q(mc_dqm_pad_o[3]) );
  dffs1  \u7_mc_dqm_r2_reg[0]  ( .DIN1(n9109), .CLK(clk_i),         .QN(n4996) );
  dffs1  \u7_mc_dqm_r2_reg[1]  ( .DIN1(n9110), .CLK(clk_i),         .QN(n4995) );
  dffs1  \u7_mc_dqm_r2_reg[2]  ( .DIN1(n9111), .CLK(clk_i),         .QN(n4994) );
  dffs1  \u7_mc_dqm_r2_reg[3]  ( .DIN1(n9112), .CLK(clk_i),         .QN(n4993) );
  dffs1  \u7_mc_dqm_r_reg[0]  ( .DIN1(n9113), .CLK(clk_i),         .Q(n9109) );
  dffs1  \u7_mc_dqm_r_reg[1]  ( .DIN1(n9114), .CLK(clk_i),         .Q(n9110) );
  dffs1  \u7_mc_dqm_r_reg[2]  ( .DIN1(n9115), .CLK(clk_i),         .Q(n9111) );
  dffs1  \u7_mc_dqm_r_reg[3]  ( .DIN1(n9116), .CLK(clk_i),         .Q(n9112) );
  dffs1  \u7_mc_addr_reg[0]  ( .DIN1(n9117), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[0]) );
  dffs1  \u7_mc_addr_reg[1]  ( .DIN1(n9118), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[1]) );
  dffs1  \u7_mc_addr_reg[2]  ( .DIN1(n9119), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[2]) );
  dffs1  \u7_mc_addr_reg[3]  ( .DIN1(n9120), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[3]) );
  dffs1  \u7_mc_addr_reg[4]  ( .DIN1(n9121), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[4]) );
  dffs1  \u7_mc_addr_reg[5]  ( .DIN1(n9122), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[5]) );
  dffs1  \u7_mc_addr_reg[6]  ( .DIN1(n9123), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[6]) );
  dffs1  \u7_mc_addr_reg[7]  ( .DIN1(n9124), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[7]) );
  dffs1  \u7_mc_addr_reg[8]  ( .DIN1(n9125), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[8]) );
  dffs1  \u7_mc_addr_reg[9]  ( .DIN1(n9126), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[9]) );
  dffs1  \u7_mc_addr_reg[10]  ( .DIN1(n9127), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[10]) );
  dffs1  \u7_mc_addr_reg[11]  ( .DIN1(n9128), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[11]) );
  dffs1  \u7_mc_addr_reg[12]  ( .DIN1(n9129), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[12]) );
  dffs1  \u7_mc_addr_reg[13]  ( .DIN1(n9130), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[13]) );
  dffs1  \u7_mc_addr_reg[14]  ( .DIN1(n9131), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[14]) );
  dffs1  \u7_mc_addr_reg[15]  ( .DIN1(n9132), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[15]) );
  dffs1  \u7_mc_addr_reg[16]  ( .DIN1(n9133), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[16]) );
  dffs1  \u7_mc_addr_reg[17]  ( .DIN1(n9134), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[17]) );
  dffs1  \u7_mc_addr_reg[18]  ( .DIN1(n9135), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[18]) );
  dffs1  \u7_mc_addr_reg[19]  ( .DIN1(n9136), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[19]) );
  dffs1  \u7_mc_addr_reg[20]  ( .DIN1(n9137), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[20]) );
  dffs1  \u7_mc_addr_reg[21]  ( .DIN1(n9138), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[21]) );
  dffs1  \u7_mc_addr_reg[22]  ( .DIN1(n9139), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[22]) );
  dffs1  \u7_mc_addr_reg[23]  ( .DIN1(n9140), .CLK(mc_clk_i),         .Q(mc_addr_pad_o[23]) );
  dffs1  \u7_mc_dp_o_reg[0]  ( .DIN1(n9141), .CLK(mc_clk_i),         .Q(mc_dp_pad_o[0]) );
  dffs1  \u7_mc_dp_o_reg[1]  ( .DIN1(n9142), .CLK(mc_clk_i),         .Q(mc_dp_pad_o[1]) );
  dffs1  \u7_mc_dp_o_reg[2]  ( .DIN1(n9143), .CLK(mc_clk_i),         .Q(mc_dp_pad_o[2]) );
  dffs1  \u7_mc_dp_o_reg[3]  ( .DIN1(n9144), .CLK(mc_clk_i),         .Q(mc_dp_pad_o[3]) );
  dffs1  \u7_mc_data_o_reg[0]  ( .DIN1(n9145), .CLK(mc_clk_i), .Q(
        mc_data_pad_o[0]) );
  dffs1  \u7_mc_data_o_reg[1]  ( .DIN1(n9146), .CLK(mc_clk_i), .Q(
        mc_data_pad_o[1]) );
  dffs1  \u7_mc_data_o_reg[2]  ( .DIN1(n9147), .CLK(mc_clk_i), .Q(
        mc_data_pad_o[2]) );
  dffs1  \u7_mc_data_o_reg[3]  ( .DIN1(n9148), .CLK(mc_clk_i), .Q(
        mc_data_pad_o[3]) );
  dffs1  \u7_mc_data_o_reg[4]  ( .DIN1(n9149), .CLK(mc_clk_i), .Q(
        mc_data_pad_o[4]) );
  dffs1  \u7_mc_data_o_reg[5]  ( .DIN1(n9150), .CLK(mc_clk_i), .Q(
        mc_data_pad_o[5]) );
  dffs1  \u7_mc_data_o_reg[6]  ( .DIN1(n9151), .CLK(mc_clk_i), .Q(
        mc_data_pad_o[6]) );
  dffs1  \u7_mc_data_o_reg[7]  ( .DIN1(n9152), .CLK(mc_clk_i), .Q(
        mc_data_pad_o[7]) );
  dffs1  \u7_mc_data_o_reg[8]  ( .DIN1(n9153), .CLK(mc_clk_i), .Q(
        mc_data_pad_o[8]) );
  dffs1  \u7_mc_data_o_reg[9]  ( .DIN1(n9154), .CLK(mc_clk_i), .Q(
        mc_data_pad_o[9]) );
  dffs1  \u7_mc_data_o_reg[10]  ( .DIN1(n9155), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[10]) );
  dffs1  \u7_mc_data_o_reg[11]  ( .DIN1(n9156), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[11]) );
  dffs1  \u7_mc_data_o_reg[12]  ( .DIN1(n9157), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[12]) );
  dffs1  \u7_mc_data_o_reg[13]  ( .DIN1(n9158), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[13]) );
  dffs1  \u7_mc_data_o_reg[14]  ( .DIN1(n9159), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[14]) );
  dffs1  \u7_mc_data_o_reg[15]  ( .DIN1(n9160), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[15]) );
  dffs1  \u7_mc_data_o_reg[16]  ( .DIN1(n9161), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[16]) );
  dffs1  \u7_mc_data_o_reg[17]  ( .DIN1(n9162), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[17]) );
  dffs1  \u7_mc_data_o_reg[18]  ( .DIN1(n9163), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[18]) );
  dffs1  \u7_mc_data_o_reg[19]  ( .DIN1(n9164), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[19]) );
  dffs1  \u7_mc_data_o_reg[20]  ( .DIN1(n9165), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[20]) );
  dffs1  \u7_mc_data_o_reg[21]  ( .DIN1(n9166), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[21]) );
  dffs1  \u7_mc_data_o_reg[22]  ( .DIN1(n9167), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[22]) );
  dffs1  \u7_mc_data_o_reg[23]  ( .DIN1(n9168), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[23]) );
  dffs1  \u7_mc_data_o_reg[24]  ( .DIN1(n9169), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[24]) );
  dffs1  \u7_mc_data_o_reg[25]  ( .DIN1(n9170), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[25]) );
  dffs1  \u7_mc_data_o_reg[26]  ( .DIN1(n9171), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[26]) );
  dffs1  \u7_mc_data_o_reg[27]  ( .DIN1(n9172), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[27]) );
  dffs1  \u7_mc_data_o_reg[28]  ( .DIN1(n9173), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[28]) );
  dffs1  \u7_mc_data_o_reg[29]  ( .DIN1(n9174), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[29]) );
  dffs1  \u7_mc_data_o_reg[30]  ( .DIN1(n9175), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[30]) );
  dffs1  \u7_mc_data_o_reg[31]  ( .DIN1(n9176), .CLK(mc_clk_i), 
        .Q(mc_data_pad_o[31]) );
  dffs1  u7_mc_data_oe_reg ( .DIN1(n9177), .CLK(mc_clk_i),         .Q(mc_doe_pad_doe_o) );
  dffs1  u7_mc_bg_reg ( .DIN1(n9178), .CLK(mc_clk_i),         .Q(mc_bg_pad_o) );
  dffs1  \u5_cmd_del_reg[1]  ( .DIN1(n9179), .CLK(clk_i),         .Q(n4531) );
  dffs1  \u5_cmd_r_reg[1]  ( .DIN1(n9180), .CLK(clk_i),         .Q(n9179) );
  dffs1  \u5_cmd_del_reg[0]  ( .DIN1(n9181), .CLK(clk_i),         .Q(n4532) );
  dffs1  \u5_cmd_r_reg[0]  ( .DIN1(n9182), .CLK(clk_i),         .Q(n9181) );
  dffs1  \u5_cmd_del_reg[2]  ( .DIN1(n9183), .CLK(clk_i),         .Q(n4530) );
  dffs1  \u5_cmd_r_reg[2]  ( .DIN1(n9184), .CLK(clk_i),         .Q(n9183) );
  dffs1  u5_cmd_a10_r_reg ( .DIN1(n9185), .CLK(clk_i),         .Q(n4535) );
  dffs1  \u5_timer_reg[6]  ( .DIN1(n9186), .CLK(clk_i),         .Q(u5_timer[6]) );
  dffs1  \u5_timer_reg[5]  ( .DIN1(n9187), .CLK(clk_i),         .Q(u5_timer[5]) );
  dffs1  \u5_timer_reg[4]  ( .DIN1(n9188), .CLK(clk_i),         .Q(u5_timer[4]) );
  dffs1  \u5_timer_reg[3]  ( .DIN1(n9189), .CLK(clk_i),         .Q(u5_timer[3]) );
  dffs1  \u5_timer_reg[2]  ( .DIN1(n9190), .CLK(clk_i),         .Q(u5_timer[2]) );
  dffs1  \u5_timer_reg[0]  ( .DIN1(n9191), .CLK(clk_i),         .Q(u5_timer[0]) );
  dffs1  \u5_timer_reg[7]  ( .DIN1(n9192), .CLK(clk_i),         .Q(u5_timer[7]) );
  dffs1  u5_cke_r_reg ( .DIN1(n9193), .CLK(clk_i),         .Q(u5_cke_r) );
  dffs1  u5_cnt_reg ( .DIN1(n9194), .CLK(clk_i), .Q(u5_cnt)
         );
  dffs1  u5_data_oe_reg ( .DIN1(n9195), .CLK(clk_i),         .QN(n15501) );
  dffs1  u5_data_oe_r2_reg ( .DIN1(n9196), .CLK(clk_i),         .Q(n4536) );
  dffs1  u5_data_oe_r_reg ( .DIN1(n9197), .CLK(clk_i),         .Q(n9196) );
  dffs1  \u3_mc_data_o_reg[0]  ( .DIN1(n9198), .CLK(clk_i),         .Q(n9145) );
  dffs1  \u3_mc_data_o_reg[1]  ( .DIN1(n9199), .CLK(clk_i),         .Q(n9146) );
  dffs1  \u3_mc_data_o_reg[2]  ( .DIN1(n9200), .CLK(clk_i),         .Q(n9147) );
  dffs1  \u3_mc_data_o_reg[3]  ( .DIN1(n9201), .CLK(clk_i),         .Q(n9148) );
  dffs1  \u3_mc_data_o_reg[4]  ( .DIN1(n9202), .CLK(clk_i),         .Q(n9149) );
  dffs1  \u3_mc_data_o_reg[5]  ( .DIN1(n9203), .CLK(clk_i),         .Q(n9150) );
  dffs1  \u3_mc_data_o_reg[6]  ( .DIN1(n9204), .CLK(clk_i),         .Q(n9151) );
  dffs1  \u3_mc_data_o_reg[7]  ( .DIN1(n9205), .CLK(clk_i),         .Q(n9152) );
  dffs1  \u3_mc_data_o_reg[8]  ( .DIN1(n9206), .CLK(clk_i),         .Q(n9153) );
  dffs1  \u3_mc_data_o_reg[9]  ( .DIN1(n9207), .CLK(clk_i),         .Q(n9154) );
  dffs1  \u3_mc_data_o_reg[10]  ( .DIN1(n9208), .CLK(clk_i),         .Q(n9155) );
  dffs1  \u3_mc_data_o_reg[11]  ( .DIN1(n9209), .CLK(clk_i),         .Q(n9156) );
  dffs1  \u3_mc_data_o_reg[12]  ( .DIN1(n9210), .CLK(clk_i),         .Q(n9157) );
  dffs1  \u3_mc_data_o_reg[13]  ( .DIN1(n9211), .CLK(clk_i),         .Q(n9158) );
  dffs1  \u3_mc_data_o_reg[14]  ( .DIN1(n9212), .CLK(clk_i),         .Q(n9159) );
  dffs1  \u3_mc_data_o_reg[15]  ( .DIN1(n9213), .CLK(clk_i),         .Q(n9160) );
  dffs1  \u3_mc_data_o_reg[16]  ( .DIN1(n9214), .CLK(clk_i),         .Q(n9161) );
  dffs1  \u3_mc_data_o_reg[17]  ( .DIN1(n9215), .CLK(clk_i),         .Q(n9162) );
  dffs1  \u3_mc_data_o_reg[18]  ( .DIN1(n9216), .CLK(clk_i),         .Q(n9163) );
  dffs1  \u3_mc_data_o_reg[19]  ( .DIN1(n9217), .CLK(clk_i),         .Q(n9164) );
  dffs1  \u3_mc_data_o_reg[20]  ( .DIN1(n9218), .CLK(clk_i),         .Q(n9165) );
  dffs1  \u3_mc_data_o_reg[21]  ( .DIN1(n9219), .CLK(clk_i),         .Q(n9166) );
  dffs1  \u3_mc_data_o_reg[22]  ( .DIN1(n9220), .CLK(clk_i),         .Q(n9167) );
  dffs1  \u3_mc_data_o_reg[23]  ( .DIN1(n9221), .CLK(clk_i),         .Q(n9168) );
  dffs1  \u3_mc_data_o_reg[24]  ( .DIN1(n9222), .CLK(clk_i),         .Q(n9169) );
  dffs1  \u3_mc_data_o_reg[25]  ( .DIN1(n9223), .CLK(clk_i),         .Q(n9170) );
  dffs1  \u3_mc_data_o_reg[26]  ( .DIN1(n9224), .CLK(clk_i),         .Q(n9171) );
  dffs1  \u3_mc_data_o_reg[27]  ( .DIN1(n9225), .CLK(clk_i),         .Q(n9172) );
  dffs1  \u3_mc_data_o_reg[28]  ( .DIN1(n9226), .CLK(clk_i),         .Q(n9173) );
  dffs1  \u3_mc_data_o_reg[29]  ( .DIN1(n9227), .CLK(clk_i),         .Q(n9174) );
  dffs1  \u3_mc_data_o_reg[30]  ( .DIN1(n9228), .CLK(clk_i),         .Q(n9175) );
  dffs1  \u3_mc_data_o_reg[31]  ( .DIN1(n9229), .CLK(clk_i),         .Q(n9176) );
  dffs1  \u3_mc_dp_o_reg[3]  ( .DIN1(n9230), .CLK(clk_i),         .Q(n9144) );
  dffs1  \u3_mc_dp_o_reg[2]  ( .DIN1(n9231), .CLK(clk_i),         .Q(n9143) );
  dffs1  \u3_mc_dp_o_reg[1]  ( .DIN1(n9232), .CLK(clk_i),         .Q(n9142) );
  dffs1  \u3_mc_dp_o_reg[0]  ( .DIN1(n9233), .CLK(clk_i),         .Q(n9141) );
  dffs1  \u5_timer2_reg[6]  ( .DIN1(n9234), .CLK(clk_i),         .Q(u5_timer2[6]) );
  dffs1  \u5_timer2_reg[5]  ( .DIN1(n9235), .CLK(clk_i),         .Q(u5_timer2[5]) );
  dffs1  \u5_timer2_reg[4]  ( .DIN1(n9236), .CLK(clk_i),         .Q(u5_timer2[4]) );
  dffs1  \u5_timer2_reg[3]  ( .DIN1(n9237), .CLK(clk_i),         .Q(u5_timer2[3]) );
  dffs1  \u5_timer2_reg[2]  ( .DIN1(n9238), .CLK(clk_i),         .Q(u5_timer2[2]) );
  dffs1  \u5_timer2_reg[1]  ( .DIN1(n9239), .CLK(clk_i),         .Q(u5_timer2[1]) );
  dffs1  \u5_timer2_reg[0]  ( .DIN1(n9240), .CLK(clk_i),         .Q(u5_timer2[0]) );
  dffs1  \u5_timer2_reg[7]  ( .DIN1(n9241), .CLK(clk_i),         .Q(u5_timer2[7]) );
  dffs1  \u1_col_adr_reg[9]  ( .DIN1(n9242), .CLK(clk_i),         .QN(n36685) );
  dffs1  \u1_col_adr_reg[8]  ( .DIN1(n9243), .CLK(clk_i),         .QN(n36688) );
  dffs1  \u1_col_adr_reg[7]  ( .DIN1(n9244), .CLK(clk_i),         .QN(n36691) );
  dffs1  \u1_col_adr_reg[6]  ( .DIN1(n9245), .CLK(clk_i),         .QN(n36694) );
  dffs1  \u1_col_adr_reg[5]  ( .DIN1(n9246), .CLK(clk_i),         .QN(n36697) );
  dffs1  \u1_col_adr_reg[4]  ( .DIN1(n9247), .CLK(clk_i),         .QN(n36700) );
  dffs1  \u1_col_adr_reg[3]  ( .DIN1(n9248), .CLK(clk_i),         .QN(n36703) );
  dffs1  \u1_col_adr_reg[2]  ( .DIN1(n9249), .CLK(clk_i),         .QN(n36706) );
  dffs1  \u1_col_adr_reg[1]  ( .DIN1(n9250), .CLK(clk_i),         .QN(n36709) );
  dffs1  \u1_col_adr_reg[0]  ( .DIN1(n9251), .CLK(clk_i),         .QN(n36712) );
  dffs1  u5_wr_cycle_reg ( .DIN1(n9252), .CLK(clk_i),         .QN(n15502) );
  dffs1  \u0_spec_req_cs_reg[7]  ( .DIN1(n9253), .CLK(clk_i),         .QN(n15489) );
  dffs1  \u0_spec_req_cs_reg[6]  ( .DIN1(n9254), .CLK(clk_i),         .QN(n15490) );
  dffs1  \u0_spec_req_cs_reg[5]  ( .DIN1(n9255), .CLK(clk_i),         .QN(n15491) );
  dffs1  \u0_spec_req_cs_reg[4]  ( .DIN1(n9256), .CLK(clk_i),         .QN(n15492) );
  dffs1  \u0_spec_req_cs_reg[3]  ( .DIN1(n9257), .CLK(clk_i),         .QN(n15493) );
  dffs1  \u0_spec_req_cs_reg[2]  ( .DIN1(n9258), .CLK(clk_i),         .QN(n15494) );
  dffs1  \u0_sp_csc_reg[1]  ( .DIN1(n9259), .CLK(clk_i),         .Q(u0_sp_csc[1]) );
  dffs1  \u0_sp_csc_reg[2]  ( .DIN1(n9260), .CLK(clk_i),         .Q(u0_sp_csc[2]) );
  dffs1  \u0_sp_csc_reg[3]  ( .DIN1(n9261), .CLK(clk_i),         .Q(u0_sp_csc[3]) );
  dffs1  \u1_row_adr_reg[0]  ( .DIN1(n9262), .CLK(clk_i),         .QN(n36711) );
  dffs1  \u1_row_adr_reg[1]  ( .DIN1(n9263), .CLK(clk_i),         .QN(n36708) );
  dffs1  \u1_row_adr_reg[2]  ( .DIN1(n9264), .CLK(clk_i),         .QN(n36705) );
  dffs1  \u1_row_adr_reg[3]  ( .DIN1(n9265), .CLK(clk_i),         .QN(n36702) );
  dffs1  \u1_row_adr_reg[4]  ( .DIN1(n9266), .CLK(clk_i),         .QN(n36699) );
  dffs1  \u1_row_adr_reg[5]  ( .DIN1(n9267), .CLK(clk_i),         .QN(n36696) );
  dffs1  \u1_row_adr_reg[6]  ( .DIN1(n9268), .CLK(clk_i),         .QN(n36693) );
  dffs1  \u1_row_adr_reg[7]  ( .DIN1(n9269), .CLK(clk_i),         .QN(n36690) );
  dffs1  \u1_row_adr_reg[8]  ( .DIN1(n9270), .CLK(clk_i),         .QN(n36687) );
  dffs1  \u1_row_adr_reg[9]  ( .DIN1(n9271), .CLK(clk_i),         .QN(n36684) );
  dffs1  \u1_row_adr_reg[10]  ( .DIN1(n9272), .CLK(clk_i),         .QN(n36682) );
  dffs1  \u1_row_adr_reg[11]  ( .DIN1(n9273), .CLK(clk_i),         .QN(n36680) );
  dffs1  \u1_row_adr_reg[12]  ( .DIN1(n9274), .CLK(clk_i),         .QN(n36678) );
  dffs1  \u1_bank_adr_reg[1]  ( .DIN1(n9275), .CLK(clk_i),         .QN(n36673) );
  dffs1  \u1_bank_adr_reg[0]  ( .DIN1(n9276), .CLK(clk_i),         .QN(n36675) );
  dffs1  \u5_burst_cnt_reg[8]  ( .DIN1(n9277), .CLK(clk_i),         .Q(u5_burst_cnt[8]) );
  dffs1  \u5_burst_cnt_reg[7]  ( .DIN1(n9278), .CLK(clk_i),         .Q(u5_burst_cnt[7]) );
  dffs1  \u5_burst_cnt_reg[6]  ( .DIN1(n9279), .CLK(clk_i),         .Q(u5_burst_cnt[6]) );
  dffs1  \u5_burst_cnt_reg[5]  ( .DIN1(n9280), .CLK(clk_i),         .Q(u5_burst_cnt[5]) );
  dffs1  \u5_burst_cnt_reg[4]  ( .DIN1(n9281), .CLK(clk_i),         .Q(u5_burst_cnt[4]) );
  dffs1  \u5_burst_cnt_reg[3]  ( .DIN1(n9282), .CLK(clk_i),         .Q(u5_burst_cnt[3]) );
  dffs1  \u5_burst_cnt_reg[2]  ( .DIN1(n9283), .CLK(clk_i),         .Q(u5_burst_cnt[2]) );
  dffs1  \u5_burst_cnt_reg[1]  ( .DIN1(n9284), .CLK(clk_i),         .Q(u5_burst_cnt[1]) );
  dffs1  \u5_burst_cnt_reg[0]  ( .DIN1(n9285), .CLK(clk_i),         .Q(u5_burst_cnt[0]) );
  dffs1  \u5_burst_cnt_reg[9]  ( .DIN1(n9286), .CLK(clk_i),         .Q(u5_burst_cnt[9]) );
  dffs1  \u1_acs_addr_reg[23]  ( .DIN1(n9287), .CLK(clk_i),         .QN(n36664) );
  dffs1  \u1_acs_addr_reg[21]  ( .DIN1(n9288), .CLK(clk_i),         .Q(u1_u0_inc_in[21]) );
  dffs1  \u1_acs_addr_reg[20]  ( .DIN1(n9289), .CLK(clk_i),         .Q(u1_u0_inc_in[20]) );
  dffs1  \u1_acs_addr_reg[19]  ( .DIN1(n9290), .CLK(clk_i),         .Q(u1_u0_inc_in[19]) );
  dffs1  \u1_acs_addr_reg[18]  ( .DIN1(n9291), .CLK(clk_i),         .Q(u1_u0_inc_in[18]) );
  dffs1  \u1_acs_addr_reg[17]  ( .DIN1(n9292), .CLK(clk_i),         .Q(u1_u0_inc_in[17]) );
  dffs1  \u1_acs_addr_reg[16]  ( .DIN1(n9293), .CLK(clk_i),         .Q(u1_u0_inc_in[16]) );
  dffs1  \u1_acs_addr_reg[15]  ( .DIN1(n9294), .CLK(clk_i),         .Q(u1_u0_inc_in[15]) );
  dffs1  \u1_acs_addr_reg[14]  ( .DIN1(n9295), .CLK(clk_i),         .Q(u1_u0_inc_in[14]) );
  dffs1  \u1_acs_addr_reg[13]  ( .DIN1(n9296), .CLK(clk_i),         .Q(u1_u0_inc_in[13]) );
  dffs1  \u1_acs_addr_reg[22]  ( .DIN1(n9297), .CLK(clk_i),         .Q(u1_u0_inc_in[22]) );
  dffs1  \u1_acs_addr_reg[12]  ( .DIN1(n9298), .CLK(clk_i),         .Q(u1_u0_inc_in[12]) );
  dffs1  \u1_u0_out_r_reg[12]  ( .DIN1(N884), .CLK(clk_i),         .Q(\u1_u0_out_r[12] ) );
  dffs1  \u1_u0_out_r_reg[11]  ( .DIN1(N883), .CLK(clk_i),         .Q(n4581) );
  dffs1  \u1_acs_addr_reg[10]  ( .DIN1(n9299), .CLK(clk_i),         .Q(u1_u0_inc_in[10]) );
  dffs1  \u1_u0_out_r_reg[10]  ( .DIN1(N882), .CLK(clk_i),         .Q(n4570) );
  dffs1  \u1_acs_addr_reg[9]  ( .DIN1(n9300), .CLK(clk_i),         .Q(u1_u0_inc_in[9]) );
  dffs1  \u1_u0_out_r_reg[9]  ( .DIN1(N881), .CLK(clk_i),         .Q(n4571) );
  dffs1  \u1_acs_addr_reg[8]  ( .DIN1(n9301), .CLK(clk_i),         .Q(u1_u0_inc_in[8]) );
  dffs1  \u1_u0_out_r_reg[8]  ( .DIN1(N880), .CLK(clk_i),         .Q(n4572) );
  dffs1  \u1_acs_addr_reg[7]  ( .DIN1(n9302), .CLK(clk_i),         .Q(u1_u0_inc_in[7]) );
  dffs1  \u1_u0_out_r_reg[7]  ( .DIN1(N879), .CLK(clk_i),         .Q(n4573) );
  dffs1  \u1_acs_addr_reg[6]  ( .DIN1(n9303), .CLK(clk_i),         .Q(u1_u0_inc_in[6]) );
  dffs1  \u1_u0_out_r_reg[6]  ( .DIN1(N878), .CLK(clk_i),         .Q(n4574) );
  dffs1  \u1_acs_addr_reg[5]  ( .DIN1(n9304), .CLK(clk_i),         .Q(u1_u0_inc_in[5]) );
  dffs1  \u1_u0_out_r_reg[5]  ( .DIN1(N877), .CLK(clk_i),         .Q(n4575) );
  dffs1  \u1_acs_addr_reg[4]  ( .DIN1(n9305), .CLK(clk_i),         .Q(u1_u0_inc_in[4]) );
  dffs1  \u1_u0_out_r_reg[4]  ( .DIN1(N876), .CLK(clk_i),         .Q(n4576) );
  dffs1  \u1_acs_addr_reg[3]  ( .DIN1(n9306), .CLK(clk_i),         .Q(u1_u0_inc_in[3]) );
  dffs1  \u1_u0_out_r_reg[3]  ( .DIN1(N875), .CLK(clk_i),         .Q(n4577) );
  dffs1  \u1_acs_addr_reg[2]  ( .DIN1(n9307), .CLK(clk_i),         .Q(u1_u0_inc_in[2]) );
  dffs1  \u1_u0_out_r_reg[2]  ( .DIN1(N874), .CLK(clk_i),         .Q(n4578) );
  dffs1  \u1_acs_addr_reg[1]  ( .DIN1(n9308), .CLK(clk_i),         .Q(u1_u0_inc_in[1]) );
  dffs1  \u1_u0_out_r_reg[1]  ( .DIN1(N873), .CLK(clk_i),         .Q(n4579) );
  dffs1  \u1_acs_addr_reg[0]  ( .DIN1(n9309), .CLK(clk_i),         .Q(u1_u0_inc_in[0]) );
  dffs1  \u1_u0_out_r_reg[0]  ( .DIN1(N872), .CLK(clk_i),         .Q(n4580) );
  dffs1  \u1_acs_addr_reg[11]  ( .DIN1(n9310), .CLK(clk_i),         .Q(u1_u0_inc_in[11]) );
  dffs1  u5_oe__reg ( .DIN1(n19409), .CLK(clk_i), .Q(n4533)
         );
  dffs1  \u6_wb_data_o_reg[15]  ( .DIN1(n9312), .CLK(clk_i),         .Q(wb_data_o[15]) );
  dffs1  \u3_byte1_reg[7]  ( .DIN1(n9313), .CLK(clk_i),         .QN(n36659) );
  dffs1  \u6_wb_data_o_reg[14]  ( .DIN1(n9314), .CLK(clk_i),         .Q(wb_data_o[14]) );
  dffs1  \u3_byte1_reg[6]  ( .DIN1(n9315), .CLK(clk_i),         .QN(n36656) );
  dffs1  \u6_wb_data_o_reg[13]  ( .DIN1(n9316), .CLK(clk_i),         .Q(wb_data_o[13]) );
  dffs1  \u3_byte1_reg[5]  ( .DIN1(n9317), .CLK(clk_i),         .QN(n36653) );
  dffs1  \u6_wb_data_o_reg[12]  ( .DIN1(n9318), .CLK(clk_i),         .Q(wb_data_o[12]) );
  dffs1  \u3_byte1_reg[4]  ( .DIN1(n9319), .CLK(clk_i),         .QN(n36650) );
  dffs1  \u6_wb_data_o_reg[11]  ( .DIN1(n9320), .CLK(clk_i),         .Q(wb_data_o[11]) );
  dffs1  \u3_byte1_reg[3]  ( .DIN1(n9321), .CLK(clk_i),         .QN(n36647) );
  dffs1  \u6_wb_data_o_reg[10]  ( .DIN1(n9322), .CLK(clk_i),         .Q(wb_data_o[10]) );
  dffs1  \u3_byte1_reg[2]  ( .DIN1(n9323), .CLK(clk_i),         .QN(n36644) );
  dffs1  \u6_wb_data_o_reg[9]  ( .DIN1(n9324), .CLK(clk_i),         .Q(wb_data_o[9]) );
  dffs1  \u3_byte1_reg[1]  ( .DIN1(n9325), .CLK(clk_i),         .QN(n36641) );
  dffs1  \u6_wb_data_o_reg[8]  ( .DIN1(n9326), .CLK(clk_i),         .Q(wb_data_o[8]) );
  dffs1  \u3_byte1_reg[0]  ( .DIN1(n9327), .CLK(clk_i),         .QN(n36638) );
  dffs1  u5_pack_le1_reg ( .DIN1(n19411), .CLK(clk_i),         .QN(n15481) );
  dffs1  u5_mc_adv_r_reg ( .DIN1(n9329), .CLK(clk_i),         .QN(n36661) );
  dffs1  u5_mc_adv_r1_reg ( .DIN1(n9330), .CLK(clk_i),         .QN(n36636) );
  dffs1  \u5_state_reg[7]  ( .DIN1(n9331), .CLK(clk_i),         .Q(u5_state[7]) );
  dffs1  \u6_wb_data_o_reg[23]  ( .DIN1(n9332), .CLK(clk_i),         .Q(wb_data_o[23]) );
  dffs1  \u3_byte2_reg[7]  ( .DIN1(n9333), .CLK(clk_i),         .QN(n36635) );
  dffs1  \u6_wb_data_o_reg[22]  ( .DIN1(n9334), .CLK(clk_i),         .Q(wb_data_o[22]) );
  dffs1  \u3_byte2_reg[6]  ( .DIN1(n9335), .CLK(clk_i),         .QN(n36633) );
  dffs1  \u6_wb_data_o_reg[21]  ( .DIN1(n9336), .CLK(clk_i),         .Q(wb_data_o[21]) );
  dffs1  \u3_byte2_reg[5]  ( .DIN1(n9337), .CLK(clk_i),         .QN(n36631) );
  dffs1  \u6_wb_data_o_reg[20]  ( .DIN1(n9338), .CLK(clk_i),         .Q(wb_data_o[20]) );
  dffs1  \u3_byte2_reg[4]  ( .DIN1(n9339), .CLK(clk_i),         .QN(n36629) );
  dffs1  \u6_wb_data_o_reg[19]  ( .DIN1(n9340), .CLK(clk_i),         .Q(wb_data_o[19]) );
  dffs1  \u3_byte2_reg[3]  ( .DIN1(n9341), .CLK(clk_i),         .QN(n36627) );
  dffs1  \u6_wb_data_o_reg[18]  ( .DIN1(n9342), .CLK(clk_i),         .Q(wb_data_o[18]) );
  dffs1  \u3_byte2_reg[2]  ( .DIN1(n9343), .CLK(clk_i),         .QN(n36625) );
  dffs1  \u6_wb_data_o_reg[17]  ( .DIN1(n9344), .CLK(clk_i),         .Q(wb_data_o[17]) );
  dffs1  \u3_byte2_reg[1]  ( .DIN1(n9345), .CLK(clk_i),         .QN(n36623) );
  dffs1  \u6_wb_data_o_reg[16]  ( .DIN1(n9346), .CLK(clk_i),         .Q(wb_data_o[16]) );
  dffs1  \u3_byte2_reg[0]  ( .DIN1(n9347), .CLK(clk_i),         .QN(n36621) );
  dffs1  u5_pack_le2_reg ( .DIN1(n9348), .CLK(clk_i),         .QN(n15503) );
  dffs1  \u6_wb_data_o_reg[7]  ( .DIN1(n9349), .CLK(clk_i),         .Q(wb_data_o[7]) );
  dffs1  \u3_byte0_reg[7]  ( .DIN1(n9350), .CLK(clk_i),         .QN(n36619) );
  dffs1  \u6_wb_data_o_reg[6]  ( .DIN1(n9351), .CLK(clk_i),         .Q(wb_data_o[6]) );
  dffs1  \u3_byte0_reg[6]  ( .DIN1(n9352), .CLK(clk_i),         .QN(n36618) );
  dffs1  \u6_wb_data_o_reg[5]  ( .DIN1(n9353), .CLK(clk_i),         .Q(wb_data_o[5]) );
  dffs1  \u3_byte0_reg[5]  ( .DIN1(n9354), .CLK(clk_i),         .QN(n36617) );
  dffs1  \u6_wb_data_o_reg[4]  ( .DIN1(n9355), .CLK(clk_i),         .Q(wb_data_o[4]) );
  dffs1  \u3_byte0_reg[4]  ( .DIN1(n9356), .CLK(clk_i),         .QN(n36616) );
  dffs1  \u6_wb_data_o_reg[3]  ( .DIN1(n9357), .CLK(clk_i),         .Q(wb_data_o[3]) );
  dffs1  \u3_byte0_reg[3]  ( .DIN1(n9358), .CLK(clk_i),         .QN(n36615) );
  dffs1  \u6_wb_data_o_reg[2]  ( .DIN1(n9359), .CLK(clk_i),         .Q(wb_data_o[2]) );
  dffs1  \u3_byte0_reg[2]  ( .DIN1(n9360), .CLK(clk_i),         .QN(n36614) );
  dffs1  \u6_wb_data_o_reg[1]  ( .DIN1(n9361), .CLK(clk_i),         .Q(wb_data_o[1]) );
  dffs1  \u3_byte0_reg[1]  ( .DIN1(n9362), .CLK(clk_i),         .QN(n36613) );
  dffs1  \u6_wb_data_o_reg[0]  ( .DIN1(n9363), .CLK(clk_i),         .Q(wb_data_o[0]) );
  dffs1  \u3_byte0_reg[0]  ( .DIN1(n9364), .CLK(clk_i),         .QN(n36612) );
  dffs1  u5_pack_le0_reg ( .DIN1(n9365), .CLK(clk_i),         .QN(n15504) );
  dffs1  u7_mc_rp_reg ( .DIN1(n19407), .CLK(mc_clk_i),         .Q(mc_rp_pad_o_) );
  dffs1  u7_mc_zz_o_reg ( .DIN1(suspended_o), .CLK(mc_clk_i),         .Q(mc_zz_pad_o) );
  dffs1  u5_suspended_reg ( .DIN1(u5_suspended_d), .CLK(clk_i), .Q(suspended_o), .QN(n15470) );
  dffs1  \u5_state_reg[32]  ( .DIN1(n9367), .CLK(clk_i),         .Q(u5_state[32]) );
  dffs1  \u5_state_reg[62]  ( .DIN1(n9368), .CLK(clk_i),         .Q(u5_state[62]) );
  dffs1  u5_ap_en_reg ( .DIN1(n9369), .CLK(clk_i),         .Q(u5_ap_en) );
  dffs1  \u5_state_reg[4]  ( .DIN1(n9370), .CLK(clk_i),         .Q(u5_state[4]) );
  dffs1  \u5_state_reg[27]  ( .DIN1(n9371), .CLK(clk_i),         .Q(u5_state[27]) );
  dffs1  u5_susp_sel_r_reg ( .DIN1(n9372), .CLK(clk_i),         .Q(u5_susp_sel_r) );
  dffs1  \u5_state_reg[33]  ( .DIN1(n9373), .CLK(clk_i),         .Q(u5_state[33]) );
  dffs1  u0_lmr_req_reg ( .DIN1(n9374), .CLK(clk_i),         .Q(n36662) );
  dffs1  u0_u0_lmr_req_reg ( .DIN1(n9375), .CLK(clk_i),         .QN(n15506) );
  dffs1  u0_u1_lmr_req_reg ( .DIN1(n9376), .CLK(clk_i),         .QN(n36611) );
  dffs1  \u5_state_reg[45]  ( .DIN1(n9377), .CLK(clk_i),         .Q(u5_state[45]) );
  dffs1  u0_lmr_ack_r_reg ( .DIN1(u5_lmr_ack), .CLK(clk_i),         .QN(n4988) );
  dffs1  u5_lmr_ack_reg ( .DIN1(n9378), .CLK(clk_i),         .Q(u5_lmr_ack) );
  dffs1  \u5_state_reg[20]  ( .DIN1(n9379), .CLK(clk_i),         .Q(u5_state[20]) );
  dffs1  \u5_state_reg[19]  ( .DIN1(n9380), .CLK(clk_i),         .Q(u5_state[19]) );
  dffs1  \u5_state_reg[18]  ( .DIN1(n9381), .CLK(clk_i),         .Q(u5_state[18]) );
  dffs1  \u5_state_reg[26]  ( .DIN1(n9382), .CLK(clk_i),         .Q(u5_state[26]) );
  dffs1  \u5_state_reg[24]  ( .DIN1(n9383), .CLK(clk_i),         .Q(u5_state[24]) );
  dffs1  \u5_state_reg[28]  ( .DIN1(n9384), .CLK(clk_i),         .Q(u5_state[28]) );
  dffs1  \u5_state_reg[35]  ( .DIN1(n9385), .CLK(clk_i),         .Q(u5_state[35]) );
  dffs1  \u5_state_reg[34]  ( .DIN1(n9386), .CLK(clk_i),         .Q(u5_state[34]) );
  dffs1  \u5_state_reg[31]  ( .DIN1(n9387), .CLK(clk_i),         .Q(u5_state[31]) );
  dffs1  \u5_state_reg[5]  ( .DIN1(n9388), .CLK(clk_i),         .Q(u5_state[5]) );
  dffs1  \u5_state_reg[49]  ( .DIN1(n9389), .CLK(clk_i),         .Q(u5_state[49]) );
  dffs1  \u5_state_reg[48]  ( .DIN1(n9390), .CLK(clk_i),         .Q(u5_state[48]) );
  dffs1  \u5_state_reg[46]  ( .DIN1(n9391), .CLK(clk_i),         .Q(u5_state[46]) );
  dffs1  \u5_state_reg[61]  ( .DIN1(n9392), .CLK(clk_i),         .Q(u5_state[61]) );
  dffs1  \u5_state_reg[22]  ( .DIN1(n9393), .CLK(clk_i),         .Q(u5_state[22]) );
  dffs1  \u5_state_reg[21]  ( .DIN1(n9394), .CLK(clk_i),         .Q(u5_state[21]) );
  dffs1  u4_rfr_req_reg ( .DIN1(n9395), .CLK(clk_i),         .Q(u4_rfr_req) );
  dffs1  u4_rfr_clr_reg ( .DIN1(n9396), .CLK(clk_i),         .Q(n4611) );
  dffs1  \u4_rfr_cnt_reg[6]  ( .DIN1(n9397), .CLK(clk_i),         .Q(u4_rfr_cnt[6]) );
  dffs1  \u4_rfr_cnt_reg[5]  ( .DIN1(n9398), .CLK(clk_i),         .Q(u4_rfr_cnt[5]) );
  dffs1  \u4_rfr_cnt_reg[4]  ( .DIN1(n9399), .CLK(clk_i),         .Q(u4_rfr_cnt[4]) );
  dffs1  \u4_rfr_cnt_reg[3]  ( .DIN1(n9400), .CLK(clk_i),         .Q(u4_rfr_cnt[3]) );
  dffs1  \u4_rfr_cnt_reg[2]  ( .DIN1(n9401), .CLK(clk_i),         .Q(u4_rfr_cnt[2]) );
  dffs1  \u4_rfr_cnt_reg[1]  ( .DIN1(n9402), .CLK(clk_i),         .Q(u4_rfr_cnt[1]) );
  dffs1  \u4_rfr_cnt_reg[0]  ( .DIN1(n9403), .CLK(clk_i),         .Q(u4_rfr_cnt[0]) );
  dffs1  \u4_rfr_cnt_reg[7]  ( .DIN1(n9404), .CLK(clk_i),         .Q(u4_rfr_cnt[7]) );
  dffs1  u5_rfr_ack_r_reg ( .DIN1(u5_rfr_ack_d), .CLK(clk_i),         .Q(rfr_ack) );
  dffs1  \u5_state_reg[30]  ( .DIN1(n9405), .CLK(clk_i),         .Q(u5_state[30]) );
  dffs1  \u5_state_reg[29]  ( .DIN1(n9406), .CLK(clk_i),         .Q(u5_state[29]) );
  dffs1  \u5_state_reg[23]  ( .DIN1(n9407), .CLK(clk_i),         .Q(u5_state[23]) );
  dffs1  \u5_ir_cnt_reg[3]  ( .DIN1(n9408), .CLK(clk_i),         .QN(n15474) );
  dffs1  u5_ir_cnt_done_reg ( .DIN1(n19413), .CLK(clk_i),         .QN(n15507) );
  dffs1  \u5_ir_cnt_reg[2]  ( .DIN1(n9410), .CLK(clk_i),         .QN(n15508) );
  dffs1  \u5_ir_cnt_reg[1]  ( .DIN1(n9411), .CLK(clk_i),         .Q(u5_ir_cnt[1]) );
  dffs1  \u5_ir_cnt_reg[0]  ( .DIN1(n9412), .CLK(clk_i),         .Q(u5_ir_cnt[0]) );
  dffs1  \u5_state_reg[64]  ( .DIN1(n9413), .CLK(clk_i),         .Q(u5_state[64]) );
  dffs1  \u5_state_reg[6]  ( .DIN1(n9414), .CLK(clk_i),         .Q(u5_state[6]) );
  dffs1  \u5_state_reg[57]  ( .DIN1(n9415), .CLK(clk_i),         .Q(u5_state[57]) );
  dffs1  \u5_state_reg[55]  ( .DIN1(n9416), .CLK(clk_i),         .Q(u5_state[55]) );
  dffs1  \u5_state_reg[54]  ( .DIN1(n9417), .CLK(clk_i),         .Q(u5_state[54]) );
  dffs1  \u5_state_reg[53]  ( .DIN1(n9418), .CLK(clk_i),         .Q(u5_state[53]) );
  dffs1  \u5_state_reg[44]  ( .DIN1(n9419), .CLK(clk_i),         .Q(u5_state[44]) );
  dffs1  \u5_state_reg[43]  ( .DIN1(n9420), .CLK(clk_i),         .Q(u5_state[43]) );
  dffs1  \u5_state_reg[42]  ( .DIN1(n9421), .CLK(clk_i),         .Q(u5_state[42]) );
  dffs1  \u5_state_reg[41]  ( .DIN1(n9422), .CLK(clk_i),         .Q(u5_state[41]) );
  dffs1  \u0_sp_csc_reg[4]  ( .DIN1(n9423), .CLK(clk_i),         .Q(u0_sp_csc[4]) );
  dffs1  \u0_sp_csc_reg[5]  ( .DIN1(n9424), .CLK(clk_i),         .QN(n31263) );
  dffs1  \u0_sp_csc_reg[6]  ( .DIN1(n9425), .CLK(clk_i),         .Q(u0_sp_csc[6]) );
  dffs1  \u0_sp_csc_reg[7]  ( .DIN1(n9426), .CLK(clk_i),         .Q(u0_sp_csc[7]) );
  dffs1  \u0_sp_csc_reg[9]  ( .DIN1(n9427), .CLK(clk_i),         .Q(u0_sp_csc_9) );
  dffs1  \u0_sp_csc_reg[10]  ( .DIN1(n9428), .CLK(clk_i),         .Q(u0_sp_csc_10) );
  dffs1  \u0_sp_tms_reg[0]  ( .DIN1(n9429), .CLK(clk_i),         .Q(u0_sp_tms[0]) );
  dffs1  \u0_sp_tms_reg[1]  ( .DIN1(n9430), .CLK(clk_i),         .Q(u0_sp_tms[1]) );
  dffs1  \u0_sp_tms_reg[2]  ( .DIN1(n9431), .CLK(clk_i),         .Q(u0_sp_tms[2]) );
  dffs1  \u0_sp_tms_reg[3]  ( .DIN1(n9432), .CLK(clk_i),         .Q(u0_sp_tms[3]) );
  dffs1  \u0_sp_tms_reg[4]  ( .DIN1(n9433), .CLK(clk_i),         .Q(u0_sp_tms[4]) );
  dffs1  \u0_sp_tms_reg[5]  ( .DIN1(n9434), .CLK(clk_i),         .Q(u0_sp_tms[5]) );
  dffs1  \u0_sp_tms_reg[6]  ( .DIN1(n9435), .CLK(clk_i),         .Q(u0_sp_tms[6]) );
  dffs1  \u0_sp_tms_reg[7]  ( .DIN1(n9436), .CLK(clk_i),         .Q(u0_sp_tms[7]) );
  dffs1  \u0_sp_tms_reg[8]  ( .DIN1(n9437), .CLK(clk_i),         .Q(u0_sp_tms[8]) );
  dffs1  \u0_sp_tms_reg[9]  ( .DIN1(n9438), .CLK(clk_i),         .Q(u0_sp_tms[9]) );
  dffs1  \u0_sp_tms_reg[10]  ( .DIN1(n9439), .CLK(clk_i),         .Q(u0_sp_tms[10]) );
  dffs1  \u0_sp_tms_reg[11]  ( .DIN1(n9440), .CLK(clk_i),         .Q(u0_sp_tms[11]) );
  dffs1  \u0_sp_tms_reg[12]  ( .DIN1(n9441), .CLK(clk_i),         .Q(u0_sp_tms[12]) );
  dffs1  \u0_sp_tms_reg[13]  ( .DIN1(n9442), .CLK(clk_i),         .Q(u0_sp_tms[13]) );
  dffs1  \u0_sp_tms_reg[14]  ( .DIN1(n9443), .CLK(clk_i),         .Q(u0_sp_tms[14]) );
  dffs1  \u0_sp_tms_reg[15]  ( .DIN1(n9444), .CLK(clk_i),         .Q(u0_sp_tms[15]) );
  dffs1  \u0_sp_tms_reg[16]  ( .DIN1(n9445), .CLK(clk_i),         .Q(u0_sp_tms[16]) );
  dffs1  \u0_sp_tms_reg[17]  ( .DIN1(n9446), .CLK(clk_i),         .Q(u0_sp_tms[17]) );
  dffs1  \u0_sp_tms_reg[18]  ( .DIN1(n9447), .CLK(clk_i),         .Q(u0_sp_tms[18]) );
  dffs1  \u0_sp_tms_reg[19]  ( .DIN1(n9448), .CLK(clk_i),         .Q(u0_sp_tms[19]) );
  dffs1  \u0_sp_tms_reg[20]  ( .DIN1(n9449), .CLK(clk_i),         .Q(u0_sp_tms[20]) );
  dffs1  \u0_sp_tms_reg[21]  ( .DIN1(n9450), .CLK(clk_i),         .Q(u0_sp_tms[21]) );
  dffs1  \u0_sp_tms_reg[22]  ( .DIN1(n9451), .CLK(clk_i),         .Q(u0_sp_tms[22]) );
  dffs1  \u0_sp_tms_reg[23]  ( .DIN1(n9452), .CLK(clk_i),         .Q(u0_sp_tms[23]) );
  dffs1  \u0_sp_tms_reg[24]  ( .DIN1(n9453), .CLK(clk_i),         .Q(u0_sp_tms[24]) );
  dffs1  \u0_sp_tms_reg[25]  ( .DIN1(n9454), .CLK(clk_i),         .Q(u0_sp_tms[25]) );
  dffs1  \u0_sp_tms_reg[26]  ( .DIN1(n9455), .CLK(clk_i),         .Q(u0_sp_tms[26]) );
  dffs1  \u0_sp_tms_reg[27]  ( .DIN1(n9456), .CLK(clk_i),         .Q(u0_sp_tms[27]) );
  dffs1  u0_u0_init_req_reg ( .DIN1(n9457), .CLK(clk_i),         .QN(n15509) );
  dffs1  u0_u0_inited_reg ( .DIN1(n9458), .CLK(clk_i),         .QN(n15510) );
  dffs1  \u0_spec_req_cs_reg[0]  ( .DIN1(n9459), .CLK(clk_i),         .Q(u0_spec_req_cs[0]) );
  dffs1  u0_init_req_reg ( .DIN1(n9460), .CLK(clk_i),         .Q(u0_init_req) );
  dffs1  u0_u1_init_req_reg ( .DIN1(n9461), .CLK(clk_i),         .QN(n36608) );
  dffs1  u0_u1_inited_reg ( .DIN1(n9462), .CLK(clk_i),         .QN(n15483) );
  dffs1  \u0_spec_req_cs_reg[1]  ( .DIN1(n9463), .CLK(clk_i),         .Q(u0_spec_req_cs[1]) );
  dffs1  u0_sreq_cs_le_reg ( .DIN1(n9464), .CLK(clk_i),         .QN(n15511) );
  dffs1  u0_init_ack_r_reg ( .DIN1(u5_init_ack), .CLK(clk_i),         .QN(n4989) );
  dffs1  \u5_state_reg[25]  ( .DIN1(n9465), .CLK(clk_i),         .Q(u5_state[25]) );
  dffs1  \u5_state_reg[9]  ( .DIN1(n9466), .CLK(clk_i),         .Q(u5_state[9]) );
  dffs1  \u5_state_reg[1]  ( .DIN1(n9467), .CLK(clk_i),         .Q(u5_state[1]) );
  dffs1  \u5_state_reg[3]  ( .DIN1(n9468), .CLK(clk_i),         .Q(u5_state[3]) );
  dffs1  u5_wb_stb_first_reg ( .DIN1(n9469), .CLK(clk_i),         .Q(u5_wb_stb_first) );
  dffs1  u6_wb_first_r_reg ( .DIN1(n9470), .CLK(clk_i),         .QN(n36607) );
  dffs1  u6_wb_err_reg ( .DIN1(n9471), .CLK(clk_i),         .Q(wb_err_o) );
  dffs1  \u5_state_reg[65]  ( .DIN1(n9472), .CLK(clk_i),         .Q(u5_state[65]) );
  dffs1  \u5_state_reg[51]  ( .DIN1(n9473), .CLK(clk_i),         .Q(u5_state[51]) );
  dffs1  u5_tmr2_done_reg ( .DIN1(n9474), .CLK(clk_i),         .Q(u5_tmr2_done) );
  dffs1  \u5_timer2_reg[8]  ( .DIN1(n9475), .CLK(clk_i),         .Q(u5_timer2[8]) );
  dffs1  \u0_csc_reg[1]  ( .DIN1(n9476), .CLK(clk_i),         .Q(u0_csc[1]) );
  dffs1  \u6_wb_data_o_reg[24]  ( .DIN1(n9477), .CLK(clk_i),         .Q(wb_data_o[24]) );
  dffs1  \u6_wb_data_o_reg[25]  ( .DIN1(n9478), .CLK(clk_i),         .Q(wb_data_o[25]) );
  dffs1  \u6_wb_data_o_reg[26]  ( .DIN1(n9479), .CLK(clk_i),         .Q(wb_data_o[26]) );
  dffs1  \u6_wb_data_o_reg[27]  ( .DIN1(n9480), .CLK(clk_i),         .Q(wb_data_o[27]) );
  dffs1  \u6_wb_data_o_reg[28]  ( .DIN1(n9481), .CLK(clk_i),         .Q(wb_data_o[28]) );
  dffs1  \u6_wb_data_o_reg[29]  ( .DIN1(n9482), .CLK(clk_i),         .Q(wb_data_o[29]) );
  dffs1  \u6_wb_data_o_reg[30]  ( .DIN1(n9483), .CLK(clk_i),         .Q(wb_data_o[30]) );
  dffs1  \u6_wb_data_o_reg[31]  ( .DIN1(n9484), .CLK(clk_i),         .Q(wb_data_o[31]) );
  dffs1  \u0_csc_reg[2]  ( .DIN1(n9485), .CLK(clk_i),         .Q(u0_csc[2]) );
  dffs1  \u0_csc_reg[3]  ( .DIN1(n9486), .CLK(clk_i),         .Q(u0_csc[3]) );
  dffs1  \u0_csc_reg[4]  ( .DIN1(n9487), .CLK(clk_i),         .Q(u0_csc[4]) );
  dffs1  \u0_csc_reg[5]  ( .DIN1(n9488), .CLK(clk_i),         .Q(u0_csc[5]) );
  dffs1  \u0_csc_reg[6]  ( .DIN1(n9489), .CLK(clk_i),         .Q(u0_csc[6]) );
  dffs1  \u0_csc_reg[7]  ( .DIN1(n9490), .CLK(clk_i),         .Q(u0_csc[7]) );
  dffs1  \u0_csc_reg[9]  ( .DIN1(n9491), .CLK(clk_i),         .Q(u0_csc_9) );
  dffs1  \u0_csc_reg[10]  ( .DIN1(n9492), .CLK(clk_i),         .Q(u0_csc_10) );
  dffs1  \u0_tms_reg[0]  ( .DIN1(n9493), .CLK(clk_i),         .Q(u0_tms[0]) );
  dffs1  \u0_tms_reg[1]  ( .DIN1(n9494), .CLK(clk_i),         .Q(u0_tms[1]) );
  dffs1  \u0_tms_reg[2]  ( .DIN1(n9495), .CLK(clk_i),         .Q(u0_tms[2]) );
  dffs1  \u0_tms_reg[3]  ( .DIN1(n9496), .CLK(clk_i),         .Q(u0_tms[3]) );
  dffs1  \u0_tms_reg[4]  ( .DIN1(n9497), .CLK(clk_i),         .Q(u0_tms[4]) );
  dffs1  \u0_tms_reg[5]  ( .DIN1(n9498), .CLK(clk_i),         .Q(u0_tms[5]) );
  dffs1  \u0_tms_reg[6]  ( .DIN1(n9499), .CLK(clk_i),         .Q(u0_tms[6]) );
  dffs1  \u0_tms_reg[7]  ( .DIN1(n9500), .CLK(clk_i),         .Q(u0_tms[7]) );
  dffs1  \u0_tms_reg[8]  ( .DIN1(n9501), .CLK(clk_i),         .Q(u0_tms[8]) );
  dffs1  \u0_tms_reg[9]  ( .DIN1(n9502), .CLK(clk_i),         .Q(u0_tms[9]) );
  dffs1  \u0_tms_reg[10]  ( .DIN1(n9503), .CLK(clk_i),         .Q(u0_tms[10]) );
  dffs1  \u0_tms_reg[11]  ( .DIN1(n9504), .CLK(clk_i),         .Q(u0_tms[11]) );
  dffs1  \u0_tms_reg[12]  ( .DIN1(n9505), .CLK(clk_i),         .Q(u0_tms[12]) );
  dffs1  \u0_tms_reg[13]  ( .DIN1(n9506), .CLK(clk_i),         .Q(u0_tms[13]) );
  dffs1  \u0_tms_reg[14]  ( .DIN1(n9507), .CLK(clk_i),         .Q(u0_tms[14]) );
  dffs1  \u0_tms_reg[15]  ( .DIN1(n9508), .CLK(clk_i),         .Q(u0_tms[15]) );
  dffs1  \u0_tms_reg[16]  ( .DIN1(n9509), .CLK(clk_i),         .Q(u0_tms[16]) );
  dffs1  \u0_tms_reg[17]  ( .DIN1(n9510), .CLK(clk_i),         .Q(u0_tms[17]) );
  dffs1  \u0_tms_reg[18]  ( .DIN1(n9511), .CLK(clk_i),         .Q(u0_tms[18]) );
  dffs1  \u0_tms_reg[19]  ( .DIN1(n9512), .CLK(clk_i),         .Q(u0_tms[19]) );
  dffs1  \u0_tms_reg[20]  ( .DIN1(n9513), .CLK(clk_i),         .Q(u0_tms[20]) );
  dffs1  \u0_tms_reg[21]  ( .DIN1(n9514), .CLK(clk_i),         .Q(u0_tms[21]) );
  dffs1  \u0_tms_reg[22]  ( .DIN1(n9515), .CLK(clk_i),         .Q(u0_tms[22]) );
  dffs1  \u0_tms_reg[23]  ( .DIN1(n9516), .CLK(clk_i),         .Q(u0_tms[23]) );
  dffs1  \u0_tms_reg[24]  ( .DIN1(n9517), .CLK(clk_i),         .Q(u0_tms[24]) );
  dffs1  \u0_tms_reg[25]  ( .DIN1(n9518), .CLK(clk_i),         .Q(u0_tms[25]) );
  dffs1  \u0_tms_reg[26]  ( .DIN1(n9519), .CLK(clk_i),         .Q(u0_tms[26]) );
  dffs1  \u0_tms_reg[27]  ( .DIN1(n9520), .CLK(clk_i),         .Q(u0_tms[27]) );
  dffs1  u0_wp_err_reg ( .DIN1(n9521), .CLK(clk_i),         .QN(n36606) );
  dffs1  u5_lookup_ready2_reg ( .DIN1(n9522), .CLK(clk_i),         .QN(n4990) );
  dffs1  u5_lookup_ready1_reg ( .DIN1(n9523), .CLK(clk_i),         .Q(n4629) );
  dffs1  \u0_cs_reg[7]  ( .DIN1(n9524), .CLK(clk_i),         .QN(n15495) );
  dffs1  \u0_cs_reg[6]  ( .DIN1(n9525), .CLK(clk_i),         .QN(n15496) );
  dffs1  \u0_cs_reg[5]  ( .DIN1(n9526), .CLK(clk_i),         .QN(n15497) );
  dffs1  \u0_cs_reg[4]  ( .DIN1(n9527), .CLK(clk_i),         .QN(n15498) );
  dffs1  \u0_cs_reg[3]  ( .DIN1(n9528), .CLK(clk_i),         .QN(n15499) );
  dffs1  \u0_cs_reg[2]  ( .DIN1(n9529), .CLK(clk_i),         .QN(n15500) );
  dffs1  \u0_cs_reg[1]  ( .DIN1(n9530), .CLK(clk_i),         .Q(u0_cs[1]) );
  dffs1  \u0_cs_reg[0]  ( .DIN1(n9531), .CLK(clk_i),         .Q(u0_cs[0]) );
  dffs1  u5_cs_le_r_reg ( .DIN1(n9532), .CLK(clk_i),         .Q(n4625) );
  dffs1  u5_cs_le_r1_reg ( .DIN1(u5_cs_le), .CLK(clk_i),         .Q(n9532) );
  dffs1  u5_cs_le_reg ( .DIN1(n9533), .CLK(clk_i),         .Q(u5_cs_le) );
  dffs1  \u5_state_reg[17]  ( .DIN1(n9534), .CLK(clk_i),         .Q(u5_state[17]) );
  dffs1  \u5_state_reg[50]  ( .DIN1(n9535), .CLK(clk_i),         .Q(u5_state[50]) );
  dffs1  \u5_state_reg[12]  ( .DIN1(n9536), .CLK(clk_i),         .Q(u5_state[12]) );
  dffs1  u5_burst_act_rd_reg ( .DIN1(n9537), .CLK(clk_i),         .Q(n4771) );
  dffs1  \u5_burst_cnt_reg[10]  ( .DIN1(n9538), .CLK(clk_i),         .Q(u5_burst_cnt[10]) );
  dffs1  \u5_ack_cnt_reg[2]  ( .DIN1(n9539), .CLK(clk_i),         .Q(u5_ack_cnt[2]) );
  dffs1  \u5_ack_cnt_reg[1]  ( .DIN1(n9540), .CLK(clk_i),         .Q(u5_ack_cnt[1]) );
  dffs1  \u5_ack_cnt_reg[3]  ( .DIN1(n9541), .CLK(clk_i),         .Q(u5_ack_cnt[3]) );
  dffs1  \u5_ack_cnt_reg[0]  ( .DIN1(n9542), .CLK(clk_i),         .Q(u5_ack_cnt[0]) );
  dffs1  \u3_u0_r3_reg[31]  ( .DIN1(n9543), .CLK(clk_i),         .QN(n31259) );
  dffs1  \u3_u0_r3_reg[30]  ( .DIN1(n9544), .CLK(clk_i),         .QN(n31255) );
  dffs1  \u3_u0_r3_reg[29]  ( .DIN1(n9545), .CLK(clk_i),         .QN(n31251) );
  dffs1  \u3_u0_r3_reg[28]  ( .DIN1(n9546), .CLK(clk_i),         .QN(n31247) );
  dffs1  \u3_u0_r3_reg[27]  ( .DIN1(n9547), .CLK(clk_i),         .QN(n31243) );
  dffs1  \u3_u0_r3_reg[26]  ( .DIN1(n9548), .CLK(clk_i),         .QN(n31239) );
  dffs1  \u3_u0_r3_reg[25]  ( .DIN1(n9549), .CLK(clk_i),         .QN(n31235) );
  dffs1  \u3_u0_r3_reg[24]  ( .DIN1(n9550), .CLK(clk_i),         .QN(n31231) );
  dffs1  \u3_u0_r3_reg[23]  ( .DIN1(n9551), .CLK(clk_i),         .QN(n31227) );
  dffs1  \u3_u0_r3_reg[22]  ( .DIN1(n9552), .CLK(clk_i),         .QN(n31223) );
  dffs1  \u3_u0_r3_reg[21]  ( .DIN1(n9553), .CLK(clk_i),         .QN(n31219) );
  dffs1  \u3_u0_r3_reg[20]  ( .DIN1(n9554), .CLK(clk_i),         .QN(n31215) );
  dffs1  \u3_u0_r3_reg[19]  ( .DIN1(n9555), .CLK(clk_i),         .QN(n31211) );
  dffs1  \u3_u0_r3_reg[18]  ( .DIN1(n9556), .CLK(clk_i),         .QN(n31207) );
  dffs1  \u3_u0_r3_reg[17]  ( .DIN1(n9557), .CLK(clk_i),         .QN(n31203) );
  dffs1  \u3_u0_r3_reg[16]  ( .DIN1(n9558), .CLK(clk_i),         .QN(n31199) );
  dffs1  \u3_u0_r3_reg[15]  ( .DIN1(n9559), .CLK(clk_i),         .QN(n31195) );
  dffs1  \u3_u0_r3_reg[14]  ( .DIN1(n9560), .CLK(clk_i),         .QN(n31191) );
  dffs1  \u3_u0_r3_reg[13]  ( .DIN1(n9561), .CLK(clk_i),         .QN(n31187) );
  dffs1  \u3_u0_r3_reg[12]  ( .DIN1(n9562), .CLK(clk_i),         .QN(n31183) );
  dffs1  \u3_u0_r3_reg[11]  ( .DIN1(n9563), .CLK(clk_i),         .QN(n31179) );
  dffs1  \u3_u0_r3_reg[10]  ( .DIN1(n9564), .CLK(clk_i),         .QN(n31175) );
  dffs1  \u3_u0_r3_reg[9]  ( .DIN1(n9565), .CLK(clk_i),         .QN(n31171) );
  dffs1  \u3_u0_r3_reg[8]  ( .DIN1(n9566), .CLK(clk_i),         .QN(n31167) );
  dffs1  \u3_u0_r3_reg[7]  ( .DIN1(n9567), .CLK(clk_i),         .QN(n31163) );
  dffs1  \u3_u0_r3_reg[6]  ( .DIN1(n9568), .CLK(clk_i),         .QN(n31159) );
  dffs1  \u3_u0_r3_reg[5]  ( .DIN1(n9569), .CLK(clk_i),         .QN(n31155) );
  dffs1  \u3_u0_r3_reg[4]  ( .DIN1(n9570), .CLK(clk_i),         .QN(n31151) );
  dffs1  \u3_u0_r3_reg[3]  ( .DIN1(n9571), .CLK(clk_i),         .QN(n31147) );
  dffs1  \u3_u0_r3_reg[2]  ( .DIN1(n9572), .CLK(clk_i),         .QN(n31143) );
  dffs1  \u3_u0_r3_reg[1]  ( .DIN1(n9573), .CLK(clk_i),         .QN(n31139) );
  dffs1  \u3_u0_r3_reg[0]  ( .DIN1(n9574), .CLK(clk_i),         .QN(n31135) );
  dffs1  \u3_u0_r2_reg[31]  ( .DIN1(n9575), .CLK(clk_i),         .QN(n31260) );
  dffs1  \u3_u0_r2_reg[30]  ( .DIN1(n9576), .CLK(clk_i),         .QN(n31256) );
  dffs1  \u3_u0_r2_reg[29]  ( .DIN1(n9577), .CLK(clk_i),         .QN(n31252) );
  dffs1  \u3_u0_r2_reg[28]  ( .DIN1(n9578), .CLK(clk_i),         .QN(n31248) );
  dffs1  \u3_u0_r2_reg[27]  ( .DIN1(n9579), .CLK(clk_i),         .QN(n31244) );
  dffs1  \u3_u0_r2_reg[26]  ( .DIN1(n9580), .CLK(clk_i),         .QN(n31240) );
  dffs1  \u3_u0_r2_reg[25]  ( .DIN1(n9581), .CLK(clk_i),         .QN(n31236) );
  dffs1  \u3_u0_r2_reg[24]  ( .DIN1(n9582), .CLK(clk_i),         .QN(n31232) );
  dffs1  \u3_u0_r2_reg[23]  ( .DIN1(n9583), .CLK(clk_i),         .QN(n31228) );
  dffs1  \u3_u0_r2_reg[22]  ( .DIN1(n9584), .CLK(clk_i),         .QN(n31224) );
  dffs1  \u3_u0_r2_reg[21]  ( .DIN1(n9585), .CLK(clk_i),         .QN(n31220) );
  dffs1  \u3_u0_r2_reg[20]  ( .DIN1(n9586), .CLK(clk_i),         .QN(n31216) );
  dffs1  \u3_u0_r2_reg[19]  ( .DIN1(n9587), .CLK(clk_i),         .QN(n31212) );
  dffs1  \u3_u0_r2_reg[18]  ( .DIN1(n9588), .CLK(clk_i),         .QN(n31208) );
  dffs1  \u3_u0_r2_reg[17]  ( .DIN1(n9589), .CLK(clk_i),         .QN(n31204) );
  dffs1  \u3_u0_r2_reg[16]  ( .DIN1(n9590), .CLK(clk_i),         .QN(n31200) );
  dffs1  \u3_u0_r2_reg[15]  ( .DIN1(n9591), .CLK(clk_i),         .QN(n31196) );
  dffs1  \u3_u0_r2_reg[14]  ( .DIN1(n9592), .CLK(clk_i),         .QN(n31192) );
  dffs1  \u3_u0_r2_reg[13]  ( .DIN1(n9593), .CLK(clk_i),         .QN(n31188) );
  dffs1  \u3_u0_r2_reg[12]  ( .DIN1(n9594), .CLK(clk_i),         .QN(n31184) );
  dffs1  \u3_u0_r2_reg[11]  ( .DIN1(n9595), .CLK(clk_i),         .QN(n31180) );
  dffs1  \u3_u0_r2_reg[10]  ( .DIN1(n9596), .CLK(clk_i),         .QN(n31176) );
  dffs1  \u3_u0_r2_reg[9]  ( .DIN1(n9597), .CLK(clk_i),         .QN(n31172) );
  dffs1  \u3_u0_r2_reg[8]  ( .DIN1(n9598), .CLK(clk_i),         .QN(n31168) );
  dffs1  \u3_u0_r2_reg[7]  ( .DIN1(n9599), .CLK(clk_i),         .QN(n31164) );
  dffs1  \u3_u0_r2_reg[6]  ( .DIN1(n9600), .CLK(clk_i),         .QN(n31160) );
  dffs1  \u3_u0_r2_reg[5]  ( .DIN1(n9601), .CLK(clk_i),         .QN(n31156) );
  dffs1  \u3_u0_r2_reg[4]  ( .DIN1(n9602), .CLK(clk_i),         .QN(n31152) );
  dffs1  \u3_u0_r2_reg[3]  ( .DIN1(n9603), .CLK(clk_i),         .QN(n31148) );
  dffs1  \u3_u0_r2_reg[2]  ( .DIN1(n9604), .CLK(clk_i),         .QN(n31144) );
  dffs1  \u3_u0_r2_reg[1]  ( .DIN1(n9605), .CLK(clk_i),         .QN(n31140) );
  dffs1  \u3_u0_r2_reg[0]  ( .DIN1(n9606), .CLK(clk_i),         .QN(n31136) );
  dffs1  \u3_u0_r1_reg[31]  ( .DIN1(n9607), .CLK(clk_i),         .QN(n31261) );
  dffs1  \u3_u0_r1_reg[30]  ( .DIN1(n9608), .CLK(clk_i),         .QN(n31257) );
  dffs1  \u3_u0_r1_reg[29]  ( .DIN1(n9609), .CLK(clk_i),         .QN(n31253) );
  dffs1  \u3_u0_r1_reg[28]  ( .DIN1(n9610), .CLK(clk_i),         .QN(n31249) );
  dffs1  \u3_u0_r1_reg[27]  ( .DIN1(n9611), .CLK(clk_i),         .QN(n31245) );
  dffs1  \u3_u0_r1_reg[26]  ( .DIN1(n9612), .CLK(clk_i),         .QN(n31241) );
  dffs1  \u3_u0_r1_reg[25]  ( .DIN1(n9613), .CLK(clk_i),         .QN(n31237) );
  dffs1  \u3_u0_r1_reg[24]  ( .DIN1(n9614), .CLK(clk_i),         .QN(n31233) );
  dffs1  \u3_u0_r1_reg[23]  ( .DIN1(n9615), .CLK(clk_i),         .QN(n31229) );
  dffs1  \u3_u0_r1_reg[22]  ( .DIN1(n9616), .CLK(clk_i),         .QN(n31225) );
  dffs1  \u3_u0_r1_reg[21]  ( .DIN1(n9617), .CLK(clk_i),         .QN(n31221) );
  dffs1  \u3_u0_r1_reg[20]  ( .DIN1(n9618), .CLK(clk_i),         .QN(n31217) );
  dffs1  \u3_u0_r1_reg[19]  ( .DIN1(n9619), .CLK(clk_i),         .QN(n31213) );
  dffs1  \u3_u0_r1_reg[18]  ( .DIN1(n9620), .CLK(clk_i),         .QN(n31209) );
  dffs1  \u3_u0_r1_reg[17]  ( .DIN1(n9621), .CLK(clk_i),         .QN(n31205) );
  dffs1  \u3_u0_r1_reg[16]  ( .DIN1(n9622), .CLK(clk_i),         .QN(n31201) );
  dffs1  \u3_u0_r1_reg[15]  ( .DIN1(n9623), .CLK(clk_i),         .QN(n31197) );
  dffs1  \u3_u0_r1_reg[14]  ( .DIN1(n9624), .CLK(clk_i),         .QN(n31193) );
  dffs1  \u3_u0_r1_reg[13]  ( .DIN1(n9625), .CLK(clk_i),         .QN(n31189) );
  dffs1  \u3_u0_r1_reg[12]  ( .DIN1(n9626), .CLK(clk_i),         .QN(n31185) );
  dffs1  \u3_u0_r1_reg[11]  ( .DIN1(n9627), .CLK(clk_i),         .QN(n31181) );
  dffs1  \u3_u0_r1_reg[10]  ( .DIN1(n9628), .CLK(clk_i),         .QN(n31177) );
  dffs1  \u3_u0_r1_reg[9]  ( .DIN1(n9629), .CLK(clk_i),         .QN(n31173) );
  dffs1  \u3_u0_r1_reg[8]  ( .DIN1(n9630), .CLK(clk_i),         .QN(n31169) );
  dffs1  \u3_u0_r1_reg[7]  ( .DIN1(n9631), .CLK(clk_i),         .QN(n31165) );
  dffs1  \u3_u0_r1_reg[6]  ( .DIN1(n9632), .CLK(clk_i),         .QN(n31161) );
  dffs1  \u3_u0_r1_reg[5]  ( .DIN1(n9633), .CLK(clk_i),         .QN(n31157) );
  dffs1  \u3_u0_r1_reg[4]  ( .DIN1(n9634), .CLK(clk_i),         .QN(n31153) );
  dffs1  \u3_u0_r1_reg[3]  ( .DIN1(n9635), .CLK(clk_i),         .QN(n31149) );
  dffs1  \u3_u0_r1_reg[2]  ( .DIN1(n9636), .CLK(clk_i),         .QN(n31145) );
  dffs1  \u3_u0_r1_reg[1]  ( .DIN1(n9637), .CLK(clk_i),         .QN(n31141) );
  dffs1  \u3_u0_r1_reg[0]  ( .DIN1(n9638), .CLK(clk_i),         .QN(n31137) );
  dffs1  \u3_u0_r0_reg[31]  ( .DIN1(n9639), .CLK(clk_i),         .QN(n31262) );
  dffs1  \u3_u0_r0_reg[30]  ( .DIN1(n9640), .CLK(clk_i),         .QN(n31258) );
  dffs1  \u3_u0_r0_reg[29]  ( .DIN1(n9641), .CLK(clk_i),         .QN(n31254) );
  dffs1  \u3_u0_r0_reg[28]  ( .DIN1(n9642), .CLK(clk_i),         .QN(n31250) );
  dffs1  \u3_u0_r0_reg[27]  ( .DIN1(n9643), .CLK(clk_i),         .QN(n31246) );
  dffs1  \u3_u0_r0_reg[26]  ( .DIN1(n9644), .CLK(clk_i),         .QN(n31242) );
  dffs1  \u3_u0_r0_reg[25]  ( .DIN1(n9645), .CLK(clk_i),         .QN(n31238) );
  dffs1  \u3_u0_r0_reg[24]  ( .DIN1(n9646), .CLK(clk_i),         .QN(n31234) );
  dffs1  \u3_u0_r0_reg[23]  ( .DIN1(n9647), .CLK(clk_i),         .QN(n31230) );
  dffs1  \u3_u0_r0_reg[22]  ( .DIN1(n9648), .CLK(clk_i),         .QN(n31226) );
  dffs1  \u3_u0_r0_reg[21]  ( .DIN1(n9649), .CLK(clk_i),         .QN(n31222) );
  dffs1  \u3_u0_r0_reg[20]  ( .DIN1(n9650), .CLK(clk_i),         .QN(n31218) );
  dffs1  \u3_u0_r0_reg[19]  ( .DIN1(n9651), .CLK(clk_i),         .QN(n31214) );
  dffs1  \u3_u0_r0_reg[18]  ( .DIN1(n9652), .CLK(clk_i),         .QN(n31210) );
  dffs1  \u3_u0_r0_reg[17]  ( .DIN1(n9653), .CLK(clk_i),         .QN(n31206) );
  dffs1  \u3_u0_r0_reg[16]  ( .DIN1(n9654), .CLK(clk_i),         .QN(n31202) );
  dffs1  \u3_u0_r0_reg[15]  ( .DIN1(n9655), .CLK(clk_i),         .QN(n31198) );
  dffs1  \u3_u0_r0_reg[14]  ( .DIN1(n9656), .CLK(clk_i),         .QN(n31194) );
  dffs1  \u3_u0_r0_reg[13]  ( .DIN1(n9657), .CLK(clk_i),         .QN(n31190) );
  dffs1  \u3_u0_r0_reg[12]  ( .DIN1(n9658), .CLK(clk_i),         .QN(n31186) );
  dffs1  \u3_u0_r0_reg[11]  ( .DIN1(n9659), .CLK(clk_i),         .QN(n31182) );
  dffs1  \u3_u0_r0_reg[10]  ( .DIN1(n9660), .CLK(clk_i),         .QN(n31178) );
  dffs1  \u3_u0_r0_reg[9]  ( .DIN1(n9661), .CLK(clk_i),         .QN(n31174) );
  dffs1  \u3_u0_r0_reg[8]  ( .DIN1(n9662), .CLK(clk_i),         .QN(n31170) );
  dffs1  \u3_u0_r0_reg[7]  ( .DIN1(n9663), .CLK(clk_i),         .QN(n31166) );
  dffs1  \u3_u0_r0_reg[6]  ( .DIN1(n9664), .CLK(clk_i),         .QN(n31162) );
  dffs1  \u3_u0_r0_reg[5]  ( .DIN1(n9665), .CLK(clk_i),         .QN(n31158) );
  dffs1  \u3_u0_r0_reg[4]  ( .DIN1(n9666), .CLK(clk_i),         .QN(n31154) );
  dffs1  \u3_u0_r0_reg[3]  ( .DIN1(n9667), .CLK(clk_i),         .QN(n31150) );
  dffs1  \u3_u0_r0_reg[2]  ( .DIN1(n9668), .CLK(clk_i),         .QN(n31146) );
  dffs1  \u3_u0_r0_reg[1]  ( .DIN1(n9669), .CLK(clk_i),         .QN(n31142) );
  dffs1  \u3_u0_r0_reg[0]  ( .DIN1(n9670), .CLK(clk_i),         .QN(n31138) );
  dffs1  \u3_u0_wr_adr_reg[2]  ( .DIN1(n9671), .CLK(clk_i),         .QN(n15478) );
  dffs1  \u3_u0_wr_adr_reg[1]  ( .DIN1(n9672), .CLK(clk_i),         .QN(n15479) );
  dffs1  \u3_u0_wr_adr_reg[0]  ( .DIN1(n9673), .CLK(clk_i),         .Q(n36595) );
  dffs1  \u3_u0_wr_adr_reg[3]  ( .DIN1(n9674), .CLK(clk_i),         .QN(n15477) );
  dffs1  u5_dv_r_reg ( .DIN1(u5_dv), .CLK(clk_i), .QN(n4987)
         );
  dffs1  u5_cke_o_del_reg ( .DIN1(n9675), .CLK(clk_i),         .Q(n4770) );
  dffs1  u5_cke_o_r2_reg ( .DIN1(n9676), .CLK(clk_i),         .Q(n9675) );
  dffs1  u5_cke_o_r1_reg ( .DIN1(mc_cke_pad_o_), .CLK(clk_i),         .Q(n9676) );
  dffs1  u5_cke__reg ( .DIN1(n9677), .CLK(clk_i), .Q(
        mc_cke_pad_o_) );
  dffs1  \u5_state_reg[2]  ( .DIN1(n9678), .CLK(clk_i),         .Q(u5_state[2]) );
  dffs1  u5_cmd_asserted2_reg ( .DIN1(n9679), .CLK(clk_i),         .Q(u5_cmd_asserted2) );
  dffs1  u5_cmd_asserted_reg ( .DIN1(n9680), .CLK(clk_i),         .QN(n15512) );
  dffs1  \u5_cmd_del_reg[3]  ( .DIN1(n9681), .CLK(clk_i),         .QN(n4997) );
  dffs1  \u5_cmd_r_reg[3]  ( .DIN1(n9682), .CLK(clk_i),         .Q(n9681) );
  dffs1  \u5_state_reg[16]  ( .DIN1(n9683), .CLK(clk_i),         .Q(u5_state[16]) );
  dffs1  \u5_state_reg[15]  ( .DIN1(n9684), .CLK(clk_i),         .Q(u5_state[15]) );
  dffs1  \u5_state_reg[11]  ( .DIN1(n9685), .CLK(clk_i),         .Q(u5_state[11]) );
  dffs1  \u5_state_reg[10]  ( .DIN1(n9686), .CLK(clk_i),         .Q(u5_state[10]) );
  dffs1  u5_tmr_done_reg ( .DIN1(n19412), .CLK(clk_i),         .Q(u5_tmr_done) );
  dffs1  \u5_timer_reg[1]  ( .DIN1(n9688), .CLK(clk_i),         .Q(u5_timer[1]) );
  dffs1  u7_mc_c_oe_reg ( .DIN1(n9689), .CLK(mc_clk_i),         .Q(mc_coe_pad_coe_o) );
  dffs1  u5_mc_c_oe_reg ( .DIN1(n9690), .CLK(clk_i),         .Q(n9689) );
  dffs1  \u5_state_reg[40]  ( .DIN1(n9691), .CLK(clk_i),         .Q(u5_state[40]) );
  dffs1  \u5_state_reg[39]  ( .DIN1(n9692), .CLK(clk_i),         .Q(u5_state[39]) );
  dffs1  \u5_state_reg[38]  ( .DIN1(n9693), .CLK(clk_i),         .Q(u5_state[38]) );
  dffs1  \u5_state_reg[37]  ( .DIN1(n9694), .CLK(clk_i),         .Q(u5_state[37]) );
  dffs1  \u5_state_reg[0]  ( .DIN1(n9695), .CLK(clk_i),         .Q(u5_state[0]) );
  dffs1  \u5_state_reg[13]  ( .DIN1(n9696), .CLK(clk_i),         .Q(u5_state[13]) );
  dffs1  \u5_state_reg[14]  ( .DIN1(n9697), .CLK(clk_i),         .Q(u5_state[14]) );
  dffs1  \u5_state_reg[36]  ( .DIN1(n9698), .CLK(clk_i),         .Q(u5_state[36]) );
  dffs1  \u5_state_reg[47]  ( .DIN1(n9699), .CLK(clk_i),         .Q(u5_state[47]) );
  dffs1  \u5_state_reg[52]  ( .DIN1(n9700), .CLK(clk_i),         .Q(u5_state[52]) );
  dffs1  \u5_state_reg[56]  ( .DIN1(n9701), .CLK(clk_i),         .Q(u5_state[56]) );
  dffs1  \u5_state_reg[58]  ( .DIN1(n9702), .CLK(clk_i),         .Q(u5_state[58]) );
  dffs1  \u5_state_reg[59]  ( .DIN1(n9703), .CLK(clk_i),         .Q(u5_state[59]) );
  dffs1  \u5_state_reg[60]  ( .DIN1(n9704), .CLK(clk_i),         .Q(u5_state[60]) );
  dffs1  \u5_state_reg[63]  ( .DIN1(n9705), .CLK(clk_i),         .Q(u5_state[63]) );
  dffs1  \u5_state_reg[8]  ( .DIN1(n9706), .CLK(clk_i),         .Q(u5_state[8]) );
  dffs1  u7_mc_ack_r_reg ( .DIN1(mc_ack_pad_i), .CLK(mc_clk_i), 
        .QN(n15513) );
  dffs1  u7_mc_br_r_reg ( .DIN1(mc_br_pad_i), .CLK(mc_clk_i),         .Q(u7_mc_br_r) );
  dffs1  \u0_u0_csc_reg[4]  ( .DIN1(n9707), .CLK(clk_i),         .QN(n31132) );
  dffs1  \u0_poc_reg[0]  ( .DIN1(n9708), .CLK(clk_i),         .Q(poc_o[0]) );
  dffs1  \u7_mc_data_ir_reg[0]  ( .DIN1(mc_data_pad_i[0]), 
        .CLK(mc_clk_i), .QN(n36637) );
  dffs1  \u0_u0_csc_reg[5]  ( .DIN1(n9709), .CLK(clk_i),         .QN(n31124) );
  dffs1  \u0_poc_reg[1]  ( .DIN1(n9710), .CLK(clk_i),         .Q(poc_o[1]) );
  dffs1  \u7_mc_data_ir_reg[1]  ( .DIN1(mc_data_pad_i[1]), 
        .CLK(mc_clk_i), .QN(n36640) );
  dffs1  u4_rfr_ce_reg ( .DIN1(n9711), .CLK(clk_i),         .Q(n36610) );
  dffs1  u4_rfr_early_reg ( .DIN1(N1549), .CLK(clk_i),         .Q(n4612) );
  dffs1  \u4_ps_cnt_reg[6]  ( .DIN1(n9712), .CLK(clk_i),         .Q(u4_ps_cnt[6]) );
  dffs1  \u4_ps_cnt_reg[5]  ( .DIN1(n9713), .CLK(clk_i),         .Q(u4_ps_cnt[5]) );
  dffs1  \u4_ps_cnt_reg[4]  ( .DIN1(n9714), .CLK(clk_i),         .Q(u4_ps_cnt[4]) );
  dffs1  \u4_ps_cnt_reg[3]  ( .DIN1(n9715), .CLK(clk_i),         .Q(u4_ps_cnt[3]) );
  dffs1  \u4_ps_cnt_reg[2]  ( .DIN1(n9716), .CLK(clk_i),         .Q(u4_ps_cnt[2]) );
  dffs1  \u4_ps_cnt_reg[1]  ( .DIN1(n9717), .CLK(clk_i),         .Q(u4_ps_cnt[1]) );
  dffs1  \u4_ps_cnt_reg[0]  ( .DIN1(n9718), .CLK(clk_i),         .Q(u4_ps_cnt[0]) );
  dffs1  \u4_ps_cnt_reg[7]  ( .DIN1(n9719), .CLK(clk_i),         .Q(u4_ps_cnt[7]) );
  dffs1  u4_rfr_en_reg ( .DIN1(n9720), .CLK(clk_i),         .QN(n4986) );
  dffs1  \u0_u0_csc_reg[1]  ( .DIN1(n9721), .CLK(clk_i),         .QN(n31119) );
  dffs1  \u0_u0_csc_reg[0]  ( .DIN1(n9722), .CLK(clk_i),         .Q(u0_csc0[0]) );
  dffs1  \u0_poc_reg[2]  ( .DIN1(n9723), .CLK(clk_i),         .Q(poc_o[2]) );
  dffs1  \u7_mc_data_ir_reg[2]  ( .DIN1(mc_data_pad_i[2]), 
        .CLK(mc_clk_i), .QN(n36643) );
  dffs1  \u0_u0_csc_reg[2]  ( .DIN1(n9724), .CLK(clk_i),         .Q(u0_csc0[2]) );
  dffs1  \u0_poc_reg[3]  ( .DIN1(n9725), .CLK(clk_i),         .Q(poc_o[3]) );
  dffs1  \u7_mc_data_ir_reg[3]  ( .DIN1(mc_data_pad_i[3]), 
        .CLK(mc_clk_i), .QN(n36646) );
  dffs1  \u0_poc_reg[4]  ( .DIN1(n9726), .CLK(clk_i),         .Q(poc_o[4]) );
  dffs1  \u7_mc_data_ir_reg[4]  ( .DIN1(mc_data_pad_i[4]), 
        .CLK(mc_clk_i), .QN(n36649) );
  dffs1  \u0_poc_reg[5]  ( .DIN1(n9727), .CLK(clk_i),         .Q(poc_o[5]) );
  dffs1  \u7_mc_data_ir_reg[5]  ( .DIN1(mc_data_pad_i[5]), 
        .CLK(mc_clk_i), .QN(n36652) );
  dffs1  \u0_poc_reg[6]  ( .DIN1(n9728), .CLK(clk_i),         .Q(poc_o[6]) );
  dffs1  \u7_mc_data_ir_reg[6]  ( .DIN1(mc_data_pad_i[6]), 
        .CLK(mc_clk_i), .QN(n36655) );
  dffs1  \u0_poc_reg[7]  ( .DIN1(n9729), .CLK(clk_i),         .Q(poc_o[7]) );
  dffs1  \u7_mc_data_ir_reg[7]  ( .DIN1(mc_data_pad_i[7]), 
        .CLK(mc_clk_i), .QN(n36658) );
  dffs1  \u0_poc_reg[8]  ( .DIN1(n9730), .CLK(clk_i),         .Q(poc_o[8]) );
  dffs1  \u7_mc_data_ir_reg[8]  ( .DIN1(mc_data_pad_i[8]), 
        .CLK(mc_clk_i), .QN(n36639) );
  dffs1  \u0_poc_reg[9]  ( .DIN1(n9731), .CLK(clk_i),         .Q(poc_o[9]) );
  dffs1  \u7_mc_data_ir_reg[9]  ( .DIN1(mc_data_pad_i[9]), 
        .CLK(mc_clk_i), .QN(n36642) );
  dffs1  \u0_poc_reg[10]  ( .DIN1(n9732), .CLK(clk_i),         .Q(poc_o[10]) );
  dffs1  \u7_mc_data_ir_reg[10]  ( .DIN1(mc_data_pad_i[10]), 
        .CLK(mc_clk_i), .QN(n36645) );
  dffs1  \u0_poc_reg[11]  ( .DIN1(n9733), .CLK(clk_i),         .Q(poc_o[11]) );
  dffs1  \u7_mc_data_ir_reg[11]  ( .DIN1(mc_data_pad_i[11]), 
        .CLK(mc_clk_i), .QN(n36648) );
  dffs1  \u0_poc_reg[12]  ( .DIN1(n9734), .CLK(clk_i),         .Q(poc_o[12]) );
  dffs1  \u7_mc_data_ir_reg[12]  ( .DIN1(mc_data_pad_i[12]), 
        .CLK(mc_clk_i), .QN(n36651) );
  dffs1  \u0_poc_reg[13]  ( .DIN1(n9735), .CLK(clk_i),         .Q(poc_o[13]) );
  dffs1  \u7_mc_data_ir_reg[13]  ( .DIN1(mc_data_pad_i[13]), 
        .CLK(mc_clk_i), .QN(n36654) );
  dffs1  \u0_poc_reg[14]  ( .DIN1(n9736), .CLK(clk_i),         .Q(poc_o[14]) );
  dffs1  \u7_mc_data_ir_reg[14]  ( .DIN1(mc_data_pad_i[14]), 
        .CLK(mc_clk_i), .QN(n36657) );
  dffs1  \u0_poc_reg[15]  ( .DIN1(n9737), .CLK(clk_i),         .Q(poc_o[15]) );
  dffs1  \u7_mc_data_ir_reg[15]  ( .DIN1(mc_data_pad_i[15]), 
        .CLK(mc_clk_i), .QN(n36660) );
  dffs1  \u0_poc_reg[16]  ( .DIN1(n9738), .CLK(clk_i),         .Q(poc_o[16]) );
  dffs1  \u7_mc_data_ir_reg[16]  ( .DIN1(mc_data_pad_i[16]), 
        .CLK(mc_clk_i), .QN(n36620) );
  dffs1  \u0_poc_reg[17]  ( .DIN1(n9739), .CLK(clk_i),         .Q(poc_o[17]) );
  dffs1  \u7_mc_data_ir_reg[17]  ( .DIN1(mc_data_pad_i[17]), 
        .CLK(mc_clk_i), .QN(n36622) );
  dffs1  \u0_poc_reg[18]  ( .DIN1(n9740), .CLK(clk_i),         .Q(poc_o[18]) );
  dffs1  \u7_mc_data_ir_reg[18]  ( .DIN1(mc_data_pad_i[18]), 
        .CLK(mc_clk_i), .QN(n36624) );
  dffs1  \u0_poc_reg[19]  ( .DIN1(n9741), .CLK(clk_i),         .Q(poc_o[19]) );
  dffs1  \u7_mc_data_ir_reg[19]  ( .DIN1(mc_data_pad_i[19]), 
        .CLK(mc_clk_i), .QN(n36626) );
  dffs1  \u0_poc_reg[20]  ( .DIN1(n9742), .CLK(clk_i),         .Q(poc_o[20]) );
  dffs1  \u7_mc_data_ir_reg[20]  ( .DIN1(mc_data_pad_i[20]), 
        .CLK(mc_clk_i), .QN(n36628) );
  dffs1  \u0_poc_reg[21]  ( .DIN1(n9743), .CLK(clk_i),         .Q(poc_o[21]) );
  dffs1  \u7_mc_data_ir_reg[21]  ( .DIN1(mc_data_pad_i[21]), 
        .CLK(mc_clk_i), .QN(n36630) );
  dffs1  \u0_poc_reg[22]  ( .DIN1(n9744), .CLK(clk_i),         .Q(poc_o[22]) );
  dffs1  \u7_mc_data_ir_reg[22]  ( .DIN1(mc_data_pad_i[22]), 
        .CLK(mc_clk_i), .QN(n36632) );
  dffs1  \u0_poc_reg[23]  ( .DIN1(n9745), .CLK(clk_i),         .Q(poc_o[23]) );
  dffs1  \u7_mc_data_ir_reg[23]  ( .DIN1(mc_data_pad_i[23]), 
        .CLK(mc_clk_i), .QN(n36634) );
  dffs1  \u0_poc_reg[24]  ( .DIN1(n9746), .CLK(clk_i),         .Q(poc_o[24]) );
  dffs1  \u7_mc_data_ir_reg[24]  ( .DIN1(mc_data_pad_i[24]), 
        .CLK(mc_clk_i), .QN(n36605) );
  dffs1  \u0_poc_reg[25]  ( .DIN1(n9747), .CLK(clk_i),         .Q(poc_o[25]) );
  dffs1  \u7_mc_data_ir_reg[25]  ( .DIN1(mc_data_pad_i[25]), 
        .CLK(mc_clk_i), .QN(n36604) );
  dffs1  \u0_poc_reg[26]  ( .DIN1(n9748), .CLK(clk_i),         .Q(poc_o[26]) );
  dffs1  \u7_mc_data_ir_reg[26]  ( .DIN1(mc_data_pad_i[26]), 
        .CLK(mc_clk_i), .QN(n36603) );
  dffs1  \u0_poc_reg[27]  ( .DIN1(n9749), .CLK(clk_i),         .Q(poc_o[27]) );
  dffs1  \u7_mc_data_ir_reg[27]  ( .DIN1(mc_data_pad_i[27]), 
        .CLK(mc_clk_i), .QN(n36602) );
  dffs1  \u0_poc_reg[28]  ( .DIN1(n9750), .CLK(clk_i),         .Q(poc_o[28]) );
  dffs1  \u7_mc_data_ir_reg[28]  ( .DIN1(mc_data_pad_i[28]), 
        .CLK(mc_clk_i), .QN(n36601) );
  dffs1  \u0_poc_reg[29]  ( .DIN1(n9751), .CLK(clk_i),         .Q(poc_o[29]) );
  dffs1  \u7_mc_data_ir_reg[29]  ( .DIN1(mc_data_pad_i[29]), 
        .CLK(mc_clk_i), .QN(n36600) );
  dffs1  \u0_poc_reg[30]  ( .DIN1(n9752), .CLK(clk_i),         .Q(poc_o[30]) );
  dffs1  \u7_mc_data_ir_reg[30]  ( .DIN1(mc_data_pad_i[30]), 
        .CLK(mc_clk_i), .QN(n36599) );
  dffs1  \u0_poc_reg[31]  ( .DIN1(n9753), .CLK(clk_i),         .Q(poc_o[31]) );
  dffs1  \u7_mc_data_ir_reg[31]  ( .DIN1(mc_data_pad_i[31]), 
        .CLK(mc_clk_i), .QN(n36598) );
  dffs1  \u0_csr_r_reg[0]  ( .DIN1(n9754), .CLK(clk_i),         .QN(n31128) );
  dffs1  u7_mc_sts_ir_reg ( .DIN1(mc_sts_pad_i), .CLK(mc_clk_i), 
        .Q(n4814) );
  dffs1  u6_read_go_r_reg ( .DIN1(n19404), .CLK(clk_i),         .QN(n15473) );
  dffs1  u6_read_go_r1_reg ( .DIN1(n9755), .CLK(clk_i),         .QN(n36597) );
  dffs1  u6_rmw_r_reg ( .DIN1(n9756), .CLK(clk_i),         .QN(n15475) );
  dffs1  u6_rmw_en_reg ( .DIN1(n9757), .CLK(clk_i),         .QN(n15471) );
  dffs1  u6_wb_ack_o_reg ( .DIN1(n9758), .CLK(clk_i),         .Q(wb_ack_o) );
  dffs1  u6_wr_hold_reg ( .DIN1(n9759), .CLK(clk_i),         .QN(n15514) );
  dffs1  u6_write_go_r1_reg ( .DIN1(n9760), .CLK(clk_i),         .Q(n4820) );
  dffs1  u6_write_go_r_reg ( .DIN1(n9761), .CLK(clk_i),         .QN(n15472) );
  dffs1  u5_wb_write_go_r_reg ( .DIN1(1'b0), .CLK(clk_i),         .Q(u5_wb_write_go_r) );
  dffs1  u5_resume_req_r_reg ( .DIN1(resume_req_i), .CLK(clk_i), .Q(u5_resume_req_r) );
  dffs1  u5_susp_req_r_reg ( .DIN1(susp_req_i), .CLK(clk_i),         .QN(n15515) );
  dffs1  u5_no_wb_cycle_reg ( .DIN1(1'b1), .CLK(clk_i),         .Q(n36596) );
  dffs1  u5_wb_cycle_reg ( .DIN1(n9762), .CLK(clk_i),         .Q(u5_wb_cycle) );
  dffs1  u5_wb_wait_r_reg ( .DIN1(n9763), .CLK(clk_i),         .Q(u5_wb_wait_r) );
  dffs1  u5_wb_wait_r2_reg ( .DIN1(1'b0), .CLK(clk_i),         .Q(n9763) );
  dffs1  u5_mem_ack_r_reg ( .DIN1(1'b0), .CLK(clk_i),         .Q(u5_mem_ack_r) );
  dffs1  u5_mc_le_reg ( .DIN1(n9764), .CLK(clk_i), .QN(n9764) );
  dffs1  u5_rsts_reg ( .DIN1(n9765), .CLK(clk_i), .Q(u5_rsts)
         );
  dffs1  u5_rsts1_reg ( .DIN1(1'b0), .CLK(mc_clk_i),         .Q(n9765) );
  dffs1  \u3_u0_rd_adr_reg[0]  ( .DIN1(n9766), .CLK(clk_i),         .Q(u3_u0_rd_adr[0]) );
  dffs1  \u3_u0_rd_adr_reg[1]  ( .DIN1(n9767), .CLK(clk_i),         .Q(u3_u0_rd_adr[1]) );
  dffs1  \u3_u0_rd_adr_reg[2]  ( .DIN1(n9768), .CLK(clk_i),         .Q(u3_u0_rd_adr[2]) );
  dffs1  \u3_u0_rd_adr_reg[3]  ( .DIN1(n9769), .CLK(clk_i),         .Q(u3_u0_rd_adr[3]) );
  dffs1  \u1_sram_addr_reg[0]  ( .DIN1(n9770), .CLK(clk_i),         .QN(n36710) );
  dffs1  \u1_sram_addr_reg[1]  ( .DIN1(n9771), .CLK(clk_i),         .QN(n36707) );
  dffs1  \u1_sram_addr_reg[2]  ( .DIN1(n9772), .CLK(clk_i),         .QN(n36704) );
  dffs1  \u1_sram_addr_reg[3]  ( .DIN1(n9773), .CLK(clk_i),         .QN(n36701) );
  dffs1  \u1_sram_addr_reg[4]  ( .DIN1(n9774), .CLK(clk_i),         .QN(n36698) );
  dffs1  \u1_sram_addr_reg[5]  ( .DIN1(n9775), .CLK(clk_i),         .QN(n36695) );
  dffs1  \u1_sram_addr_reg[6]  ( .DIN1(n9776), .CLK(clk_i),         .QN(n36692) );
  dffs1  \u1_sram_addr_reg[7]  ( .DIN1(n9777), .CLK(clk_i),         .QN(n36689) );
  dffs1  \u1_sram_addr_reg[8]  ( .DIN1(n9778), .CLK(clk_i),         .QN(n36686) );
  dffs1  \u1_sram_addr_reg[9]  ( .DIN1(n9779), .CLK(clk_i),         .QN(n36683) );
  dffs1  \u1_sram_addr_reg[10]  ( .DIN1(n9780), .CLK(clk_i),         .QN(n36681) );
  dffs1  \u1_sram_addr_reg[11]  ( .DIN1(n9781), .CLK(clk_i),         .QN(n36679) );
  dffs1  \u1_sram_addr_reg[12]  ( .DIN1(n9782), .CLK(clk_i),         .QN(n36677) );
  dffs1  \u1_sram_addr_reg[13]  ( .DIN1(n9783), .CLK(clk_i),         .QN(n36676) );
  dffs1  \u1_sram_addr_reg[14]  ( .DIN1(n9784), .CLK(clk_i),         .QN(n36674) );
  dffs1  \u1_sram_addr_reg[15]  ( .DIN1(n9785), .CLK(clk_i),         .QN(n36672) );
  dffs1  \u1_sram_addr_reg[16]  ( .DIN1(n9786), .CLK(clk_i),         .QN(n36671) );
  dffs1  \u1_sram_addr_reg[17]  ( .DIN1(n9787), .CLK(clk_i),         .QN(n36670) );
  dffs1  \u1_sram_addr_reg[18]  ( .DIN1(n9788), .CLK(clk_i),         .QN(n36669) );
  dffs1  \u1_sram_addr_reg[19]  ( .DIN1(n9789), .CLK(clk_i),         .QN(n36668) );
  dffs1  \u1_sram_addr_reg[20]  ( .DIN1(n9790), .CLK(clk_i),         .QN(n36667) );
  dffs1  \u1_sram_addr_reg[21]  ( .DIN1(n9791), .CLK(clk_i),         .QN(n36666) );
  dffs1  \u1_sram_addr_reg[22]  ( .DIN1(n9792), .CLK(clk_i),         .QN(n36665) );
  dffs1  \u1_sram_addr_reg[23]  ( .DIN1(n9793), .CLK(clk_i),         .QN(n36663) );
  dffs1  u0_u1_init_req_we_reg ( .DIN1(n9794), .CLK(clk_i),         .Q(n4618) );
  dffs1  u0_u1_lmr_req_we_reg ( .DIN1(n9795), .CLK(clk_i),         .QN(n4991) );
  dffs1  \u0_u1_tms_reg[0]  ( .DIN1(n9796), .CLK(clk_i),         .QN(n31129) );
  dffs1  \u0_u1_tms_reg[1]  ( .DIN1(n9797), .CLK(clk_i),         .QN(n31121) );
  dffs1  \u0_u1_tms_reg[2]  ( .DIN1(n9798), .CLK(clk_i),         .QN(n31116) );
  dffs1  \u0_u1_tms_reg[3]  ( .DIN1(n9799), .CLK(clk_i),         .QN(n31114) );
  dffs1  \u0_u1_tms_reg[4]  ( .DIN1(n9800), .CLK(clk_i),         .QN(n31134) );
  dffs1  \u0_u1_tms_reg[5]  ( .DIN1(n9801), .CLK(clk_i),         .QN(n31126) );
  dffs1  \u0_u1_tms_reg[6]  ( .DIN1(n9802), .CLK(clk_i),         .QN(n31111) );
  dffs1  \u0_u1_tms_reg[7]  ( .DIN1(n9803), .CLK(clk_i),         .QN(n31106) );
  dffs1  \u0_u1_tms_reg[8]  ( .DIN1(n9804), .CLK(clk_i),         .QN(n31100) );
  dffs1  \u0_u1_tms_reg[9]  ( .DIN1(n9805), .CLK(clk_i),         .QN(n31097) );
  dffs1  \u0_u1_tms_reg[10]  ( .DIN1(n9806), .CLK(clk_i),         .QN(n31092) );
  dffs1  \u0_u1_tms_reg[11]  ( .DIN1(n9807), .CLK(clk_i),         .QN(n31088) );
  dffs1  \u0_u1_tms_reg[12]  ( .DIN1(n9808), .CLK(clk_i),         .QN(n31084) );
  dffs1  \u0_u1_tms_reg[13]  ( .DIN1(n9809), .CLK(clk_i),         .QN(n31080) );
  dffs1  \u0_u1_tms_reg[14]  ( .DIN1(n9810), .CLK(clk_i),         .QN(n31076) );
  dffs1  \u0_u1_tms_reg[15]  ( .DIN1(n9811), .CLK(clk_i),         .QN(n31072) );
  dffs1  \u0_u1_tms_reg[16]  ( .DIN1(n9812), .CLK(clk_i),         .QN(n31068) );
  dffs1  \u0_u1_tms_reg[17]  ( .DIN1(n9813), .CLK(clk_i),         .QN(n31066) );
  dffs1  \u0_u1_tms_reg[18]  ( .DIN1(n9814), .CLK(clk_i),         .QN(n31064) );
  dffs1  \u0_u1_tms_reg[19]  ( .DIN1(n9815), .CLK(clk_i),         .QN(n31062) );
  dffs1  \u0_u1_tms_reg[20]  ( .DIN1(n9816), .CLK(clk_i),         .QN(n31060) );
  dffs1  \u0_u1_tms_reg[21]  ( .DIN1(n9817), .CLK(clk_i),         .QN(n31058) );
  dffs1  \u0_u1_tms_reg[22]  ( .DIN1(n9818), .CLK(clk_i),         .QN(n31056) );
  dffs1  \u0_u1_tms_reg[23]  ( .DIN1(n9819), .CLK(clk_i),         .QN(n31054) );
  dffs1  \u0_u1_tms_reg[24]  ( .DIN1(n9820), .CLK(clk_i),         .QN(n31052) );
  dffs1  \u0_u1_tms_reg[25]  ( .DIN1(n9821), .CLK(clk_i),         .QN(n31048) );
  dffs1  \u0_u1_tms_reg[26]  ( .DIN1(n9822), .CLK(clk_i),         .QN(n31044) );
  dffs1  \u0_u1_tms_reg[27]  ( .DIN1(n9823), .CLK(clk_i),         .QN(n31040) );
  dffs1  \u0_u1_tms_reg[28]  ( .DIN1(n9824), .CLK(clk_i),         .QN(n31036) );
  dffs1  \u0_u1_tms_reg[29]  ( .DIN1(n9825), .CLK(clk_i),         .QN(n31032) );
  dffs1  \u0_u1_tms_reg[30]  ( .DIN1(n9826), .CLK(clk_i),         .QN(n31028) );
  dffs1  \u0_u1_tms_reg[31]  ( .DIN1(n9827), .CLK(clk_i),         .QN(n31024) );
  dffs1  \u0_u1_csc_reg[0]  ( .DIN1(n9828), .CLK(clk_i),         .Q(u0_csc1[0]) );
  dffs1  \u0_u1_csc_reg[1]  ( .DIN1(n9829), .CLK(clk_i),         .QN(n31120) );
  dffs1  \u0_u1_csc_reg[2]  ( .DIN1(n9830), .CLK(clk_i),         .Q(u0_csc1[2]) );
  dffs1  \u0_u1_csc_reg[3]  ( .DIN1(n9831), .CLK(clk_i),         .Q(u0_csc1[3]) );
  dffs1  \u0_u1_csc_reg[4]  ( .DIN1(n9832), .CLK(clk_i),         .QN(n31133) );
  dffs1  \u0_u1_csc_reg[5]  ( .DIN1(n9833), .CLK(clk_i),         .QN(n31125) );
  dffs1  \u0_u1_csc_reg[6]  ( .DIN1(n9834), .CLK(clk_i),         .QN(n31110) );
  dffs1  \u0_u1_csc_reg[7]  ( .DIN1(n9835), .CLK(clk_i),         .QN(n31105) );
  dffs1  \u0_u1_csc_reg[8]  ( .DIN1(n9836), .CLK(clk_i),         .Q(u0_csc1[8]) );
  dffs1  \u0_u1_csc_reg[9]  ( .DIN1(n9837), .CLK(clk_i),         .QN(n31096) );
  dffs1  \u0_u1_csc_reg[10]  ( .DIN1(n9838), .CLK(clk_i),         .QN(n31091) );
  dffs1  \u0_u1_csc_reg[11]  ( .DIN1(n9839), .CLK(clk_i),         .QN(n31087) );
  dffs1  \u0_u1_csc_reg[12]  ( .DIN1(n9840), .CLK(clk_i),         .QN(n31083) );
  dffs1  \u0_u1_csc_reg[13]  ( .DIN1(n9841), .CLK(clk_i),         .QN(n31079) );
  dffs1  \u0_u1_csc_reg[14]  ( .DIN1(n9842), .CLK(clk_i),         .QN(n31075) );
  dffs1  \u0_u1_csc_reg[15]  ( .DIN1(n9843), .CLK(clk_i),         .QN(n31071) );
  dffs1  \u0_u1_csc_reg[16]  ( .DIN1(n9844), .CLK(clk_i),         .Q(u0_csc1[16]) );
  dffs1  \u0_u1_csc_reg[17]  ( .DIN1(n9845), .CLK(clk_i),         .Q(u0_csc1[17]) );
  dffs1  \u0_u1_csc_reg[18]  ( .DIN1(n9846), .CLK(clk_i),         .Q(u0_csc1[18]) );
  dffs1  \u0_u1_csc_reg[19]  ( .DIN1(n9847), .CLK(clk_i),         .Q(u0_csc1[19]) );
  dffs1  \u0_u1_csc_reg[20]  ( .DIN1(n9848), .CLK(clk_i),         .Q(u0_csc1[20]) );
  dffs1  \u0_u1_csc_reg[21]  ( .DIN1(n9849), .CLK(clk_i),         .Q(u0_csc1[21]) );
  dffs1  \u0_u1_csc_reg[22]  ( .DIN1(n9850), .CLK(clk_i),         .Q(u0_csc1[22]) );
  dffs1  \u0_u1_csc_reg[23]  ( .DIN1(n9851), .CLK(clk_i),         .Q(u0_csc1[23]) );
  dffs1  \u0_u1_csc_reg[24]  ( .DIN1(n9852), .CLK(clk_i),         .QN(n31051) );
  dffs1  \u0_u1_csc_reg[25]  ( .DIN1(n9853), .CLK(clk_i),         .QN(n31047) );
  dffs1  \u0_u1_csc_reg[26]  ( .DIN1(n9854), .CLK(clk_i),         .QN(n31043) );
  dffs1  \u0_u1_csc_reg[27]  ( .DIN1(n9855), .CLK(clk_i),         .QN(n31039) );
  dffs1  \u0_u1_csc_reg[28]  ( .DIN1(n9856), .CLK(clk_i),         .QN(n31035) );
  dffs1  \u0_u1_csc_reg[29]  ( .DIN1(n9857), .CLK(clk_i),         .QN(n31031) );
  dffs1  \u0_u1_csc_reg[30]  ( .DIN1(n9858), .CLK(clk_i),         .QN(n31027) );
  dffs1  \u0_u1_csc_reg[31]  ( .DIN1(n9859), .CLK(clk_i),         .QN(n31023) );
  dffs1  \u0_u1_addr_r_reg[2]  ( .DIN1(wb_addr_i[2]), .CLK(clk_i), .QN(n15486) );
  dffs1  \u0_u1_addr_r_reg[3]  ( .DIN1(wb_addr_i[3]), .CLK(clk_i), .Q(n36589) );
  dffs1  \u0_u1_addr_r_reg[4]  ( .DIN1(wb_addr_i[4]), .CLK(clk_i), .Q(n36588) );
  dffs1  \u0_u1_addr_r_reg[5]  ( .DIN1(wb_addr_i[5]), .CLK(clk_i), .QN(n36586) );
  dffs1  \u0_u1_addr_r_reg[6]  ( .DIN1(wb_addr_i[6]), .CLK(clk_i), .QN(n36587) );
  dffs1  u0_u1_rst_r2_reg ( .DIN1(n9860), .CLK(clk_i),         .Q(n36585) );
  dffs1  u0_u1_rst_r1_reg ( .DIN1(1'b0), .CLK(clk_i),         .Q(n9860) );
  dffs1  u0_u0_init_req_we_reg ( .DIN1(n19405), .CLK(clk_i),         .Q(n4616) );
  dffs1  u0_u0_lmr_req_we_reg ( .DIN1(n19406), .CLK(clk_i),         .QN(n4992) );
  dffs1  \u0_u0_tms_reg[0]  ( .DIN1(n9863), .CLK(clk_i),         .QN(n31127) );
  dffs1  \u0_u0_tms_reg[1]  ( .DIN1(n9864), .CLK(clk_i),         .QN(n31117) );
  dffs1  \u0_u0_tms_reg[2]  ( .DIN1(n9865), .CLK(clk_i),         .QN(n31115) );
  dffs1  \u0_u0_tms_reg[3]  ( .DIN1(n9866), .CLK(clk_i),         .QN(n31112) );
  dffs1  \u0_u0_tms_reg[4]  ( .DIN1(n9867), .CLK(clk_i),         .QN(n31130) );
  dffs1  \u0_u0_tms_reg[5]  ( .DIN1(n9868), .CLK(clk_i),         .QN(n31122) );
  dffs1  \u0_u0_tms_reg[6]  ( .DIN1(n9869), .CLK(clk_i),         .QN(n31107) );
  dffs1  \u0_u0_tms_reg[7]  ( .DIN1(n9870), .CLK(clk_i),         .QN(n31102) );
  dffs1  \u0_u0_tms_reg[8]  ( .DIN1(n9871), .CLK(clk_i),         .QN(n31099) );
  dffs1  \u0_u0_tms_reg[9]  ( .DIN1(n9872), .CLK(clk_i),         .QN(n31094) );
  dffs1  \u0_u0_tms_reg[10]  ( .DIN1(n9873), .CLK(clk_i),         .QN(n31089) );
  dffs1  \u0_u0_tms_reg[11]  ( .DIN1(n9874), .CLK(clk_i),         .QN(n31086) );
  dffs1  \u0_u0_tms_reg[12]  ( .DIN1(n9875), .CLK(clk_i),         .QN(n31082) );
  dffs1  \u0_u0_tms_reg[13]  ( .DIN1(n9876), .CLK(clk_i),         .QN(n31078) );
  dffs1  \u0_u0_tms_reg[14]  ( .DIN1(n9877), .CLK(clk_i),         .QN(n31074) );
  dffs1  \u0_u0_tms_reg[15]  ( .DIN1(n9878), .CLK(clk_i),         .QN(n31070) );
  dffs1  \u0_u0_tms_reg[16]  ( .DIN1(n9879), .CLK(clk_i),         .QN(n31067) );
  dffs1  \u0_u0_tms_reg[17]  ( .DIN1(n9880), .CLK(clk_i),         .QN(n31065) );
  dffs1  \u0_u0_tms_reg[18]  ( .DIN1(n9881), .CLK(clk_i),         .QN(n31063) );
  dffs1  \u0_u0_tms_reg[19]  ( .DIN1(n9882), .CLK(clk_i),         .QN(n31061) );
  dffs1  \u0_u0_tms_reg[20]  ( .DIN1(n9883), .CLK(clk_i),         .QN(n31059) );
  dffs1  \u0_u0_tms_reg[21]  ( .DIN1(n9884), .CLK(clk_i),         .QN(n31057) );
  dffs1  \u0_u0_tms_reg[22]  ( .DIN1(n9885), .CLK(clk_i),         .QN(n31055) );
  dffs1  \u0_u0_tms_reg[23]  ( .DIN1(n9886), .CLK(clk_i),         .QN(n31053) );
  dffs1  \u0_u0_tms_reg[24]  ( .DIN1(n9887), .CLK(clk_i),         .QN(n31049) );
  dffs1  \u0_u0_tms_reg[25]  ( .DIN1(n9888), .CLK(clk_i),         .QN(n31045) );
  dffs1  \u0_u0_tms_reg[26]  ( .DIN1(n9889), .CLK(clk_i),         .QN(n31041) );
  dffs1  \u0_u0_tms_reg[27]  ( .DIN1(n9890), .CLK(clk_i),         .QN(n31037) );
  dffs1  \u0_u0_tms_reg[28]  ( .DIN1(n9891), .CLK(clk_i),         .QN(n31033) );
  dffs1  \u0_u0_tms_reg[29]  ( .DIN1(n9892), .CLK(clk_i),         .QN(n31029) );
  dffs1  \u0_u0_tms_reg[30]  ( .DIN1(n9893), .CLK(clk_i),         .QN(n31025) );
  dffs1  \u0_u0_tms_reg[31]  ( .DIN1(n9894), .CLK(clk_i),         .QN(n31021) );
  dffs1  \u0_u0_csc_reg[3]  ( .DIN1(n9895), .CLK(clk_i),         .Q(u0_csc0[3]) );
  dffs1  \u0_u0_csc_reg[6]  ( .DIN1(n9896), .CLK(clk_i),         .QN(n31109) );
  dffs1  \u0_u0_csc_reg[7]  ( .DIN1(n9897), .CLK(clk_i),         .QN(n31104) );
  dffs1  \u0_u0_csc_reg[8]  ( .DIN1(n9898), .CLK(clk_i),         .Q(u0_csc0[8]) );
  dffs1  \u0_u0_csc_reg[9]  ( .DIN1(n9899), .CLK(clk_i),         .QN(n31095) );
  dffs1  \u0_u0_csc_reg[10]  ( .DIN1(n9900), .CLK(clk_i),         .QN(n31090) );
  dffs1  \u0_u0_csc_reg[11]  ( .DIN1(n9901), .CLK(clk_i),         .QN(n31085) );
  dffs1  \u0_u0_csc_reg[12]  ( .DIN1(n9902), .CLK(clk_i),         .QN(n31081) );
  dffs1  \u0_u0_csc_reg[13]  ( .DIN1(n9903), .CLK(clk_i),         .QN(n31077) );
  dffs1  \u0_u0_csc_reg[14]  ( .DIN1(n9904), .CLK(clk_i),         .QN(n31073) );
  dffs1  \u0_u0_csc_reg[15]  ( .DIN1(n9905), .CLK(clk_i),         .QN(n31069) );
  dffs1  \u0_u0_csc_reg[16]  ( .DIN1(n9906), .CLK(clk_i),         .Q(u0_csc0[16]) );
  dffs1  \u0_u0_csc_reg[17]  ( .DIN1(n9907), .CLK(clk_i),         .Q(u0_csc0[17]) );
  dffs1  \u0_u0_csc_reg[18]  ( .DIN1(n9908), .CLK(clk_i),         .Q(u0_csc0[18]) );
  dffs1  \u0_u0_csc_reg[19]  ( .DIN1(n9909), .CLK(clk_i),         .Q(u0_csc0[19]) );
  dffs1  \u0_u0_csc_reg[20]  ( .DIN1(n9910), .CLK(clk_i),         .Q(u0_csc0[20]) );
  dffs1  \u0_u0_csc_reg[21]  ( .DIN1(n9911), .CLK(clk_i),         .Q(u0_csc0[21]) );
  dffs1  \u0_u0_csc_reg[22]  ( .DIN1(n9912), .CLK(clk_i),         .Q(u0_csc0[22]) );
  dffs1  \u0_u0_csc_reg[23]  ( .DIN1(n9913), .CLK(clk_i),         .Q(u0_csc0[23]) );
  dffs1  \u0_u0_csc_reg[24]  ( .DIN1(n9914), .CLK(clk_i),         .QN(n31050) );
  dffs1  \u0_u0_csc_reg[25]  ( .DIN1(n9915), .CLK(clk_i),         .QN(n31046) );
  dffs1  \u0_u0_csc_reg[26]  ( .DIN1(n9916), .CLK(clk_i),         .QN(n31042) );
  dffs1  \u0_u0_csc_reg[27]  ( .DIN1(n9917), .CLK(clk_i),         .QN(n31038) );
  dffs1  \u0_u0_csc_reg[28]  ( .DIN1(n9918), .CLK(clk_i),         .QN(n31034) );
  dffs1  \u0_u0_csc_reg[29]  ( .DIN1(n9919), .CLK(clk_i),         .QN(n31030) );
  dffs1  \u0_u0_csc_reg[30]  ( .DIN1(n9920), .CLK(clk_i),         .QN(n31026) );
  dffs1  \u0_u0_csc_reg[31]  ( .DIN1(n9921), .CLK(clk_i),         .QN(n31022) );
  dffs1  \u0_u0_addr_r_reg[2]  ( .DIN1(wb_addr_i[2]), .CLK(clk_i), .Q(n36590) );
  dffs1  \u0_u0_addr_r_reg[3]  ( .DIN1(wb_addr_i[3]), .CLK(clk_i), .QN(n36591) );
  dffs1  \u0_u0_addr_r_reg[4]  ( .DIN1(wb_addr_i[4]), .CLK(clk_i), .Q(n36594) );
  dffs1  \u0_u0_addr_r_reg[5]  ( .DIN1(wb_addr_i[5]), .CLK(clk_i), .QN(n36592) );
  dffs1  \u0_u0_addr_r_reg[6]  ( .DIN1(wb_addr_i[6]), .CLK(clk_i), .QN(n36593) );
  dffs1  u0_u0_rst_r2_reg ( .DIN1(n9922), .CLK(clk_i),         .QN(n15487) );
  dffs1  u0_u0_rst_r1_reg ( .DIN1(1'b0), .CLK(clk_i),         .Q(n9922) );
  dffs1  u0_rst_r3_reg ( .DIN1(n9923), .CLK(clk_i),         .QN(n15521) );
  dffs1  u0_rst_r2_reg ( .DIN1(n9924), .CLK(clk_i),         .Q(n9923) );
  dffs1  u0_rst_r1_reg ( .DIN1(1'b0), .CLK(clk_i),         .Q(n9924) );
  dffs1  \u0_csc_mask_r_reg[0]  ( .DIN1(n9925), .CLK(clk_i),         .Q(u0_csc_mask_r[0]) );
  dffs1  \u0_csc_mask_r_reg[1]  ( .DIN1(n9926), .CLK(clk_i),         .Q(u0_csc_mask_r[1]) );
  dffs1  \u0_csc_mask_r_reg[2]  ( .DIN1(n9927), .CLK(clk_i),         .Q(u0_csc_mask_r[2]) );
  dffs1  \u0_csc_mask_r_reg[3]  ( .DIN1(n9928), .CLK(clk_i),         .Q(u0_csc_mask_r[3]) );
  dffs1  \u0_csc_mask_r_reg[4]  ( .DIN1(n9929), .CLK(clk_i),         .Q(u0_csc_mask_r[4]) );
  dffs1  \u0_csc_mask_r_reg[5]  ( .DIN1(n9930), .CLK(clk_i),         .Q(u0_csc_mask_r[5]) );
  dffs1  \u0_csc_mask_r_reg[6]  ( .DIN1(n9931), .CLK(clk_i),         .Q(u0_csc_mask_r[6]) );
  dffs1  \u0_csc_mask_r_reg[7]  ( .DIN1(n9932), .CLK(clk_i),         .Q(u0_csc_mask_r[7]) );
  dffs1  \u0_csc_mask_r_reg[8]  ( .DIN1(n9933), .CLK(clk_i),         .QN(n31101) );
  dffs1  \u0_csc_mask_r_reg[9]  ( .DIN1(n9934), .CLK(clk_i),         .QN(n31098) );
  dffs1  \u0_csc_mask_r_reg[10]  ( .DIN1(n9935), .CLK(clk_i),         .QN(n31093) );
  dffs1  u0_trig_reg ( .DIN1(n9936), .CLK(clk_i), .QN(n15488)
         );
  dffs1  \u0_csr_r_reg[1]  ( .DIN1(n9937), .CLK(clk_i),         .Q(mc_vpen_pad_o), .QN(n31118) );
  dffs1  \u0_csr_r_reg[2]  ( .DIN1(n9938), .CLK(clk_i),         .QN(n15523) );
  dffs1  \u0_csr_r_reg[3]  ( .DIN1(n9939), .CLK(clk_i),         .QN(n31113) );
  dffs1  \u0_csr_r_reg[4]  ( .DIN1(n9940), .CLK(clk_i),         .QN(n31131) );
  dffs1  \u0_csr_r_reg[5]  ( .DIN1(n9941), .CLK(clk_i),         .QN(n31123) );
  dffs1  \u0_csr_r_reg[6]  ( .DIN1(n9942), .CLK(clk_i),         .QN(n31108) );
  dffs1  \u0_csr_r_reg[7]  ( .DIN1(n9943), .CLK(clk_i),         .QN(n31103) );
  dffs1  \u0_csr_r_reg[8]  ( .DIN1(n9944), .CLK(clk_i),         .Q(u0_csr_r[8]) );
  dffs1  \u0_csr_r_reg[9]  ( .DIN1(n9945), .CLK(clk_i),         .Q(u0_csr_r[9]) );
  dffs1  \u0_csr_r_reg[10]  ( .DIN1(n9946), .CLK(clk_i),         .Q(u0_csr_r[10]) );
  dffs1  \u0_csr_tj_val_reg[0]  ( .DIN1(n9947), .CLK(clk_i),         .QN(n36584) );
  dffs1  \u0_csr_tj_val_reg[1]  ( .DIN1(n9948), .CLK(clk_i),         .QN(n36583) );
  dffs1  \u0_csr_tj_val_reg[2]  ( .DIN1(n9949), .CLK(clk_i),         .QN(n36582) );
  dffs1  \u0_csr_tj_val_reg[3]  ( .DIN1(n9950), .CLK(clk_i),         .Q(u0_csr_tj_val[3]) );
  dffs1  \u0_csr_tj_val_reg[4]  ( .DIN1(n9951), .CLK(clk_i),         .QN(n36581) );
  dffs1  \u0_csr_tj_val_reg[5]  ( .DIN1(n9952), .CLK(clk_i),         .QN(n36580) );
  dffs1  \u0_csr_tj_val_reg[6]  ( .DIN1(n9953), .CLK(clk_i),         .QN(n36579) );
  dffs1  \u0_csr_tj_val_reg[7]  ( .DIN1(n9954), .CLK(clk_i),         .Q(u0_csr_tj_val[7]) );
  dffs1  \u0_csr_r2_reg[0]  ( .DIN1(n9955), .CLK(clk_i),         .Q(u0_csr_r2[0]) );
  dffs1  \u0_csr_r2_reg[1]  ( .DIN1(n9956), .CLK(clk_i),         .Q(u0_csr_r2[1]) );
  dffs1  \u0_csr_r2_reg[2]  ( .DIN1(n9957), .CLK(clk_i),         .Q(u0_csr_r2[2]) );
  dffs1  \u0_csr_r2_reg[3]  ( .DIN1(n9958), .CLK(clk_i),         .Q(u0_csr_r2[3]) );
  dffs1  \u0_csr_r2_reg[4]  ( .DIN1(n9959), .CLK(clk_i),         .Q(u0_csr_r2[4]) );
  dffs1  \u0_csr_r2_reg[5]  ( .DIN1(n9960), .CLK(clk_i),         .Q(u0_csr_r2[5]) );
  dffs1  \u0_csr_r2_reg[6]  ( .DIN1(n9961), .CLK(clk_i),         .Q(u0_csr_r2[6]) );
  dffs1  \u0_csr_r2_reg[7]  ( .DIN1(n9962), .CLK(clk_i),         .Q(u0_csr_r2[7]) );
  dffs1  u0_rf_we_reg ( .DIN1(n9963), .CLK(clk_i),         .Q(n36609) );
  dffs1  \u0_wb_addr_r_reg[2]  ( .DIN1(wb_addr_i[2]), .CLK(clk_i), .Q(u0_wb_addr_r[2]) );
  dffs1  \u0_wb_addr_r_reg[3]  ( .DIN1(wb_addr_i[3]), .CLK(clk_i), .Q(u0_wb_addr_r[3]) );
  dffs1  \u0_wb_addr_r_reg[4]  ( .DIN1(wb_addr_i[4]), .CLK(clk_i), .Q(n4975) );
  dffs1  \u0_wb_addr_r_reg[5]  ( .DIN1(wb_addr_i[5]), .CLK(clk_i), .Q(u0_wb_addr_r[5]) );
  dffs1  \u0_wb_addr_r_reg[6]  ( .DIN1(wb_addr_i[6]), .CLK(clk_i), .Q(u0_wb_addr_r[6]) );
  dffs1  mem_ack_r_reg ( .DIN1(1'b0), .CLK(clk_i),         .Q(n15482) );
  and2s1 U23054 ( .DIN1(n15531), .DIN2(n31272), .Q(n5176) );
  or2s1 U23055 ( .DIN1(n31268), .DIN2(n15531), .Q(n31932) );
  hi1s1 U23056 ( .DIN1(n31932), .Q(n31930) );
  or2s1 U23057 ( .DIN1(n31930), .DIN2(n31266), .Q(n5175) );
  and2s1 U23058 ( .DIN1(n34100), .DIN2(n35360), .Q(n5504) );
  or2s1 U23059 ( .DIN1(n35285), .DIN2(n5504), .Q(n31264) );
  hi1s1 U23060 ( .DIN1(n31264), .Q(n5503) );
  and2s1 U23061 ( .DIN1(n15530), .DIN2(n31272), .Q(n19401) );
  or2s1 U23062 ( .DIN1(n31268), .DIN2(n15530), .Q(n31267) );
  hi1s1 U23063 ( .DIN1(n31267), .Q(n31265) );
  or2s1 U23064 ( .DIN1(n31265), .DIN2(n31266), .Q(n5499) );
  hi1s1 U23065 ( .DIN1(n35082), .Q(n35066) );
  and2s1 U23066 ( .DIN1(n34100), .DIN2(n35066), .Q(n35167) );
  or2s1 U23067 ( .DIN1(n34958), .DIN2(n32850), .Q(n35372) );
  hi1s1 U23068 ( .DIN1(n35372), .Q(n34296) );
  hi1s1 U23069 ( .DIN1(n35071), .Q(n35277) );
  hi1s1 U23070 ( .DIN1(n35069), .Q(n35276) );
  or2s1 U23071 ( .DIN1(n35276), .DIN2(n35277), .Q(n31271) );
  and2s1 U23072 ( .DIN1(n35082), .DIN2(n31271), .Q(n35360) );
  and2s1 U23073 ( .DIN1(n35360), .DIN2(n34296), .Q(n31270) );
  or2s1 U23074 ( .DIN1(n31270), .DIN2(n35167), .Q(n5496) );
  or2s1 U23075 ( .DIN1(n35285), .DIN2(n5496), .Q(n31269) );
  hi1s1 U23076 ( .DIN1(n31269), .Q(n5495) );
  and2s1 U23077 ( .DIN1(n15529), .DIN2(n31272), .Q(n5492) );
  or2s1 U23078 ( .DIN1(n31268), .DIN2(n15529), .Q(n31274) );
  hi1s1 U23079 ( .DIN1(n31274), .Q(n31273) );
  or2s1 U23080 ( .DIN1(n31273), .DIN2(n31266), .Q(n5491) );
  hi1s1 U23081 ( .DIN1(n31275), .Q(n19403) );
  hi1s1 U23082 ( .DIN1(n35141), .Q(n34958) );
  and2s1 U23083 ( .DIN1(n34958), .DIN2(n34957), .Q(n34100) );
  hi1s1 U23084 ( .DIN1(n32850), .Q(n34957) );
  or2s1 U23085 ( .DIN1(n35071), .DIN2(n35069), .Q(n35082) );
  and2s1 U23086 ( .DIN1(n35082), .DIN2(n34957), .Q(n35151) );
  or2s1 U23087 ( .DIN1(n35151), .DIN2(n34100), .Q(n35077) );
  or2s1 U23088 ( .DIN1(n35285), .DIN2(n35077), .Q(n31275) );
  and2s1 U23089 ( .DIN1(n19408), .DIN2(n31275), .Q(n5487) );
  and2s1 U23090 ( .DIN1(n15528), .DIN2(n31272), .Q(n5484) );
  or2s1 U23091 ( .DIN1(n31268), .DIN2(n15528), .Q(n31277) );
  hi1s1 U23092 ( .DIN1(n31277), .Q(n31276) );
  or2s1 U23093 ( .DIN1(n31276), .DIN2(n31266), .Q(n5483) );
  hi1s1 U23094 ( .DIN1(n31263), .Q(n34093) );
  and2s1 U23095 ( .DIN1(n35282), .DIN2(n34093), .Q(n31936) );
  and2s1 U23096 ( .DIN1(u0_csc[5]), .DIN2(n35283), .Q(n31935) );
  or2s1 U23097 ( .DIN1(n31935), .DIN2(n31936), .Q(n32850) );
  and2s1 U23098 ( .DIN1(u0_sp_csc[4]), .DIN2(n35282), .Q(n31938) );
  and2s1 U23099 ( .DIN1(u0_csc[4]), .DIN2(n35283), .Q(n31937) );
  or2s1 U23100 ( .DIN1(n31937), .DIN2(n31938), .Q(n35141) );
  and2s1 U23101 ( .DIN1(n35141), .DIN2(n32850), .Q(n31934) );
  and2s1 U23102 ( .DIN1(u0_sp_csc[6]), .DIN2(n35282), .Q(n31940) );
  and2s1 U23103 ( .DIN1(u0_csc[6]), .DIN2(n35283), .Q(n31939) );
  or2s1 U23104 ( .DIN1(n31939), .DIN2(n31940), .Q(n35069) );
  and2s1 U23105 ( .DIN1(u0_sp_csc[7]), .DIN2(n35282), .Q(n31942) );
  and2s1 U23106 ( .DIN1(u0_csc[7]), .DIN2(n35283), .Q(n31941) );
  or2s1 U23107 ( .DIN1(n31941), .DIN2(n31942), .Q(n35071) );
  and2s1 U23108 ( .DIN1(n35071), .DIN2(n35069), .Q(n35371) );
  or2s1 U23109 ( .DIN1(n35371), .DIN2(n31934), .Q(n35285) );
  hi1s1 U23110 ( .DIN1(n35285), .Q(n19408) );
  and2s1 U23111 ( .DIN1(n15527), .DIN2(n31272), .Q(n5477) );
  or2s1 U23112 ( .DIN1(n31268), .DIN2(n15527), .Q(n31279) );
  hi1s1 U23113 ( .DIN1(n31279), .Q(n31278) );
  or2s1 U23114 ( .DIN1(n31278), .DIN2(n31266), .Q(n5476) );
  and2s1 U23115 ( .DIN1(n15526), .DIN2(n31272), .Q(n5471) );
  or2s1 U23116 ( .DIN1(n31268), .DIN2(n15526), .Q(n31281) );
  hi1s1 U23117 ( .DIN1(n31281), .Q(n31280) );
  or2s1 U23118 ( .DIN1(n31280), .DIN2(n31266), .Q(n5470) );
  and2s1 U23119 ( .DIN1(n15525), .DIN2(n31272), .Q(n5465) );
  hi1s1 U23120 ( .DIN1(n31272), .Q(n31931) );
  and2s1 U23121 ( .DIN1(n31285), .DIN2(n31931), .Q(n31266) );
  or2s1 U23122 ( .DIN1(n31268), .DIN2(n15525), .Q(n31283) );
  hi1s1 U23123 ( .DIN1(n31283), .Q(n31282) );
  or2s1 U23124 ( .DIN1(n31282), .DIN2(n31266), .Q(n5464) );
  hi1s1 U23125 ( .DIN1(n31284), .Q(n19402) );
  or2s1 U23126 ( .DIN1(n31291), .DIN2(n31296), .Q(n31944) );
  and2s1 U23127 ( .DIN1(n35451), .DIN2(n4529), .Q(n31943) );
  or2s1 U23128 ( .DIN1(n31943), .DIN2(n31944), .Q(n31284) );
  and2s1 U23129 ( .DIN1(n31284), .DIN2(n31285), .Q(n5458) );
  and2s1 U23130 ( .DIN1(n31272), .DIN2(n5448), .Q(n31288) );
  and2s1 U23131 ( .DIN1(n31291), .DIN2(n32879), .Q(n31289) );
  and2s1 U23132 ( .DIN1(n31289), .DIN2(n31290), .Q(n31287) );
  or2s1 U23133 ( .DIN1(n31287), .DIN2(n31288), .Q(n5453) );
  or2s1 U23134 ( .DIN1(n31268), .DIN2(n5453), .Q(n31286) );
  hi1s1 U23135 ( .DIN1(n31286), .Q(n5452) );
  and2s1 U23136 ( .DIN1(n31272), .DIN2(n5441), .Q(n31294) );
  and2s1 U23137 ( .DIN1(n31296), .DIN2(n35406), .Q(n31295) );
  and2s1 U23138 ( .DIN1(n31295), .DIN2(n31290), .Q(n31293) );
  or2s1 U23139 ( .DIN1(n31293), .DIN2(n31294), .Q(n5446) );
  or2s1 U23140 ( .DIN1(n31268), .DIN2(n5446), .Q(n31292) );
  hi1s1 U23141 ( .DIN1(n31292), .Q(n5445) );
  hi1s1 U23142 ( .DIN1(n35406), .Q(n31291) );
  hi1s1 U23143 ( .DIN1(n32879), .Q(n31296) );
  and2s1 U23144 ( .DIN1(n31296), .DIN2(n31291), .Q(n31299) );
  and2s1 U23145 ( .DIN1(n31290), .DIN2(n31299), .Q(n34331) );
  and2s1 U23146 ( .DIN1(n35451), .DIN2(n35406), .Q(n31945) );
  and2s1 U23147 ( .DIN1(n32879), .DIN2(n31945), .Q(n31272) );
  and2s1 U23148 ( .DIN1(n31272), .DIN2(n5434), .Q(n31298) );
  or2s1 U23149 ( .DIN1(n31298), .DIN2(n34331), .Q(n5439) );
  and2s1 U23150 ( .DIN1(u0_sp_tms[2]), .DIN2(n35282), .Q(n31949) );
  and2s1 U23151 ( .DIN1(u0_tms[2]), .DIN2(n35283), .Q(n31948) );
  or2s1 U23152 ( .DIN1(n31948), .DIN2(n31949), .Q(n35970) );
  or2s1 U23153 ( .DIN1(n35970), .DIN2(n35415), .Q(n35451) );
  hi1s1 U23154 ( .DIN1(n35451), .Q(n31290) );
  and2s1 U23155 ( .DIN1(u0_sp_tms[0]), .DIN2(n35282), .Q(n31947) );
  and2s1 U23156 ( .DIN1(u0_tms[0]), .DIN2(n35283), .Q(n31946) );
  or2s1 U23157 ( .DIN1(n31946), .DIN2(n31947), .Q(n35999) );
  or2s1 U23158 ( .DIN1(n35999), .DIN2(n35415), .Q(n35406) );
  hi1s1 U23159 ( .DIN1(u5_susp_sel_r), .Q(n34322) );
  hi1s1 U23160 ( .DIN1(rfr_ack), .Q(n34126) );
  and2s1 U23161 ( .DIN1(n34126), .DIN2(n34322), .Q(n36216) );
  hi1s1 U23162 ( .DIN1(n36216), .Q(n36214) );
  or2s1 U23163 ( .DIN1(n36346), .DIN2(n36343), .Q(n36470) );
  or2s1 U23164 ( .DIN1(u5_state[61]), .DIN2(n36471), .Q(n31956) );
  or2s1 U23165 ( .DIN1(n31956), .DIN2(n36470), .Q(n36097) );
  or2s1 U23166 ( .DIN1(u5_state[8]), .DIN2(n36097), .Q(n31955) );
  hi1s1 U23167 ( .DIN1(u5_state[1]), .Q(n31954) );
  or2s1 U23168 ( .DIN1(n31954), .DIN2(n31955), .Q(n34315) );
  hi1s1 U23169 ( .DIN1(n34315), .Q(n32870) );
  and2s1 U23170 ( .DIN1(u4_rfr_req), .DIN2(n32870), .Q(n34327) );
  hi1s1 U23171 ( .DIN1(u5_state[5]), .Q(n31960) );
  or2s1 U23172 ( .DIN1(u5_state[51]), .DIN2(n36107), .Q(n31961) );
  or2s1 U23173 ( .DIN1(u5_state[29]), .DIN2(n36369), .Q(n31963) );
  or2s1 U23174 ( .DIN1(n31962), .DIN2(n31963), .Q(n36108) );
  or2s1 U23175 ( .DIN1(n36108), .DIN2(n31961), .Q(n36128) );
  or2s1 U23176 ( .DIN1(n36128), .DIN2(n31960), .Q(n31959) );
  or2s1 U23177 ( .DIN1(u5_state[62]), .DIN2(u5_state[57]), .Q(n31958) );
  or2s1 U23178 ( .DIN1(n31958), .DIN2(n31959), .Q(n31957) );
  hi1s1 U23179 ( .DIN1(n31957), .Q(n34125) );
  and2s1 U23180 ( .DIN1(n34125), .DIN2(rfr_ack), .Q(n33491) );
  or2s1 U23181 ( .DIN1(n33491), .DIN2(n34327), .Q(n31953) );
  or2s1 U23182 ( .DIN1(n31968), .DIN2(n36193), .Q(n31967) );
  or2s1 U23183 ( .DIN1(n36194), .DIN2(n31967), .Q(n36369) );
  or2s1 U23184 ( .DIN1(n36195), .DIN2(n36369), .Q(n31966) );
  hi1s1 U23185 ( .DIN1(n31966), .Q(n31965) );
  and2s1 U23186 ( .DIN1(u5_state[29]), .DIN2(n31965), .Q(n34161) );
  or2s1 U23187 ( .DIN1(n36202), .DIN2(n31972), .Q(n36363) );
  or2s1 U23188 ( .DIN1(n31971), .DIN2(n36363), .Q(n36373) );
  or2s1 U23189 ( .DIN1(u5_state[50]), .DIN2(n36373), .Q(n31970) );
  hi1s1 U23190 ( .DIN1(n31970), .Q(n31969) );
  and2s1 U23191 ( .DIN1(u5_state[4]), .DIN2(n31969), .Q(n34254) );
  and2s1 U23192 ( .DIN1(n34254), .DIN2(rfr_ack), .Q(n35785) );
  or2s1 U23193 ( .DIN1(n35785), .DIN2(n34161), .Q(n31964) );
  or2s1 U23194 ( .DIN1(n31978), .DIN2(n31979), .Q(n31977) );
  or2s1 U23195 ( .DIN1(u5_state[24]), .DIN2(n36346), .Q(n31976) );
  or2s1 U23196 ( .DIN1(n31976), .DIN2(n31977), .Q(n36091) );
  or2s1 U23197 ( .DIN1(u5_state[20]), .DIN2(n36091), .Q(n31975) );
  or2s1 U23198 ( .DIN1(n36291), .DIN2(n31975), .Q(n36150) );
  or2s1 U23199 ( .DIN1(n36150), .DIN2(n36289), .Q(n31974) );
  hi1s1 U23200 ( .DIN1(n31974), .Q(n31973) );
  and2s1 U23201 ( .DIN1(u5_state[17]), .DIN2(n31973), .Q(n34324) );
  or2s1 U23202 ( .DIN1(n34324), .DIN2(n31964), .Q(n31952) );
  or2s1 U23203 ( .DIN1(n31952), .DIN2(n31953), .Q(u5_rfr_ack_d) );
  or2s1 U23204 ( .DIN1(u5_rfr_ack_d), .DIN2(n36214), .Q(n31951) );
  hi1s1 U23205 ( .DIN1(n9689), .Q(n31950) );
  or2s1 U23206 ( .DIN1(n31950), .DIN2(n31951), .Q(n35415) );
  and2s1 U23207 ( .DIN1(u0_sp_tms[1]), .DIN2(n35282), .Q(n31981) );
  or2s1 U23208 ( .DIN1(n31979), .DIN2(n31986), .Q(n31985) );
  hi1s1 U23209 ( .DIN1(n31985), .Q(n31984) );
  and2s1 U23210 ( .DIN1(u5_state[24]), .DIN2(n31984), .Q(n34152) );
  hi1s1 U23211 ( .DIN1(u5_state[22]), .Q(n31989) );
  or2s1 U23212 ( .DIN1(u5_state[15]), .DIN2(n36465), .Q(n31990) );
  or2s1 U23213 ( .DIN1(u5_state[60]), .DIN2(u5_state[26]), .Q(n36314) );
  or2s1 U23214 ( .DIN1(n36314), .DIN2(n31990), .Q(n36117) );
  or2s1 U23215 ( .DIN1(n36117), .DIN2(n31989), .Q(n31988) );
  or2s1 U23216 ( .DIN1(u5_state[21]), .DIN2(u5_state[18]), .Q(n31987) );
  or2s1 U23217 ( .DIN1(n31987), .DIN2(n31988), .Q(n34150) );
  hi1s1 U23218 ( .DIN1(n34150), .Q(n34136) );
  or2s1 U23219 ( .DIN1(n34136), .DIN2(n34152), .Q(n31983) );
  or2s1 U23220 ( .DIN1(u5_state[32]), .DIN2(n36200), .Q(n31998) );
  or2s1 U23221 ( .DIN1(u5_state[28]), .DIN2(u5_state[25]), .Q(n32002) );
  or2s1 U23222 ( .DIN1(u5_state[23]), .DIN2(n32002), .Q(n31979) );
  or2s1 U23223 ( .DIN1(u5_state[24]), .DIN2(n31979), .Q(n32000) );
  or2s1 U23224 ( .DIN1(n32000), .DIN2(n32001), .Q(n36343) );
  or2s1 U23225 ( .DIN1(n31978), .DIN2(n36343), .Q(n36280) );
  or2s1 U23226 ( .DIN1(n31999), .DIN2(n36280), .Q(n36194) );
  or2s1 U23227 ( .DIN1(n36194), .DIN2(n31998), .Q(n31972) );
  or2s1 U23228 ( .DIN1(n36203), .DIN2(n31972), .Q(n36478) );
  or2s1 U23229 ( .DIN1(n31997), .DIN2(n36478), .Q(n36307) );
  or2s1 U23230 ( .DIN1(u5_state[34]), .DIN2(n36164), .Q(n31996) );
  or2s1 U23231 ( .DIN1(n31996), .DIN2(n36307), .Q(n36465) );
  or2s1 U23232 ( .DIN1(n36304), .DIN2(n36465), .Q(n36313) );
  hi1s1 U23233 ( .DIN1(u5_state[26]), .Q(n31995) );
  or2s1 U23234 ( .DIN1(n31995), .DIN2(n36313), .Q(n31994) );
  or2s1 U23235 ( .DIN1(u5_state[60]), .DIN2(u5_state[18]), .Q(n32003) );
  or2s1 U23236 ( .DIN1(u5_state[15]), .DIN2(n32003), .Q(n31993) );
  or2s1 U23237 ( .DIN1(n31993), .DIN2(n31994), .Q(n31992) );
  hi1s1 U23238 ( .DIN1(n31992), .Q(n36285) );
  or2s1 U23239 ( .DIN1(u5_state[25]), .DIN2(u5_state[24]), .Q(n32006) );
  or2s1 U23240 ( .DIN1(n31986), .DIN2(n32006), .Q(n36087) );
  or2s1 U23241 ( .DIN1(u5_state[28]), .DIN2(n36087), .Q(n32005) );
  hi1s1 U23242 ( .DIN1(u5_state[23]), .Q(n36086) );
  or2s1 U23243 ( .DIN1(n36086), .DIN2(n32005), .Q(n32004) );
  hi1s1 U23244 ( .DIN1(n32004), .Q(n34273) );
  or2s1 U23245 ( .DIN1(n34273), .DIN2(n36285), .Q(n31991) );
  hi1s1 U23246 ( .DIN1(u5_state[25]), .Q(n32010) );
  or2s1 U23247 ( .DIN1(u5_state[20]), .DIN2(u5_state[17]), .Q(n32012) );
  or2s1 U23248 ( .DIN1(u5_state[16]), .DIN2(u5_state[19]), .Q(n36289) );
  or2s1 U23249 ( .DIN1(n36289), .DIN2(n32012), .Q(n36089) );
  or2s1 U23250 ( .DIN1(u5_state[10]), .DIN2(u5_state[11]), .Q(n36291) );
  or2s1 U23251 ( .DIN1(n36291), .DIN2(n36089), .Q(n32001) );
  or2s1 U23252 ( .DIN1(u5_state[64]), .DIN2(u5_state[63]), .Q(n32014) );
  or2s1 U23253 ( .DIN1(u5_state[6]), .DIN2(u5_state[65]), .Q(n32013) );
  or2s1 U23254 ( .DIN1(n32013), .DIN2(n32014), .Q(n36471) );
  or2s1 U23255 ( .DIN1(u5_state[8]), .DIN2(u5_state[61]), .Q(n32015) );
  or2s1 U23256 ( .DIN1(u5_state[1]), .DIN2(n32015), .Q(n36345) );
  or2s1 U23257 ( .DIN1(n36345), .DIN2(n36471), .Q(n31978) );
  or2s1 U23258 ( .DIN1(u5_state[31]), .DIN2(u5_state[30]), .Q(n36180) );
  or2s1 U23259 ( .DIN1(u5_state[2]), .DIN2(n36180), .Q(n31968) );
  or2s1 U23260 ( .DIN1(u5_state[29]), .DIN2(n31968), .Q(n32016) );
  or2s1 U23261 ( .DIN1(u5_state[45]), .DIN2(u5_state[43]), .Q(n36425) );
  or2s1 U23262 ( .DIN1(u5_state[54]), .DIN2(u5_state[53]), .Q(n36461) );
  or2s1 U23263 ( .DIN1(n36461), .DIN2(n36425), .Q(n36107) );
  or2s1 U23264 ( .DIN1(u5_state[57]), .DIN2(u5_state[51]), .Q(n32018) );
  or2s1 U23265 ( .DIN1(u5_state[62]), .DIN2(u5_state[5]), .Q(n36109) );
  or2s1 U23266 ( .DIN1(n36109), .DIN2(n32018), .Q(n36370) );
  or2s1 U23267 ( .DIN1(n36370), .DIN2(n36107), .Q(n32017) );
  or2s1 U23268 ( .DIN1(u5_state[39]), .DIN2(u5_state[33]), .Q(n31962) );
  or2s1 U23269 ( .DIN1(n31962), .DIN2(n32017), .Q(n36195) );
  or2s1 U23270 ( .DIN1(n36195), .DIN2(n32016), .Q(n36200) );
  or2s1 U23271 ( .DIN1(u5_state[3]), .DIN2(u5_state[37]), .Q(n36451) );
  or2s1 U23272 ( .DIN1(u5_state[38]), .DIN2(u5_state[36]), .Q(n36141) );
  or2s1 U23273 ( .DIN1(u5_state[0]), .DIN2(n36141), .Q(n36124) );
  or2s1 U23274 ( .DIN1(n36124), .DIN2(n36451), .Q(n36421) );
  or2s1 U23275 ( .DIN1(u5_state[56]), .DIN2(u5_state[52]), .Q(n36418) );
  or2s1 U23276 ( .DIN1(u5_state[44]), .DIN2(n36418), .Q(n36351) );
  or2s1 U23277 ( .DIN1(u5_state[55]), .DIN2(n36351), .Q(n32022) );
  or2s1 U23278 ( .DIN1(u5_state[47]), .DIN2(u5_state[46]), .Q(n36403) );
  or2s1 U23279 ( .DIN1(n36403), .DIN2(n32022), .Q(n36395) );
  or2s1 U23280 ( .DIN1(n36395), .DIN2(n36421), .Q(n32021) );
  or2s1 U23281 ( .DIN1(u5_state[42]), .DIN2(u5_state[41]), .Q(n32023) );
  or2s1 U23282 ( .DIN1(u5_state[40]), .DIN2(n32023), .Q(n36452) );
  or2s1 U23283 ( .DIN1(u5_state[58]), .DIN2(u5_state[59]), .Q(n36455) );
  or2s1 U23284 ( .DIN1(n36455), .DIN2(n36452), .Q(n32020) );
  or2s1 U23285 ( .DIN1(n32020), .DIN2(n32021), .Q(n31997) );
  or2s1 U23286 ( .DIN1(u5_state[27]), .DIN2(u5_state[35]), .Q(n36164) );
  or2s1 U23287 ( .DIN1(u5_state[22]), .DIN2(u5_state[21]), .Q(n36304) );
  or2s1 U23288 ( .DIN1(u5_state[15]), .DIN2(n36304), .Q(n32027) );
  or2s1 U23289 ( .DIN1(u5_state[26]), .DIN2(u5_state[18]), .Q(n32026) );
  or2s1 U23290 ( .DIN1(n32026), .DIN2(n32027), .Q(n36308) );
  or2s1 U23291 ( .DIN1(n36308), .DIN2(n36164), .Q(n32025) );
  or2s1 U23292 ( .DIN1(u5_state[60]), .DIN2(u5_state[34]), .Q(n32024) );
  or2s1 U23293 ( .DIN1(n32024), .DIN2(n32025), .Q(n36477) );
  or2s1 U23294 ( .DIN1(n36477), .DIN2(n31997), .Q(n36202) );
  or2s1 U23295 ( .DIN1(u5_state[32]), .DIN2(n36202), .Q(n32019) );
  or2s1 U23296 ( .DIN1(u5_state[49]), .DIN2(u5_state[48]), .Q(n36334) );
  or2s1 U23297 ( .DIN1(u5_state[14]), .DIN2(n36334), .Q(n36138) );
  or2s1 U23298 ( .DIN1(u5_state[12]), .DIN2(u5_state[13]), .Q(n36356) );
  or2s1 U23299 ( .DIN1(n36356), .DIN2(n36138), .Q(n31971) );
  or2s1 U23300 ( .DIN1(u5_state[50]), .DIN2(u5_state[4]), .Q(n36362) );
  or2s1 U23301 ( .DIN1(n36362), .DIN2(n31971), .Q(n36203) );
  or2s1 U23302 ( .DIN1(n36203), .DIN2(n32019), .Q(n36193) );
  or2s1 U23303 ( .DIN1(n36193), .DIN2(n36200), .Q(n36279) );
  or2s1 U23304 ( .DIN1(u5_state[9]), .DIN2(u5_state[7]), .Q(n31999) );
  or2s1 U23305 ( .DIN1(n31999), .DIN2(n36279), .Q(n36346) );
  or2s1 U23306 ( .DIN1(n36346), .DIN2(n31978), .Q(n32011) );
  or2s1 U23307 ( .DIN1(n32011), .DIN2(n32001), .Q(n31986) );
  or2s1 U23308 ( .DIN1(n31986), .DIN2(n32010), .Q(n32009) );
  or2s1 U23309 ( .DIN1(u5_state[28]), .DIN2(u5_state[24]), .Q(n32028) );
  or2s1 U23310 ( .DIN1(u5_state[23]), .DIN2(n32028), .Q(n32008) );
  or2s1 U23311 ( .DIN1(n32008), .DIN2(n32009), .Q(n32007) );
  hi1s1 U23312 ( .DIN1(n32007), .Q(n34274) );
  or2s1 U23313 ( .DIN1(n34274), .DIN2(n31991), .Q(n31982) );
  or2s1 U23314 ( .DIN1(n31982), .DIN2(n31983), .Q(u5_init_ack) );
  or2s1 U23315 ( .DIN1(u5_lmr_ack), .DIN2(u5_init_ack), .Q(n35282) );
  hi1s1 U23316 ( .DIN1(n35282), .Q(n35283) );
  and2s1 U23317 ( .DIN1(u0_tms[1]), .DIN2(n35283), .Q(n31980) );
  or2s1 U23318 ( .DIN1(n31980), .DIN2(n31981), .Q(n35981) );
  or2s1 U23319 ( .DIN1(n35981), .DIN2(n35415), .Q(n32879) );
  and2s1 U23320 ( .DIN1(n32879), .DIN2(n35406), .Q(n31933) );
  or2s1 U23321 ( .DIN1(n31933), .DIN2(n31290), .Q(n31285) );
  hi1s1 U23322 ( .DIN1(n31285), .Q(n31268) );
  or2s1 U23323 ( .DIN1(n31268), .DIN2(n5439), .Q(n31297) );
  hi1s1 U23324 ( .DIN1(n31297), .Q(n5438) );
  hi1s1 U23325 ( .DIN1(n31259), .Q(n33423) );
  and2s1 U23326 ( .DIN1(n31306), .DIN2(n33423), .Q(n31305) );
  hi1s1 U23327 ( .DIN1(n31260), .Q(n33326) );
  and2s1 U23328 ( .DIN1(n31307), .DIN2(n33326), .Q(n31304) );
  or2s1 U23329 ( .DIN1(n31304), .DIN2(n31305), .Q(n31303) );
  hi1s1 U23330 ( .DIN1(n31261), .Q(n33229) );
  and2s1 U23331 ( .DIN1(n31310), .DIN2(n33229), .Q(n31309) );
  hi1s1 U23332 ( .DIN1(n31262), .Q(n33132) );
  and2s1 U23333 ( .DIN1(n31311), .DIN2(n33132), .Q(n31308) );
  or2s1 U23334 ( .DIN1(n31308), .DIN2(n31309), .Q(n31302) );
  or2s1 U23335 ( .DIN1(n31302), .DIN2(n31303), .Q(n5432) );
  hi1s1 U23336 ( .DIN1(n5432), .Q(n31301) );
  and2s1 U23337 ( .DIN1(n31300), .DIN2(n31301), .Q(n5431) );
  hi1s1 U23338 ( .DIN1(n31255), .Q(n33420) );
  and2s1 U23339 ( .DIN1(n31306), .DIN2(n33420), .Q(n31316) );
  hi1s1 U23340 ( .DIN1(n31256), .Q(n33323) );
  and2s1 U23341 ( .DIN1(n31307), .DIN2(n33323), .Q(n31315) );
  or2s1 U23342 ( .DIN1(n31315), .DIN2(n31316), .Q(n31314) );
  hi1s1 U23343 ( .DIN1(n31257), .Q(n33226) );
  and2s1 U23344 ( .DIN1(n31310), .DIN2(n33226), .Q(n31318) );
  hi1s1 U23345 ( .DIN1(n31258), .Q(n33129) );
  and2s1 U23346 ( .DIN1(n31311), .DIN2(n33129), .Q(n31317) );
  or2s1 U23347 ( .DIN1(n31317), .DIN2(n31318), .Q(n31313) );
  or2s1 U23348 ( .DIN1(n31313), .DIN2(n31314), .Q(n5428) );
  hi1s1 U23349 ( .DIN1(n5428), .Q(n31312) );
  and2s1 U23350 ( .DIN1(n31300), .DIN2(n31312), .Q(n5427) );
  hi1s1 U23351 ( .DIN1(n31251), .Q(n33417) );
  and2s1 U23352 ( .DIN1(n31306), .DIN2(n33417), .Q(n31323) );
  hi1s1 U23353 ( .DIN1(n31252), .Q(n33320) );
  and2s1 U23354 ( .DIN1(n31307), .DIN2(n33320), .Q(n31322) );
  or2s1 U23355 ( .DIN1(n31322), .DIN2(n31323), .Q(n31321) );
  hi1s1 U23356 ( .DIN1(n31253), .Q(n33223) );
  and2s1 U23357 ( .DIN1(n31310), .DIN2(n33223), .Q(n31325) );
  hi1s1 U23358 ( .DIN1(n31254), .Q(n33126) );
  and2s1 U23359 ( .DIN1(n31311), .DIN2(n33126), .Q(n31324) );
  or2s1 U23360 ( .DIN1(n31324), .DIN2(n31325), .Q(n31320) );
  or2s1 U23361 ( .DIN1(n31320), .DIN2(n31321), .Q(n5424) );
  hi1s1 U23362 ( .DIN1(n5424), .Q(n31319) );
  and2s1 U23363 ( .DIN1(n31300), .DIN2(n31319), .Q(n5423) );
  hi1s1 U23364 ( .DIN1(n31247), .Q(n33414) );
  and2s1 U23365 ( .DIN1(n31306), .DIN2(n33414), .Q(n31330) );
  hi1s1 U23366 ( .DIN1(n31248), .Q(n33317) );
  and2s1 U23367 ( .DIN1(n31307), .DIN2(n33317), .Q(n31329) );
  or2s1 U23368 ( .DIN1(n31329), .DIN2(n31330), .Q(n31328) );
  hi1s1 U23369 ( .DIN1(n31249), .Q(n33220) );
  and2s1 U23370 ( .DIN1(n31310), .DIN2(n33220), .Q(n31332) );
  hi1s1 U23371 ( .DIN1(n31250), .Q(n33123) );
  and2s1 U23372 ( .DIN1(n31311), .DIN2(n33123), .Q(n31331) );
  or2s1 U23373 ( .DIN1(n31331), .DIN2(n31332), .Q(n31327) );
  or2s1 U23374 ( .DIN1(n31327), .DIN2(n31328), .Q(n5420) );
  hi1s1 U23375 ( .DIN1(n5420), .Q(n31326) );
  and2s1 U23376 ( .DIN1(n31300), .DIN2(n31326), .Q(n5419) );
  hi1s1 U23377 ( .DIN1(n31243), .Q(n33411) );
  and2s1 U23378 ( .DIN1(n31306), .DIN2(n33411), .Q(n31337) );
  hi1s1 U23379 ( .DIN1(n31244), .Q(n33314) );
  and2s1 U23380 ( .DIN1(n31307), .DIN2(n33314), .Q(n31336) );
  or2s1 U23381 ( .DIN1(n31336), .DIN2(n31337), .Q(n31335) );
  hi1s1 U23382 ( .DIN1(n31245), .Q(n33217) );
  and2s1 U23383 ( .DIN1(n31310), .DIN2(n33217), .Q(n31339) );
  hi1s1 U23384 ( .DIN1(n31246), .Q(n33120) );
  and2s1 U23385 ( .DIN1(n31311), .DIN2(n33120), .Q(n31338) );
  or2s1 U23386 ( .DIN1(n31338), .DIN2(n31339), .Q(n31334) );
  or2s1 U23387 ( .DIN1(n31334), .DIN2(n31335), .Q(n5416) );
  hi1s1 U23388 ( .DIN1(n5416), .Q(n31333) );
  and2s1 U23389 ( .DIN1(n31300), .DIN2(n31333), .Q(n5415) );
  hi1s1 U23390 ( .DIN1(n31239), .Q(n33408) );
  and2s1 U23391 ( .DIN1(n31306), .DIN2(n33408), .Q(n31344) );
  hi1s1 U23392 ( .DIN1(n31240), .Q(n33311) );
  and2s1 U23393 ( .DIN1(n31307), .DIN2(n33311), .Q(n31343) );
  or2s1 U23394 ( .DIN1(n31343), .DIN2(n31344), .Q(n31342) );
  hi1s1 U23395 ( .DIN1(n31241), .Q(n33214) );
  and2s1 U23396 ( .DIN1(n31310), .DIN2(n33214), .Q(n31346) );
  hi1s1 U23397 ( .DIN1(n31242), .Q(n33117) );
  and2s1 U23398 ( .DIN1(n31311), .DIN2(n33117), .Q(n31345) );
  or2s1 U23399 ( .DIN1(n31345), .DIN2(n31346), .Q(n31341) );
  or2s1 U23400 ( .DIN1(n31341), .DIN2(n31342), .Q(n5412) );
  hi1s1 U23401 ( .DIN1(n5412), .Q(n31340) );
  and2s1 U23402 ( .DIN1(n31300), .DIN2(n31340), .Q(n5411) );
  hi1s1 U23403 ( .DIN1(n31235), .Q(n33405) );
  and2s1 U23404 ( .DIN1(n31306), .DIN2(n33405), .Q(n31351) );
  hi1s1 U23405 ( .DIN1(n31236), .Q(n33308) );
  and2s1 U23406 ( .DIN1(n31307), .DIN2(n33308), .Q(n31350) );
  or2s1 U23407 ( .DIN1(n31350), .DIN2(n31351), .Q(n31349) );
  hi1s1 U23408 ( .DIN1(n31237), .Q(n33211) );
  and2s1 U23409 ( .DIN1(n31310), .DIN2(n33211), .Q(n31353) );
  hi1s1 U23410 ( .DIN1(n31238), .Q(n33114) );
  and2s1 U23411 ( .DIN1(n31311), .DIN2(n33114), .Q(n31352) );
  or2s1 U23412 ( .DIN1(n31352), .DIN2(n31353), .Q(n31348) );
  or2s1 U23413 ( .DIN1(n31348), .DIN2(n31349), .Q(n5408) );
  hi1s1 U23414 ( .DIN1(n5408), .Q(n31347) );
  and2s1 U23415 ( .DIN1(n31300), .DIN2(n31347), .Q(n5407) );
  hi1s1 U23416 ( .DIN1(n31231), .Q(n33402) );
  and2s1 U23417 ( .DIN1(n31306), .DIN2(n33402), .Q(n31358) );
  hi1s1 U23418 ( .DIN1(n31232), .Q(n33305) );
  and2s1 U23419 ( .DIN1(n31307), .DIN2(n33305), .Q(n31357) );
  or2s1 U23420 ( .DIN1(n31357), .DIN2(n31358), .Q(n31356) );
  hi1s1 U23421 ( .DIN1(n31233), .Q(n33208) );
  and2s1 U23422 ( .DIN1(n31310), .DIN2(n33208), .Q(n31360) );
  hi1s1 U23423 ( .DIN1(n31234), .Q(n33111) );
  and2s1 U23424 ( .DIN1(n31311), .DIN2(n33111), .Q(n31359) );
  or2s1 U23425 ( .DIN1(n31359), .DIN2(n31360), .Q(n31355) );
  or2s1 U23426 ( .DIN1(n31355), .DIN2(n31356), .Q(n5404) );
  hi1s1 U23427 ( .DIN1(n5404), .Q(n31354) );
  and2s1 U23428 ( .DIN1(n31300), .DIN2(n31354), .Q(n5403) );
  hi1s1 U23429 ( .DIN1(n31227), .Q(n33399) );
  and2s1 U23430 ( .DIN1(n31306), .DIN2(n33399), .Q(n31365) );
  hi1s1 U23431 ( .DIN1(n31228), .Q(n33302) );
  and2s1 U23432 ( .DIN1(n31307), .DIN2(n33302), .Q(n31364) );
  or2s1 U23433 ( .DIN1(n31364), .DIN2(n31365), .Q(n31363) );
  hi1s1 U23434 ( .DIN1(n31229), .Q(n33205) );
  and2s1 U23435 ( .DIN1(n31310), .DIN2(n33205), .Q(n31367) );
  hi1s1 U23436 ( .DIN1(n31230), .Q(n33108) );
  and2s1 U23437 ( .DIN1(n31311), .DIN2(n33108), .Q(n31366) );
  or2s1 U23438 ( .DIN1(n31366), .DIN2(n31367), .Q(n31362) );
  or2s1 U23439 ( .DIN1(n31362), .DIN2(n31363), .Q(n5400) );
  hi1s1 U23440 ( .DIN1(n5400), .Q(n31361) );
  and2s1 U23441 ( .DIN1(n31300), .DIN2(n31361), .Q(n5399) );
  hi1s1 U23442 ( .DIN1(n31223), .Q(n33396) );
  and2s1 U23443 ( .DIN1(n31306), .DIN2(n33396), .Q(n31372) );
  hi1s1 U23444 ( .DIN1(n31224), .Q(n33299) );
  and2s1 U23445 ( .DIN1(n31307), .DIN2(n33299), .Q(n31371) );
  or2s1 U23446 ( .DIN1(n31371), .DIN2(n31372), .Q(n31370) );
  hi1s1 U23447 ( .DIN1(n31225), .Q(n33202) );
  and2s1 U23448 ( .DIN1(n31310), .DIN2(n33202), .Q(n31374) );
  hi1s1 U23449 ( .DIN1(n31226), .Q(n33105) );
  and2s1 U23450 ( .DIN1(n31311), .DIN2(n33105), .Q(n31373) );
  or2s1 U23451 ( .DIN1(n31373), .DIN2(n31374), .Q(n31369) );
  or2s1 U23452 ( .DIN1(n31369), .DIN2(n31370), .Q(n5396) );
  hi1s1 U23453 ( .DIN1(n5396), .Q(n31368) );
  and2s1 U23454 ( .DIN1(n31300), .DIN2(n31368), .Q(n5395) );
  hi1s1 U23455 ( .DIN1(n31219), .Q(n33393) );
  and2s1 U23456 ( .DIN1(n31306), .DIN2(n33393), .Q(n31379) );
  hi1s1 U23457 ( .DIN1(n31220), .Q(n33296) );
  and2s1 U23458 ( .DIN1(n31307), .DIN2(n33296), .Q(n31378) );
  or2s1 U23459 ( .DIN1(n31378), .DIN2(n31379), .Q(n31377) );
  hi1s1 U23460 ( .DIN1(n31221), .Q(n33199) );
  and2s1 U23461 ( .DIN1(n31310), .DIN2(n33199), .Q(n31381) );
  hi1s1 U23462 ( .DIN1(n31222), .Q(n33102) );
  and2s1 U23463 ( .DIN1(n31311), .DIN2(n33102), .Q(n31380) );
  or2s1 U23464 ( .DIN1(n31380), .DIN2(n31381), .Q(n31376) );
  or2s1 U23465 ( .DIN1(n31376), .DIN2(n31377), .Q(n5392) );
  hi1s1 U23466 ( .DIN1(n5392), .Q(n31375) );
  and2s1 U23467 ( .DIN1(n31300), .DIN2(n31375), .Q(n5391) );
  hi1s1 U23468 ( .DIN1(n31215), .Q(n33390) );
  and2s1 U23469 ( .DIN1(n31306), .DIN2(n33390), .Q(n31386) );
  hi1s1 U23470 ( .DIN1(n31216), .Q(n33293) );
  and2s1 U23471 ( .DIN1(n31307), .DIN2(n33293), .Q(n31385) );
  or2s1 U23472 ( .DIN1(n31385), .DIN2(n31386), .Q(n31384) );
  hi1s1 U23473 ( .DIN1(n31217), .Q(n33196) );
  and2s1 U23474 ( .DIN1(n31310), .DIN2(n33196), .Q(n31388) );
  hi1s1 U23475 ( .DIN1(n31218), .Q(n33099) );
  and2s1 U23476 ( .DIN1(n31311), .DIN2(n33099), .Q(n31387) );
  or2s1 U23477 ( .DIN1(n31387), .DIN2(n31388), .Q(n31383) );
  or2s1 U23478 ( .DIN1(n31383), .DIN2(n31384), .Q(n5388) );
  hi1s1 U23479 ( .DIN1(n5388), .Q(n31382) );
  and2s1 U23480 ( .DIN1(n31300), .DIN2(n31382), .Q(n5387) );
  hi1s1 U23481 ( .DIN1(n31211), .Q(n33387) );
  and2s1 U23482 ( .DIN1(n31306), .DIN2(n33387), .Q(n31393) );
  hi1s1 U23483 ( .DIN1(n31212), .Q(n33290) );
  and2s1 U23484 ( .DIN1(n31307), .DIN2(n33290), .Q(n31392) );
  or2s1 U23485 ( .DIN1(n31392), .DIN2(n31393), .Q(n31391) );
  hi1s1 U23486 ( .DIN1(n31213), .Q(n33193) );
  and2s1 U23487 ( .DIN1(n31310), .DIN2(n33193), .Q(n31395) );
  hi1s1 U23488 ( .DIN1(n31214), .Q(n33096) );
  and2s1 U23489 ( .DIN1(n31311), .DIN2(n33096), .Q(n31394) );
  or2s1 U23490 ( .DIN1(n31394), .DIN2(n31395), .Q(n31390) );
  or2s1 U23491 ( .DIN1(n31390), .DIN2(n31391), .Q(n5384) );
  hi1s1 U23492 ( .DIN1(n5384), .Q(n31389) );
  and2s1 U23493 ( .DIN1(n31300), .DIN2(n31389), .Q(n5383) );
  hi1s1 U23494 ( .DIN1(n31207), .Q(n33384) );
  and2s1 U23495 ( .DIN1(n31306), .DIN2(n33384), .Q(n31400) );
  hi1s1 U23496 ( .DIN1(n31208), .Q(n33287) );
  and2s1 U23497 ( .DIN1(n31307), .DIN2(n33287), .Q(n31399) );
  or2s1 U23498 ( .DIN1(n31399), .DIN2(n31400), .Q(n31398) );
  hi1s1 U23499 ( .DIN1(n31209), .Q(n33190) );
  and2s1 U23500 ( .DIN1(n31310), .DIN2(n33190), .Q(n31402) );
  hi1s1 U23501 ( .DIN1(n31210), .Q(n33093) );
  and2s1 U23502 ( .DIN1(n31311), .DIN2(n33093), .Q(n31401) );
  or2s1 U23503 ( .DIN1(n31401), .DIN2(n31402), .Q(n31397) );
  or2s1 U23504 ( .DIN1(n31397), .DIN2(n31398), .Q(n5380) );
  hi1s1 U23505 ( .DIN1(n5380), .Q(n31396) );
  and2s1 U23506 ( .DIN1(n31300), .DIN2(n31396), .Q(n5379) );
  hi1s1 U23507 ( .DIN1(n31203), .Q(n33381) );
  and2s1 U23508 ( .DIN1(n31306), .DIN2(n33381), .Q(n31407) );
  hi1s1 U23509 ( .DIN1(n31204), .Q(n33284) );
  and2s1 U23510 ( .DIN1(n31307), .DIN2(n33284), .Q(n31406) );
  or2s1 U23511 ( .DIN1(n31406), .DIN2(n31407), .Q(n31405) );
  hi1s1 U23512 ( .DIN1(n31205), .Q(n33187) );
  and2s1 U23513 ( .DIN1(n31310), .DIN2(n33187), .Q(n31409) );
  hi1s1 U23514 ( .DIN1(n31206), .Q(n33090) );
  and2s1 U23515 ( .DIN1(n31311), .DIN2(n33090), .Q(n31408) );
  or2s1 U23516 ( .DIN1(n31408), .DIN2(n31409), .Q(n31404) );
  or2s1 U23517 ( .DIN1(n31404), .DIN2(n31405), .Q(n5376) );
  hi1s1 U23518 ( .DIN1(n5376), .Q(n31403) );
  and2s1 U23519 ( .DIN1(n31300), .DIN2(n31403), .Q(n5375) );
  hi1s1 U23520 ( .DIN1(n31199), .Q(n33378) );
  and2s1 U23521 ( .DIN1(n31306), .DIN2(n33378), .Q(n31414) );
  hi1s1 U23522 ( .DIN1(n31200), .Q(n33281) );
  and2s1 U23523 ( .DIN1(n31307), .DIN2(n33281), .Q(n31413) );
  or2s1 U23524 ( .DIN1(n31413), .DIN2(n31414), .Q(n31412) );
  hi1s1 U23525 ( .DIN1(n31201), .Q(n33184) );
  and2s1 U23526 ( .DIN1(n31310), .DIN2(n33184), .Q(n31416) );
  hi1s1 U23527 ( .DIN1(n31202), .Q(n33087) );
  and2s1 U23528 ( .DIN1(n31311), .DIN2(n33087), .Q(n31415) );
  or2s1 U23529 ( .DIN1(n31415), .DIN2(n31416), .Q(n31411) );
  or2s1 U23530 ( .DIN1(n31411), .DIN2(n31412), .Q(n5372) );
  hi1s1 U23531 ( .DIN1(n5372), .Q(n31410) );
  and2s1 U23532 ( .DIN1(n31300), .DIN2(n31410), .Q(n5371) );
  hi1s1 U23533 ( .DIN1(n31195), .Q(n33375) );
  and2s1 U23534 ( .DIN1(n31306), .DIN2(n33375), .Q(n31421) );
  hi1s1 U23535 ( .DIN1(n31196), .Q(n33278) );
  and2s1 U23536 ( .DIN1(n31307), .DIN2(n33278), .Q(n31420) );
  or2s1 U23537 ( .DIN1(n31420), .DIN2(n31421), .Q(n31419) );
  hi1s1 U23538 ( .DIN1(n31197), .Q(n33181) );
  and2s1 U23539 ( .DIN1(n31310), .DIN2(n33181), .Q(n31423) );
  hi1s1 U23540 ( .DIN1(n31198), .Q(n33084) );
  and2s1 U23541 ( .DIN1(n31311), .DIN2(n33084), .Q(n31422) );
  or2s1 U23542 ( .DIN1(n31422), .DIN2(n31423), .Q(n31418) );
  or2s1 U23543 ( .DIN1(n31418), .DIN2(n31419), .Q(n5368) );
  hi1s1 U23544 ( .DIN1(n5368), .Q(n31417) );
  and2s1 U23545 ( .DIN1(n31300), .DIN2(n31417), .Q(n5367) );
  hi1s1 U23546 ( .DIN1(n31191), .Q(n33372) );
  and2s1 U23547 ( .DIN1(n31306), .DIN2(n33372), .Q(n31428) );
  hi1s1 U23548 ( .DIN1(n31192), .Q(n33275) );
  and2s1 U23549 ( .DIN1(n31307), .DIN2(n33275), .Q(n31427) );
  or2s1 U23550 ( .DIN1(n31427), .DIN2(n31428), .Q(n31426) );
  hi1s1 U23551 ( .DIN1(n31193), .Q(n33178) );
  and2s1 U23552 ( .DIN1(n31310), .DIN2(n33178), .Q(n31430) );
  hi1s1 U23553 ( .DIN1(n31194), .Q(n33081) );
  and2s1 U23554 ( .DIN1(n31311), .DIN2(n33081), .Q(n31429) );
  or2s1 U23555 ( .DIN1(n31429), .DIN2(n31430), .Q(n31425) );
  or2s1 U23556 ( .DIN1(n31425), .DIN2(n31426), .Q(n5364) );
  hi1s1 U23557 ( .DIN1(n5364), .Q(n31424) );
  and2s1 U23558 ( .DIN1(n31300), .DIN2(n31424), .Q(n5363) );
  hi1s1 U23559 ( .DIN1(n31187), .Q(n33369) );
  and2s1 U23560 ( .DIN1(n31306), .DIN2(n33369), .Q(n31435) );
  hi1s1 U23561 ( .DIN1(n31188), .Q(n33272) );
  and2s1 U23562 ( .DIN1(n31307), .DIN2(n33272), .Q(n31434) );
  or2s1 U23563 ( .DIN1(n31434), .DIN2(n31435), .Q(n31433) );
  hi1s1 U23564 ( .DIN1(n31189), .Q(n33175) );
  and2s1 U23565 ( .DIN1(n31310), .DIN2(n33175), .Q(n31437) );
  hi1s1 U23566 ( .DIN1(n31190), .Q(n33078) );
  and2s1 U23567 ( .DIN1(n31311), .DIN2(n33078), .Q(n31436) );
  or2s1 U23568 ( .DIN1(n31436), .DIN2(n31437), .Q(n31432) );
  or2s1 U23569 ( .DIN1(n31432), .DIN2(n31433), .Q(n5360) );
  hi1s1 U23570 ( .DIN1(n5360), .Q(n31431) );
  and2s1 U23571 ( .DIN1(n31300), .DIN2(n31431), .Q(n5359) );
  hi1s1 U23572 ( .DIN1(n31183), .Q(n33366) );
  and2s1 U23573 ( .DIN1(n31306), .DIN2(n33366), .Q(n31442) );
  hi1s1 U23574 ( .DIN1(n31184), .Q(n33269) );
  and2s1 U23575 ( .DIN1(n31307), .DIN2(n33269), .Q(n31441) );
  or2s1 U23576 ( .DIN1(n31441), .DIN2(n31442), .Q(n31440) );
  hi1s1 U23577 ( .DIN1(n31185), .Q(n33172) );
  and2s1 U23578 ( .DIN1(n31310), .DIN2(n33172), .Q(n31444) );
  hi1s1 U23579 ( .DIN1(n31186), .Q(n33075) );
  and2s1 U23580 ( .DIN1(n31311), .DIN2(n33075), .Q(n31443) );
  or2s1 U23581 ( .DIN1(n31443), .DIN2(n31444), .Q(n31439) );
  or2s1 U23582 ( .DIN1(n31439), .DIN2(n31440), .Q(n5356) );
  hi1s1 U23583 ( .DIN1(n5356), .Q(n31438) );
  and2s1 U23584 ( .DIN1(n31300), .DIN2(n31438), .Q(n5355) );
  hi1s1 U23585 ( .DIN1(n31179), .Q(n33363) );
  and2s1 U23586 ( .DIN1(n31306), .DIN2(n33363), .Q(n31449) );
  hi1s1 U23587 ( .DIN1(n31180), .Q(n33266) );
  and2s1 U23588 ( .DIN1(n31307), .DIN2(n33266), .Q(n31448) );
  or2s1 U23589 ( .DIN1(n31448), .DIN2(n31449), .Q(n31447) );
  hi1s1 U23590 ( .DIN1(n31181), .Q(n33169) );
  and2s1 U23591 ( .DIN1(n31310), .DIN2(n33169), .Q(n31451) );
  hi1s1 U23592 ( .DIN1(n31182), .Q(n33072) );
  and2s1 U23593 ( .DIN1(n31311), .DIN2(n33072), .Q(n31450) );
  or2s1 U23594 ( .DIN1(n31450), .DIN2(n31451), .Q(n31446) );
  or2s1 U23595 ( .DIN1(n31446), .DIN2(n31447), .Q(n5352) );
  hi1s1 U23596 ( .DIN1(n5352), .Q(n31445) );
  and2s1 U23597 ( .DIN1(n31300), .DIN2(n31445), .Q(n5351) );
  hi1s1 U23598 ( .DIN1(n31175), .Q(n33360) );
  and2s1 U23599 ( .DIN1(n31306), .DIN2(n33360), .Q(n31456) );
  hi1s1 U23600 ( .DIN1(n31176), .Q(n33263) );
  and2s1 U23601 ( .DIN1(n31307), .DIN2(n33263), .Q(n31455) );
  or2s1 U23602 ( .DIN1(n31455), .DIN2(n31456), .Q(n31454) );
  hi1s1 U23603 ( .DIN1(n31177), .Q(n33166) );
  and2s1 U23604 ( .DIN1(n31310), .DIN2(n33166), .Q(n31458) );
  hi1s1 U23605 ( .DIN1(n31178), .Q(n33069) );
  and2s1 U23606 ( .DIN1(n31311), .DIN2(n33069), .Q(n31457) );
  or2s1 U23607 ( .DIN1(n31457), .DIN2(n31458), .Q(n31453) );
  or2s1 U23608 ( .DIN1(n31453), .DIN2(n31454), .Q(n5348) );
  hi1s1 U23609 ( .DIN1(n5348), .Q(n31452) );
  and2s1 U23610 ( .DIN1(n31300), .DIN2(n31452), .Q(n5347) );
  hi1s1 U23611 ( .DIN1(n31171), .Q(n33357) );
  and2s1 U23612 ( .DIN1(n31306), .DIN2(n33357), .Q(n31463) );
  hi1s1 U23613 ( .DIN1(n31172), .Q(n33260) );
  and2s1 U23614 ( .DIN1(n31307), .DIN2(n33260), .Q(n31462) );
  or2s1 U23615 ( .DIN1(n31462), .DIN2(n31463), .Q(n31461) );
  hi1s1 U23616 ( .DIN1(n31173), .Q(n33163) );
  and2s1 U23617 ( .DIN1(n31310), .DIN2(n33163), .Q(n31465) );
  hi1s1 U23618 ( .DIN1(n31174), .Q(n33066) );
  and2s1 U23619 ( .DIN1(n31311), .DIN2(n33066), .Q(n31464) );
  or2s1 U23620 ( .DIN1(n31464), .DIN2(n31465), .Q(n31460) );
  or2s1 U23621 ( .DIN1(n31460), .DIN2(n31461), .Q(n5344) );
  hi1s1 U23622 ( .DIN1(n5344), .Q(n31459) );
  and2s1 U23623 ( .DIN1(n31300), .DIN2(n31459), .Q(n5343) );
  hi1s1 U23624 ( .DIN1(n31167), .Q(n33354) );
  and2s1 U23625 ( .DIN1(n31306), .DIN2(n33354), .Q(n31470) );
  hi1s1 U23626 ( .DIN1(n31168), .Q(n33257) );
  and2s1 U23627 ( .DIN1(n31307), .DIN2(n33257), .Q(n31469) );
  or2s1 U23628 ( .DIN1(n31469), .DIN2(n31470), .Q(n31468) );
  hi1s1 U23629 ( .DIN1(n31169), .Q(n33160) );
  and2s1 U23630 ( .DIN1(n31310), .DIN2(n33160), .Q(n31472) );
  hi1s1 U23631 ( .DIN1(n31170), .Q(n33063) );
  and2s1 U23632 ( .DIN1(n31311), .DIN2(n33063), .Q(n31471) );
  or2s1 U23633 ( .DIN1(n31471), .DIN2(n31472), .Q(n31467) );
  or2s1 U23634 ( .DIN1(n31467), .DIN2(n31468), .Q(n5340) );
  hi1s1 U23635 ( .DIN1(n5340), .Q(n31466) );
  and2s1 U23636 ( .DIN1(n31300), .DIN2(n31466), .Q(n5339) );
  hi1s1 U23637 ( .DIN1(n31163), .Q(n33351) );
  and2s1 U23638 ( .DIN1(n31306), .DIN2(n33351), .Q(n31477) );
  hi1s1 U23639 ( .DIN1(n31164), .Q(n33254) );
  and2s1 U23640 ( .DIN1(n31307), .DIN2(n33254), .Q(n31476) );
  or2s1 U23641 ( .DIN1(n31476), .DIN2(n31477), .Q(n31475) );
  hi1s1 U23642 ( .DIN1(n31165), .Q(n33157) );
  and2s1 U23643 ( .DIN1(n31310), .DIN2(n33157), .Q(n31479) );
  hi1s1 U23644 ( .DIN1(n31166), .Q(n33060) );
  and2s1 U23645 ( .DIN1(n31311), .DIN2(n33060), .Q(n31478) );
  or2s1 U23646 ( .DIN1(n31478), .DIN2(n31479), .Q(n31474) );
  or2s1 U23647 ( .DIN1(n31474), .DIN2(n31475), .Q(n5336) );
  hi1s1 U23648 ( .DIN1(n5336), .Q(n31473) );
  and2s1 U23649 ( .DIN1(n31300), .DIN2(n31473), .Q(n5335) );
  hi1s1 U23650 ( .DIN1(n31159), .Q(n33348) );
  and2s1 U23651 ( .DIN1(n31306), .DIN2(n33348), .Q(n31484) );
  hi1s1 U23652 ( .DIN1(n31160), .Q(n33251) );
  and2s1 U23653 ( .DIN1(n31307), .DIN2(n33251), .Q(n31483) );
  or2s1 U23654 ( .DIN1(n31483), .DIN2(n31484), .Q(n31482) );
  hi1s1 U23655 ( .DIN1(n31161), .Q(n33154) );
  and2s1 U23656 ( .DIN1(n31310), .DIN2(n33154), .Q(n31486) );
  hi1s1 U23657 ( .DIN1(n31162), .Q(n33057) );
  and2s1 U23658 ( .DIN1(n31311), .DIN2(n33057), .Q(n31485) );
  or2s1 U23659 ( .DIN1(n31485), .DIN2(n31486), .Q(n31481) );
  or2s1 U23660 ( .DIN1(n31481), .DIN2(n31482), .Q(n5332) );
  hi1s1 U23661 ( .DIN1(n5332), .Q(n31480) );
  and2s1 U23662 ( .DIN1(n31300), .DIN2(n31480), .Q(n5331) );
  hi1s1 U23663 ( .DIN1(n31155), .Q(n33345) );
  and2s1 U23664 ( .DIN1(n31306), .DIN2(n33345), .Q(n31491) );
  hi1s1 U23665 ( .DIN1(n31156), .Q(n33248) );
  and2s1 U23666 ( .DIN1(n31307), .DIN2(n33248), .Q(n31490) );
  or2s1 U23667 ( .DIN1(n31490), .DIN2(n31491), .Q(n31489) );
  hi1s1 U23668 ( .DIN1(n31157), .Q(n33151) );
  and2s1 U23669 ( .DIN1(n31310), .DIN2(n33151), .Q(n31493) );
  hi1s1 U23670 ( .DIN1(n31158), .Q(n33054) );
  and2s1 U23671 ( .DIN1(n31311), .DIN2(n33054), .Q(n31492) );
  or2s1 U23672 ( .DIN1(n31492), .DIN2(n31493), .Q(n31488) );
  or2s1 U23673 ( .DIN1(n31488), .DIN2(n31489), .Q(n5328) );
  hi1s1 U23674 ( .DIN1(n5328), .Q(n31487) );
  and2s1 U23675 ( .DIN1(n31300), .DIN2(n31487), .Q(n5327) );
  hi1s1 U23676 ( .DIN1(n31151), .Q(n33342) );
  and2s1 U23677 ( .DIN1(n31306), .DIN2(n33342), .Q(n31498) );
  hi1s1 U23678 ( .DIN1(n31152), .Q(n33245) );
  and2s1 U23679 ( .DIN1(n31307), .DIN2(n33245), .Q(n31497) );
  or2s1 U23680 ( .DIN1(n31497), .DIN2(n31498), .Q(n31496) );
  hi1s1 U23681 ( .DIN1(n31153), .Q(n33148) );
  and2s1 U23682 ( .DIN1(n31310), .DIN2(n33148), .Q(n31500) );
  hi1s1 U23683 ( .DIN1(n31154), .Q(n33051) );
  and2s1 U23684 ( .DIN1(n31311), .DIN2(n33051), .Q(n31499) );
  or2s1 U23685 ( .DIN1(n31499), .DIN2(n31500), .Q(n31495) );
  or2s1 U23686 ( .DIN1(n31495), .DIN2(n31496), .Q(n5324) );
  hi1s1 U23687 ( .DIN1(n5324), .Q(n31494) );
  and2s1 U23688 ( .DIN1(n31300), .DIN2(n31494), .Q(n5323) );
  hi1s1 U23689 ( .DIN1(n31147), .Q(n33339) );
  and2s1 U23690 ( .DIN1(n31306), .DIN2(n33339), .Q(n31505) );
  hi1s1 U23691 ( .DIN1(n31148), .Q(n33242) );
  and2s1 U23692 ( .DIN1(n31307), .DIN2(n33242), .Q(n31504) );
  or2s1 U23693 ( .DIN1(n31504), .DIN2(n31505), .Q(n31503) );
  hi1s1 U23694 ( .DIN1(n31149), .Q(n33145) );
  and2s1 U23695 ( .DIN1(n31310), .DIN2(n33145), .Q(n31507) );
  hi1s1 U23696 ( .DIN1(n31150), .Q(n33048) );
  and2s1 U23697 ( .DIN1(n31311), .DIN2(n33048), .Q(n31506) );
  or2s1 U23698 ( .DIN1(n31506), .DIN2(n31507), .Q(n31502) );
  or2s1 U23699 ( .DIN1(n31502), .DIN2(n31503), .Q(n5320) );
  hi1s1 U23700 ( .DIN1(n5320), .Q(n31501) );
  and2s1 U23701 ( .DIN1(n31300), .DIN2(n31501), .Q(n5319) );
  hi1s1 U23702 ( .DIN1(n31143), .Q(n33336) );
  and2s1 U23703 ( .DIN1(n31306), .DIN2(n33336), .Q(n31512) );
  hi1s1 U23704 ( .DIN1(n31144), .Q(n33239) );
  and2s1 U23705 ( .DIN1(n31307), .DIN2(n33239), .Q(n31511) );
  or2s1 U23706 ( .DIN1(n31511), .DIN2(n31512), .Q(n31510) );
  hi1s1 U23707 ( .DIN1(n31145), .Q(n33142) );
  and2s1 U23708 ( .DIN1(n31310), .DIN2(n33142), .Q(n31514) );
  hi1s1 U23709 ( .DIN1(n31146), .Q(n33045) );
  and2s1 U23710 ( .DIN1(n31311), .DIN2(n33045), .Q(n31513) );
  or2s1 U23711 ( .DIN1(n31513), .DIN2(n31514), .Q(n31509) );
  or2s1 U23712 ( .DIN1(n31509), .DIN2(n31510), .Q(n5316) );
  hi1s1 U23713 ( .DIN1(n5316), .Q(n31508) );
  and2s1 U23714 ( .DIN1(n31300), .DIN2(n31508), .Q(n5315) );
  hi1s1 U23715 ( .DIN1(n31139), .Q(n33333) );
  and2s1 U23716 ( .DIN1(n31306), .DIN2(n33333), .Q(n31519) );
  hi1s1 U23717 ( .DIN1(n31140), .Q(n33236) );
  and2s1 U23718 ( .DIN1(n31307), .DIN2(n33236), .Q(n31518) );
  or2s1 U23719 ( .DIN1(n31518), .DIN2(n31519), .Q(n31517) );
  hi1s1 U23720 ( .DIN1(n31141), .Q(n33139) );
  and2s1 U23721 ( .DIN1(n31310), .DIN2(n33139), .Q(n31521) );
  hi1s1 U23722 ( .DIN1(n31142), .Q(n33042) );
  and2s1 U23723 ( .DIN1(n31311), .DIN2(n33042), .Q(n31520) );
  or2s1 U23724 ( .DIN1(n31520), .DIN2(n31521), .Q(n31516) );
  or2s1 U23725 ( .DIN1(n31516), .DIN2(n31517), .Q(n5312) );
  hi1s1 U23726 ( .DIN1(n5312), .Q(n31515) );
  and2s1 U23727 ( .DIN1(n31300), .DIN2(n31515), .Q(n5311) );
  hi1s1 U23728 ( .DIN1(n31135), .Q(n33330) );
  and2s1 U23729 ( .DIN1(n31306), .DIN2(n33330), .Q(n31526) );
  hi1s1 U23730 ( .DIN1(n31136), .Q(n33233) );
  and2s1 U23731 ( .DIN1(n31307), .DIN2(n33233), .Q(n31525) );
  or2s1 U23732 ( .DIN1(n31525), .DIN2(n31526), .Q(n31524) );
  hi1s1 U23733 ( .DIN1(n31137), .Q(n33136) );
  and2s1 U23734 ( .DIN1(n31310), .DIN2(n33136), .Q(n31528) );
  hi1s1 U23735 ( .DIN1(n31138), .Q(n33039) );
  and2s1 U23736 ( .DIN1(n31311), .DIN2(n33039), .Q(n31527) );
  or2s1 U23737 ( .DIN1(n31527), .DIN2(n31528), .Q(n31523) );
  or2s1 U23738 ( .DIN1(n31523), .DIN2(n31524), .Q(n5308) );
  hi1s1 U23739 ( .DIN1(n5308), .Q(n31522) );
  or2s1 U23740 ( .DIN1(u3_u0_rd_adr[0]), .DIN2(n31534), .Q(n31533) );
  or2s1 U23741 ( .DIN1(u3_u0_rd_adr[3]), .DIN2(u3_u0_rd_adr[2]), .Q(n31532) );
  or2s1 U23742 ( .DIN1(n31532), .DIN2(n31533), .Q(n31531) );
  hi1s1 U23743 ( .DIN1(n31531), .Q(n31310) );
  or2s1 U23744 ( .DIN1(u3_u0_rd_adr[0]), .DIN2(n31538), .Q(n31537) );
  or2s1 U23745 ( .DIN1(u3_u0_rd_adr[3]), .DIN2(u3_u0_rd_adr[1]), .Q(n31536) );
  or2s1 U23746 ( .DIN1(n31536), .DIN2(n31537), .Q(n31535) );
  hi1s1 U23747 ( .DIN1(n31535), .Q(n31307) );
  or2s1 U23748 ( .DIN1(n31307), .DIN2(n31310), .Q(n31530) );
  or2s1 U23749 ( .DIN1(u3_u0_rd_adr[0]), .DIN2(n31542), .Q(n31541) );
  or2s1 U23750 ( .DIN1(u3_u0_rd_adr[2]), .DIN2(u3_u0_rd_adr[1]), .Q(n31540) );
  or2s1 U23751 ( .DIN1(n31540), .DIN2(n31541), .Q(n31539) );
  hi1s1 U23752 ( .DIN1(n31539), .Q(n31306) );
  hi1s1 U23753 ( .DIN1(u3_u0_rd_adr[1]), .Q(n31534) );
  and2s1 U23754 ( .DIN1(n31534), .DIN2(u3_u0_rd_adr[0]), .Q(n31544) );
  hi1s1 U23755 ( .DIN1(u3_u0_rd_adr[2]), .Q(n31538) );
  hi1s1 U23756 ( .DIN1(u3_u0_rd_adr[3]), .Q(n31542) );
  and2s1 U23757 ( .DIN1(n31542), .DIN2(n31538), .Q(n31543) );
  and2s1 U23758 ( .DIN1(n31543), .DIN2(n31544), .Q(n31311) );
  or2s1 U23759 ( .DIN1(n31311), .DIN2(n31306), .Q(n31529) );
  or2s1 U23760 ( .DIN1(n31529), .DIN2(n31530), .Q(n31300) );
  and2s1 U23761 ( .DIN1(n31300), .DIN2(n31522), .Q(n5307) );
  hi1s1 U23762 ( .DIN1(n31130), .Q(n32326) );
  and2s1 U23763 ( .DIN1(n31553), .DIN2(n32326), .Q(n31552) );
  hi1s1 U23764 ( .DIN1(n31131), .Q(n32092) );
  and2s1 U23765 ( .DIN1(n31554), .DIN2(n32092), .Q(n31551) );
  or2s1 U23766 ( .DIN1(n31551), .DIN2(n31552), .Q(n31550) );
  hi1s1 U23767 ( .DIN1(n31132), .Q(n32842) );
  and2s1 U23768 ( .DIN1(n31555), .DIN2(n32842), .Q(n31549) );
  or2s1 U23769 ( .DIN1(n31549), .DIN2(n31550), .Q(n31548) );
  and2s1 U23770 ( .DIN1(n31560), .DIN2(poc_o[4]), .Q(n31559) );
  hi1s1 U23771 ( .DIN1(n31133), .Q(n32419) );
  and2s1 U23772 ( .DIN1(n31561), .DIN2(n32419), .Q(n31558) );
  or2s1 U23773 ( .DIN1(n31558), .DIN2(n31559), .Q(n31557) );
  hi1s1 U23774 ( .DIN1(n31134), .Q(n32516) );
  and2s1 U23775 ( .DIN1(n31564), .DIN2(n32516), .Q(n31563) );
  and2s1 U23776 ( .DIN1(n31565), .DIN2(u0_csc_mask_r[4]), .Q(n31562) );
  or2s1 U23777 ( .DIN1(n31562), .DIN2(n31563), .Q(n31556) );
  or2s1 U23778 ( .DIN1(n31556), .DIN2(n31557), .Q(n31547) );
  or2s1 U23779 ( .DIN1(n31547), .DIN2(n31548), .Q(n5304) );
  hi1s1 U23780 ( .DIN1(n5304), .Q(n31546) );
  and2s1 U23781 ( .DIN1(n31545), .DIN2(n31546), .Q(n5303) );
  hi1s1 U23782 ( .DIN1(n31127), .Q(n32342) );
  and2s1 U23783 ( .DIN1(n31553), .DIN2(n32342), .Q(n31572) );
  hi1s1 U23784 ( .DIN1(n31128), .Q(n32642) );
  and2s1 U23785 ( .DIN1(n31554), .DIN2(n32642), .Q(n31571) );
  or2s1 U23786 ( .DIN1(n31571), .DIN2(n31572), .Q(n31570) );
  and2s1 U23787 ( .DIN1(n31555), .DIN2(u0_csc0[0]), .Q(n31569) );
  or2s1 U23788 ( .DIN1(n31569), .DIN2(n31570), .Q(n31568) );
  and2s1 U23789 ( .DIN1(n31560), .DIN2(poc_o[0]), .Q(n31576) );
  and2s1 U23790 ( .DIN1(n31561), .DIN2(u0_csc1[0]), .Q(n31575) );
  or2s1 U23791 ( .DIN1(n31575), .DIN2(n31576), .Q(n31574) );
  hi1s1 U23792 ( .DIN1(n31129), .Q(n32528) );
  and2s1 U23793 ( .DIN1(n31564), .DIN2(n32528), .Q(n31578) );
  and2s1 U23794 ( .DIN1(n31565), .DIN2(u0_csc_mask_r[0]), .Q(n31577) );
  or2s1 U23795 ( .DIN1(n31577), .DIN2(n31578), .Q(n31573) );
  or2s1 U23796 ( .DIN1(n31573), .DIN2(n31574), .Q(n31567) );
  or2s1 U23797 ( .DIN1(n31567), .DIN2(n31568), .Q(n5300) );
  hi1s1 U23798 ( .DIN1(n5300), .Q(n31566) );
  and2s1 U23799 ( .DIN1(n31545), .DIN2(n31566), .Q(n5299) );
  hi1s1 U23800 ( .DIN1(n31122), .Q(n32322) );
  and2s1 U23801 ( .DIN1(n31553), .DIN2(n32322), .Q(n31585) );
  hi1s1 U23802 ( .DIN1(n31123), .Q(n32089) );
  and2s1 U23803 ( .DIN1(n31554), .DIN2(n32089), .Q(n31584) );
  or2s1 U23804 ( .DIN1(n31584), .DIN2(n31585), .Q(n31583) );
  hi1s1 U23805 ( .DIN1(n31124), .Q(n32834) );
  and2s1 U23806 ( .DIN1(n31555), .DIN2(n32834), .Q(n31582) );
  or2s1 U23807 ( .DIN1(n31582), .DIN2(n31583), .Q(n31581) );
  and2s1 U23808 ( .DIN1(n31560), .DIN2(poc_o[5]), .Q(n31589) );
  hi1s1 U23809 ( .DIN1(n31125), .Q(n32416) );
  and2s1 U23810 ( .DIN1(n31561), .DIN2(n32416), .Q(n31588) );
  or2s1 U23811 ( .DIN1(n31588), .DIN2(n31589), .Q(n31587) );
  hi1s1 U23812 ( .DIN1(n31126), .Q(n32513) );
  and2s1 U23813 ( .DIN1(n31564), .DIN2(n32513), .Q(n31591) );
  and2s1 U23814 ( .DIN1(n31565), .DIN2(u0_csc_mask_r[5]), .Q(n31590) );
  or2s1 U23815 ( .DIN1(n31590), .DIN2(n31591), .Q(n31586) );
  or2s1 U23816 ( .DIN1(n31586), .DIN2(n31587), .Q(n31580) );
  or2s1 U23817 ( .DIN1(n31580), .DIN2(n31581), .Q(n5296) );
  hi1s1 U23818 ( .DIN1(n5296), .Q(n31579) );
  and2s1 U23819 ( .DIN1(n31545), .DIN2(n31579), .Q(n5295) );
  hi1s1 U23820 ( .DIN1(n31117), .Q(n32338) );
  and2s1 U23821 ( .DIN1(n31553), .DIN2(n32338), .Q(n31598) );
  hi1s1 U23822 ( .DIN1(n31118), .Q(n32101) );
  and2s1 U23823 ( .DIN1(n31554), .DIN2(n32101), .Q(n31597) );
  or2s1 U23824 ( .DIN1(n31597), .DIN2(n31598), .Q(n31596) );
  hi1s1 U23825 ( .DIN1(n31119), .Q(n32750) );
  and2s1 U23826 ( .DIN1(n31555), .DIN2(n32750), .Q(n31595) );
  or2s1 U23827 ( .DIN1(n31595), .DIN2(n31596), .Q(n31594) );
  and2s1 U23828 ( .DIN1(n31560), .DIN2(poc_o[1]), .Q(n31602) );
  hi1s1 U23829 ( .DIN1(n31120), .Q(n32426) );
  and2s1 U23830 ( .DIN1(n31561), .DIN2(n32426), .Q(n31601) );
  or2s1 U23831 ( .DIN1(n31601), .DIN2(n31602), .Q(n31600) );
  hi1s1 U23832 ( .DIN1(n31121), .Q(n32525) );
  and2s1 U23833 ( .DIN1(n31564), .DIN2(n32525), .Q(n31604) );
  and2s1 U23834 ( .DIN1(n31565), .DIN2(u0_csc_mask_r[1]), .Q(n31603) );
  or2s1 U23835 ( .DIN1(n31603), .DIN2(n31604), .Q(n31599) );
  or2s1 U23836 ( .DIN1(n31599), .DIN2(n31600), .Q(n31593) );
  or2s1 U23837 ( .DIN1(n31593), .DIN2(n31594), .Q(n5292) );
  hi1s1 U23838 ( .DIN1(n5292), .Q(n31592) );
  and2s1 U23839 ( .DIN1(n31545), .DIN2(n31592), .Q(n5291) );
  hi1s1 U23840 ( .DIN1(n31115), .Q(n32334) );
  and2s1 U23841 ( .DIN1(n31553), .DIN2(n32334), .Q(n31611) );
  hi1s1 U23842 ( .DIN1(n15523), .Q(n32098) );
  and2s1 U23843 ( .DIN1(n31554), .DIN2(n32098), .Q(n31610) );
  or2s1 U23844 ( .DIN1(n31610), .DIN2(n31611), .Q(n31609) );
  and2s1 U23845 ( .DIN1(n31555), .DIN2(u0_csc0[2]), .Q(n31608) );
  or2s1 U23846 ( .DIN1(n31608), .DIN2(n31609), .Q(n31607) );
  and2s1 U23847 ( .DIN1(n31560), .DIN2(poc_o[2]), .Q(n31615) );
  and2s1 U23848 ( .DIN1(n31561), .DIN2(u0_csc1[2]), .Q(n31614) );
  or2s1 U23849 ( .DIN1(n31614), .DIN2(n31615), .Q(n31613) );
  hi1s1 U23850 ( .DIN1(n31116), .Q(n32522) );
  and2s1 U23851 ( .DIN1(n31564), .DIN2(n32522), .Q(n31617) );
  and2s1 U23852 ( .DIN1(n31565), .DIN2(u0_csc_mask_r[2]), .Q(n31616) );
  or2s1 U23853 ( .DIN1(n31616), .DIN2(n31617), .Q(n31612) );
  or2s1 U23854 ( .DIN1(n31612), .DIN2(n31613), .Q(n31606) );
  or2s1 U23855 ( .DIN1(n31606), .DIN2(n31607), .Q(n5288) );
  hi1s1 U23856 ( .DIN1(n5288), .Q(n31605) );
  and2s1 U23857 ( .DIN1(n31545), .DIN2(n31605), .Q(n5287) );
  hi1s1 U23858 ( .DIN1(n31112), .Q(n32330) );
  and2s1 U23859 ( .DIN1(n31553), .DIN2(n32330), .Q(n31624) );
  hi1s1 U23860 ( .DIN1(n31113), .Q(n32095) );
  and2s1 U23861 ( .DIN1(n31554), .DIN2(n32095), .Q(n31623) );
  or2s1 U23862 ( .DIN1(n31623), .DIN2(n31624), .Q(n31622) );
  and2s1 U23863 ( .DIN1(n31555), .DIN2(u0_csc0[3]), .Q(n31621) );
  or2s1 U23864 ( .DIN1(n31621), .DIN2(n31622), .Q(n31620) );
  and2s1 U23865 ( .DIN1(n31560), .DIN2(poc_o[3]), .Q(n31628) );
  and2s1 U23866 ( .DIN1(n31561), .DIN2(u0_csc1[3]), .Q(n31627) );
  or2s1 U23867 ( .DIN1(n31627), .DIN2(n31628), .Q(n31626) );
  hi1s1 U23868 ( .DIN1(n31114), .Q(n32519) );
  and2s1 U23869 ( .DIN1(n31564), .DIN2(n32519), .Q(n31630) );
  and2s1 U23870 ( .DIN1(n31565), .DIN2(u0_csc_mask_r[3]), .Q(n31629) );
  or2s1 U23871 ( .DIN1(n31629), .DIN2(n31630), .Q(n31625) );
  or2s1 U23872 ( .DIN1(n31625), .DIN2(n31626), .Q(n31619) );
  or2s1 U23873 ( .DIN1(n31619), .DIN2(n31620), .Q(n5284) );
  hi1s1 U23874 ( .DIN1(n5284), .Q(n31618) );
  and2s1 U23875 ( .DIN1(n31545), .DIN2(n31618), .Q(n5283) );
  hi1s1 U23876 ( .DIN1(n31107), .Q(n32318) );
  and2s1 U23877 ( .DIN1(n31553), .DIN2(n32318), .Q(n31637) );
  hi1s1 U23878 ( .DIN1(n31108), .Q(n32086) );
  and2s1 U23879 ( .DIN1(n31554), .DIN2(n32086), .Q(n31636) );
  or2s1 U23880 ( .DIN1(n31636), .DIN2(n31637), .Q(n31635) );
  hi1s1 U23881 ( .DIN1(n31109), .Q(n32210) );
  and2s1 U23882 ( .DIN1(n31555), .DIN2(n32210), .Q(n31634) );
  or2s1 U23883 ( .DIN1(n31634), .DIN2(n31635), .Q(n31633) );
  and2s1 U23884 ( .DIN1(n31560), .DIN2(poc_o[6]), .Q(n31641) );
  hi1s1 U23885 ( .DIN1(n31110), .Q(n32413) );
  and2s1 U23886 ( .DIN1(n31561), .DIN2(n32413), .Q(n31640) );
  or2s1 U23887 ( .DIN1(n31640), .DIN2(n31641), .Q(n31639) );
  hi1s1 U23888 ( .DIN1(n31111), .Q(n32510) );
  and2s1 U23889 ( .DIN1(n31564), .DIN2(n32510), .Q(n31643) );
  and2s1 U23890 ( .DIN1(n31565), .DIN2(u0_csc_mask_r[6]), .Q(n31642) );
  or2s1 U23891 ( .DIN1(n31642), .DIN2(n31643), .Q(n31638) );
  or2s1 U23892 ( .DIN1(n31638), .DIN2(n31639), .Q(n31632) );
  or2s1 U23893 ( .DIN1(n31632), .DIN2(n31633), .Q(n5280) );
  hi1s1 U23894 ( .DIN1(n5280), .Q(n31631) );
  and2s1 U23895 ( .DIN1(n31545), .DIN2(n31631), .Q(n5279) );
  hi1s1 U23896 ( .DIN1(n31102), .Q(n32314) );
  and2s1 U23897 ( .DIN1(n31553), .DIN2(n32314), .Q(n31650) );
  hi1s1 U23898 ( .DIN1(n31103), .Q(n32083) );
  and2s1 U23899 ( .DIN1(n31554), .DIN2(n32083), .Q(n31649) );
  or2s1 U23900 ( .DIN1(n31649), .DIN2(n31650), .Q(n31648) );
  hi1s1 U23901 ( .DIN1(n31104), .Q(n32207) );
  and2s1 U23902 ( .DIN1(n31555), .DIN2(n32207), .Q(n31647) );
  or2s1 U23903 ( .DIN1(n31647), .DIN2(n31648), .Q(n31646) );
  and2s1 U23904 ( .DIN1(n31560), .DIN2(poc_o[7]), .Q(n31654) );
  hi1s1 U23905 ( .DIN1(n31105), .Q(n32410) );
  and2s1 U23906 ( .DIN1(n31561), .DIN2(n32410), .Q(n31653) );
  or2s1 U23907 ( .DIN1(n31653), .DIN2(n31654), .Q(n31652) );
  hi1s1 U23908 ( .DIN1(n31106), .Q(n32507) );
  and2s1 U23909 ( .DIN1(n31564), .DIN2(n32507), .Q(n31656) );
  and2s1 U23910 ( .DIN1(n31565), .DIN2(u0_csc_mask_r[7]), .Q(n31655) );
  or2s1 U23911 ( .DIN1(n31655), .DIN2(n31656), .Q(n31651) );
  or2s1 U23912 ( .DIN1(n31651), .DIN2(n31652), .Q(n31645) );
  or2s1 U23913 ( .DIN1(n31645), .DIN2(n31646), .Q(n5276) );
  hi1s1 U23914 ( .DIN1(n5276), .Q(n31644) );
  and2s1 U23915 ( .DIN1(n31545), .DIN2(n31644), .Q(n5275) );
  hi1s1 U23916 ( .DIN1(n31099), .Q(n32310) );
  and2s1 U23917 ( .DIN1(n31553), .DIN2(n32310), .Q(n31663) );
  and2s1 U23918 ( .DIN1(n31554), .DIN2(u0_csr_r[8]), .Q(n31662) );
  or2s1 U23919 ( .DIN1(n31662), .DIN2(n31663), .Q(n31661) );
  and2s1 U23920 ( .DIN1(n31555), .DIN2(u0_csc0[8]), .Q(n31660) );
  or2s1 U23921 ( .DIN1(n31660), .DIN2(n31661), .Q(n31659) );
  and2s1 U23922 ( .DIN1(n31560), .DIN2(poc_o[8]), .Q(n31667) );
  and2s1 U23923 ( .DIN1(n31561), .DIN2(u0_csc1[8]), .Q(n31666) );
  or2s1 U23924 ( .DIN1(n31666), .DIN2(n31667), .Q(n31665) );
  hi1s1 U23925 ( .DIN1(n31100), .Q(n32504) );
  and2s1 U23926 ( .DIN1(n31564), .DIN2(n32504), .Q(n31669) );
  hi1s1 U23927 ( .DIN1(n31101), .Q(n32121) );
  and2s1 U23928 ( .DIN1(n31565), .DIN2(n32121), .Q(n31668) );
  or2s1 U23929 ( .DIN1(n31668), .DIN2(n31669), .Q(n31664) );
  or2s1 U23930 ( .DIN1(n31664), .DIN2(n31665), .Q(n31658) );
  or2s1 U23931 ( .DIN1(n31658), .DIN2(n31659), .Q(n5272) );
  hi1s1 U23932 ( .DIN1(n5272), .Q(n31657) );
  and2s1 U23933 ( .DIN1(n31545), .DIN2(n31657), .Q(n5271) );
  hi1s1 U23934 ( .DIN1(n31094), .Q(n32306) );
  and2s1 U23935 ( .DIN1(n31553), .DIN2(n32306), .Q(n31676) );
  and2s1 U23936 ( .DIN1(n31554), .DIN2(u0_csr_r[9]), .Q(n31675) );
  or2s1 U23937 ( .DIN1(n31675), .DIN2(n31676), .Q(n31674) );
  hi1s1 U23938 ( .DIN1(n31095), .Q(n32202) );
  and2s1 U23939 ( .DIN1(n31555), .DIN2(n32202), .Q(n31673) );
  or2s1 U23940 ( .DIN1(n31673), .DIN2(n31674), .Q(n31672) );
  and2s1 U23941 ( .DIN1(n31560), .DIN2(poc_o[9]), .Q(n31680) );
  hi1s1 U23942 ( .DIN1(n31096), .Q(n32405) );
  and2s1 U23943 ( .DIN1(n31561), .DIN2(n32405), .Q(n31679) );
  or2s1 U23944 ( .DIN1(n31679), .DIN2(n31680), .Q(n31678) );
  hi1s1 U23945 ( .DIN1(n31097), .Q(n32501) );
  and2s1 U23946 ( .DIN1(n31564), .DIN2(n32501), .Q(n31682) );
  hi1s1 U23947 ( .DIN1(n31098), .Q(n32118) );
  and2s1 U23948 ( .DIN1(n31565), .DIN2(n32118), .Q(n31681) );
  or2s1 U23949 ( .DIN1(n31681), .DIN2(n31682), .Q(n31677) );
  or2s1 U23950 ( .DIN1(n31677), .DIN2(n31678), .Q(n31671) );
  or2s1 U23951 ( .DIN1(n31671), .DIN2(n31672), .Q(n5268) );
  hi1s1 U23952 ( .DIN1(n5268), .Q(n31670) );
  and2s1 U23953 ( .DIN1(n31545), .DIN2(n31670), .Q(n5267) );
  hi1s1 U23954 ( .DIN1(n31089), .Q(n32302) );
  and2s1 U23955 ( .DIN1(n31553), .DIN2(n32302), .Q(n31689) );
  and2s1 U23956 ( .DIN1(n31554), .DIN2(u0_csr_r[10]), .Q(n31688) );
  or2s1 U23957 ( .DIN1(n31688), .DIN2(n31689), .Q(n31687) );
  hi1s1 U23958 ( .DIN1(n31090), .Q(n32199) );
  and2s1 U23959 ( .DIN1(n31555), .DIN2(n32199), .Q(n31686) );
  or2s1 U23960 ( .DIN1(n31686), .DIN2(n31687), .Q(n31685) );
  and2s1 U23961 ( .DIN1(n31560), .DIN2(poc_o[10]), .Q(n31693) );
  hi1s1 U23962 ( .DIN1(n31091), .Q(n32402) );
  and2s1 U23963 ( .DIN1(n31561), .DIN2(n32402), .Q(n31692) );
  or2s1 U23964 ( .DIN1(n31692), .DIN2(n31693), .Q(n31691) );
  hi1s1 U23965 ( .DIN1(n31092), .Q(n32498) );
  and2s1 U23966 ( .DIN1(n31564), .DIN2(n32498), .Q(n31695) );
  hi1s1 U23967 ( .DIN1(n31093), .Q(n32114) );
  and2s1 U23968 ( .DIN1(n31565), .DIN2(n32114), .Q(n31694) );
  or2s1 U23969 ( .DIN1(n31694), .DIN2(n31695), .Q(n31690) );
  or2s1 U23970 ( .DIN1(n31690), .DIN2(n31691), .Q(n31684) );
  or2s1 U23971 ( .DIN1(n31684), .DIN2(n31685), .Q(n5264) );
  hi1s1 U23972 ( .DIN1(n5264), .Q(n31683) );
  and2s1 U23973 ( .DIN1(n31545), .DIN2(n31683), .Q(n5263) );
  hi1s1 U23974 ( .DIN1(n31085), .Q(n32196) );
  and2s1 U23975 ( .DIN1(n31555), .DIN2(n32196), .Q(n31700) );
  hi1s1 U23976 ( .DIN1(n31086), .Q(n32298) );
  and2s1 U23977 ( .DIN1(n31553), .DIN2(n32298), .Q(n31699) );
  or2s1 U23978 ( .DIN1(n31699), .DIN2(n31700), .Q(n31698) );
  hi1s1 U23979 ( .DIN1(n31087), .Q(n32399) );
  and2s1 U23980 ( .DIN1(n31561), .DIN2(n32399), .Q(n31704) );
  hi1s1 U23981 ( .DIN1(n31088), .Q(n32495) );
  and2s1 U23982 ( .DIN1(n31564), .DIN2(n32495), .Q(n31703) );
  or2s1 U23983 ( .DIN1(n31703), .DIN2(n31704), .Q(n31702) );
  and2s1 U23984 ( .DIN1(n31560), .DIN2(poc_o[11]), .Q(n31701) );
  or2s1 U23985 ( .DIN1(n31701), .DIN2(n31702), .Q(n31697) );
  or2s1 U23986 ( .DIN1(n31697), .DIN2(n31698), .Q(n5260) );
  hi1s1 U23987 ( .DIN1(n5260), .Q(n31696) );
  and2s1 U23988 ( .DIN1(n31545), .DIN2(n31696), .Q(n5259) );
  hi1s1 U23989 ( .DIN1(n31081), .Q(n32193) );
  and2s1 U23990 ( .DIN1(n31555), .DIN2(n32193), .Q(n31709) );
  hi1s1 U23991 ( .DIN1(n31082), .Q(n32294) );
  and2s1 U23992 ( .DIN1(n31553), .DIN2(n32294), .Q(n31708) );
  or2s1 U23993 ( .DIN1(n31708), .DIN2(n31709), .Q(n31707) );
  hi1s1 U23994 ( .DIN1(n31083), .Q(n32396) );
  and2s1 U23995 ( .DIN1(n31561), .DIN2(n32396), .Q(n31713) );
  hi1s1 U23996 ( .DIN1(n31084), .Q(n32492) );
  and2s1 U23997 ( .DIN1(n31564), .DIN2(n32492), .Q(n31712) );
  or2s1 U23998 ( .DIN1(n31712), .DIN2(n31713), .Q(n31711) );
  and2s1 U23999 ( .DIN1(n31560), .DIN2(poc_o[12]), .Q(n31710) );
  or2s1 U24000 ( .DIN1(n31710), .DIN2(n31711), .Q(n31706) );
  or2s1 U24001 ( .DIN1(n31706), .DIN2(n31707), .Q(n5256) );
  hi1s1 U24002 ( .DIN1(n5256), .Q(n31705) );
  and2s1 U24003 ( .DIN1(n31545), .DIN2(n31705), .Q(n5255) );
  hi1s1 U24004 ( .DIN1(n31077), .Q(n32190) );
  and2s1 U24005 ( .DIN1(n31555), .DIN2(n32190), .Q(n31718) );
  hi1s1 U24006 ( .DIN1(n31078), .Q(n32290) );
  and2s1 U24007 ( .DIN1(n31553), .DIN2(n32290), .Q(n31717) );
  or2s1 U24008 ( .DIN1(n31717), .DIN2(n31718), .Q(n31716) );
  hi1s1 U24009 ( .DIN1(n31079), .Q(n32393) );
  and2s1 U24010 ( .DIN1(n31561), .DIN2(n32393), .Q(n31722) );
  hi1s1 U24011 ( .DIN1(n31080), .Q(n32489) );
  and2s1 U24012 ( .DIN1(n31564), .DIN2(n32489), .Q(n31721) );
  or2s1 U24013 ( .DIN1(n31721), .DIN2(n31722), .Q(n31720) );
  and2s1 U24014 ( .DIN1(n31560), .DIN2(poc_o[13]), .Q(n31719) );
  or2s1 U24015 ( .DIN1(n31719), .DIN2(n31720), .Q(n31715) );
  or2s1 U24016 ( .DIN1(n31715), .DIN2(n31716), .Q(n5252) );
  hi1s1 U24017 ( .DIN1(n5252), .Q(n31714) );
  and2s1 U24018 ( .DIN1(n31545), .DIN2(n31714), .Q(n5251) );
  hi1s1 U24019 ( .DIN1(n31073), .Q(n32187) );
  and2s1 U24020 ( .DIN1(n31555), .DIN2(n32187), .Q(n31727) );
  hi1s1 U24021 ( .DIN1(n31074), .Q(n32286) );
  and2s1 U24022 ( .DIN1(n31553), .DIN2(n32286), .Q(n31726) );
  or2s1 U24023 ( .DIN1(n31726), .DIN2(n31727), .Q(n31725) );
  hi1s1 U24024 ( .DIN1(n31075), .Q(n32390) );
  and2s1 U24025 ( .DIN1(n31561), .DIN2(n32390), .Q(n31731) );
  hi1s1 U24026 ( .DIN1(n31076), .Q(n32486) );
  and2s1 U24027 ( .DIN1(n31564), .DIN2(n32486), .Q(n31730) );
  or2s1 U24028 ( .DIN1(n31730), .DIN2(n31731), .Q(n31729) );
  and2s1 U24029 ( .DIN1(n31560), .DIN2(poc_o[14]), .Q(n31728) );
  or2s1 U24030 ( .DIN1(n31728), .DIN2(n31729), .Q(n31724) );
  or2s1 U24031 ( .DIN1(n31724), .DIN2(n31725), .Q(n5248) );
  hi1s1 U24032 ( .DIN1(n5248), .Q(n31723) );
  and2s1 U24033 ( .DIN1(n31545), .DIN2(n31723), .Q(n5247) );
  hi1s1 U24034 ( .DIN1(n31069), .Q(n32184) );
  and2s1 U24035 ( .DIN1(n31555), .DIN2(n32184), .Q(n31736) );
  hi1s1 U24036 ( .DIN1(n31070), .Q(n32282) );
  and2s1 U24037 ( .DIN1(n31553), .DIN2(n32282), .Q(n31735) );
  or2s1 U24038 ( .DIN1(n31735), .DIN2(n31736), .Q(n31734) );
  hi1s1 U24039 ( .DIN1(n31071), .Q(n32387) );
  and2s1 U24040 ( .DIN1(n31561), .DIN2(n32387), .Q(n31740) );
  hi1s1 U24041 ( .DIN1(n31072), .Q(n32483) );
  and2s1 U24042 ( .DIN1(n31564), .DIN2(n32483), .Q(n31739) );
  or2s1 U24043 ( .DIN1(n31739), .DIN2(n31740), .Q(n31738) );
  and2s1 U24044 ( .DIN1(n31560), .DIN2(poc_o[15]), .Q(n31737) );
  or2s1 U24045 ( .DIN1(n31737), .DIN2(n31738), .Q(n31733) );
  or2s1 U24046 ( .DIN1(n31733), .DIN2(n31734), .Q(n5244) );
  hi1s1 U24047 ( .DIN1(n5244), .Q(n31732) );
  and2s1 U24048 ( .DIN1(n31545), .DIN2(n31732), .Q(n5243) );
  and2s1 U24049 ( .DIN1(n31555), .DIN2(u0_csc0[16]), .Q(n31745) );
  hi1s1 U24050 ( .DIN1(n31067), .Q(n32278) );
  and2s1 U24051 ( .DIN1(n31553), .DIN2(n32278), .Q(n31744) );
  or2s1 U24052 ( .DIN1(n31744), .DIN2(n31745), .Q(n31743) );
  and2s1 U24053 ( .DIN1(n31561), .DIN2(u0_csc1[16]), .Q(n31749) );
  hi1s1 U24054 ( .DIN1(n31068), .Q(n32480) );
  and2s1 U24055 ( .DIN1(n31564), .DIN2(n32480), .Q(n31748) );
  or2s1 U24056 ( .DIN1(n31748), .DIN2(n31749), .Q(n31747) );
  and2s1 U24057 ( .DIN1(n31560), .DIN2(poc_o[16]), .Q(n31746) );
  or2s1 U24058 ( .DIN1(n31746), .DIN2(n31747), .Q(n31742) );
  or2s1 U24059 ( .DIN1(n31742), .DIN2(n31743), .Q(n5240) );
  hi1s1 U24060 ( .DIN1(n5240), .Q(n31741) );
  and2s1 U24061 ( .DIN1(n31545), .DIN2(n31741), .Q(n5239) );
  and2s1 U24062 ( .DIN1(n31555), .DIN2(u0_csc0[17]), .Q(n31754) );
  hi1s1 U24063 ( .DIN1(n31065), .Q(n32274) );
  and2s1 U24064 ( .DIN1(n31553), .DIN2(n32274), .Q(n31753) );
  or2s1 U24065 ( .DIN1(n31753), .DIN2(n31754), .Q(n31752) );
  and2s1 U24066 ( .DIN1(n31561), .DIN2(u0_csc1[17]), .Q(n31758) );
  hi1s1 U24067 ( .DIN1(n31066), .Q(n32477) );
  and2s1 U24068 ( .DIN1(n31564), .DIN2(n32477), .Q(n31757) );
  or2s1 U24069 ( .DIN1(n31757), .DIN2(n31758), .Q(n31756) );
  and2s1 U24070 ( .DIN1(n31560), .DIN2(poc_o[17]), .Q(n31755) );
  or2s1 U24071 ( .DIN1(n31755), .DIN2(n31756), .Q(n31751) );
  or2s1 U24072 ( .DIN1(n31751), .DIN2(n31752), .Q(n5236) );
  hi1s1 U24073 ( .DIN1(n5236), .Q(n31750) );
  and2s1 U24074 ( .DIN1(n31545), .DIN2(n31750), .Q(n5235) );
  and2s1 U24075 ( .DIN1(n31555), .DIN2(u0_csc0[18]), .Q(n31763) );
  hi1s1 U24076 ( .DIN1(n31063), .Q(n32270) );
  and2s1 U24077 ( .DIN1(n31553), .DIN2(n32270), .Q(n31762) );
  or2s1 U24078 ( .DIN1(n31762), .DIN2(n31763), .Q(n31761) );
  and2s1 U24079 ( .DIN1(n31561), .DIN2(u0_csc1[18]), .Q(n31767) );
  hi1s1 U24080 ( .DIN1(n31064), .Q(n32474) );
  and2s1 U24081 ( .DIN1(n31564), .DIN2(n32474), .Q(n31766) );
  or2s1 U24082 ( .DIN1(n31766), .DIN2(n31767), .Q(n31765) );
  and2s1 U24083 ( .DIN1(n31560), .DIN2(poc_o[18]), .Q(n31764) );
  or2s1 U24084 ( .DIN1(n31764), .DIN2(n31765), .Q(n31760) );
  or2s1 U24085 ( .DIN1(n31760), .DIN2(n31761), .Q(n5232) );
  hi1s1 U24086 ( .DIN1(n5232), .Q(n31759) );
  and2s1 U24087 ( .DIN1(n31545), .DIN2(n31759), .Q(n5231) );
  and2s1 U24088 ( .DIN1(n31555), .DIN2(u0_csc0[19]), .Q(n31772) );
  hi1s1 U24089 ( .DIN1(n31061), .Q(n32266) );
  and2s1 U24090 ( .DIN1(n31553), .DIN2(n32266), .Q(n31771) );
  or2s1 U24091 ( .DIN1(n31771), .DIN2(n31772), .Q(n31770) );
  and2s1 U24092 ( .DIN1(n31561), .DIN2(u0_csc1[19]), .Q(n31776) );
  hi1s1 U24093 ( .DIN1(n31062), .Q(n32471) );
  and2s1 U24094 ( .DIN1(n31564), .DIN2(n32471), .Q(n31775) );
  or2s1 U24095 ( .DIN1(n31775), .DIN2(n31776), .Q(n31774) );
  and2s1 U24096 ( .DIN1(n31560), .DIN2(poc_o[19]), .Q(n31773) );
  or2s1 U24097 ( .DIN1(n31773), .DIN2(n31774), .Q(n31769) );
  or2s1 U24098 ( .DIN1(n31769), .DIN2(n31770), .Q(n5228) );
  hi1s1 U24099 ( .DIN1(n5228), .Q(n31768) );
  and2s1 U24100 ( .DIN1(n31545), .DIN2(n31768), .Q(n5227) );
  and2s1 U24101 ( .DIN1(n31555), .DIN2(u0_csc0[20]), .Q(n31781) );
  hi1s1 U24102 ( .DIN1(n31059), .Q(n32262) );
  and2s1 U24103 ( .DIN1(n31553), .DIN2(n32262), .Q(n31780) );
  or2s1 U24104 ( .DIN1(n31780), .DIN2(n31781), .Q(n31779) );
  and2s1 U24105 ( .DIN1(n31561), .DIN2(u0_csc1[20]), .Q(n31785) );
  hi1s1 U24106 ( .DIN1(n31060), .Q(n32468) );
  and2s1 U24107 ( .DIN1(n31564), .DIN2(n32468), .Q(n31784) );
  or2s1 U24108 ( .DIN1(n31784), .DIN2(n31785), .Q(n31783) );
  and2s1 U24109 ( .DIN1(n31560), .DIN2(poc_o[20]), .Q(n31782) );
  or2s1 U24110 ( .DIN1(n31782), .DIN2(n31783), .Q(n31778) );
  or2s1 U24111 ( .DIN1(n31778), .DIN2(n31779), .Q(n5224) );
  hi1s1 U24112 ( .DIN1(n5224), .Q(n31777) );
  and2s1 U24113 ( .DIN1(n31545), .DIN2(n31777), .Q(n5223) );
  and2s1 U24114 ( .DIN1(n31555), .DIN2(u0_csc0[21]), .Q(n31790) );
  hi1s1 U24115 ( .DIN1(n31057), .Q(n32258) );
  and2s1 U24116 ( .DIN1(n31553), .DIN2(n32258), .Q(n31789) );
  or2s1 U24117 ( .DIN1(n31789), .DIN2(n31790), .Q(n31788) );
  and2s1 U24118 ( .DIN1(n31561), .DIN2(u0_csc1[21]), .Q(n31794) );
  hi1s1 U24119 ( .DIN1(n31058), .Q(n32465) );
  and2s1 U24120 ( .DIN1(n31564), .DIN2(n32465), .Q(n31793) );
  or2s1 U24121 ( .DIN1(n31793), .DIN2(n31794), .Q(n31792) );
  and2s1 U24122 ( .DIN1(n31560), .DIN2(poc_o[21]), .Q(n31791) );
  or2s1 U24123 ( .DIN1(n31791), .DIN2(n31792), .Q(n31787) );
  or2s1 U24124 ( .DIN1(n31787), .DIN2(n31788), .Q(n5220) );
  hi1s1 U24125 ( .DIN1(n5220), .Q(n31786) );
  and2s1 U24126 ( .DIN1(n31545), .DIN2(n31786), .Q(n5219) );
  and2s1 U24127 ( .DIN1(n31555), .DIN2(u0_csc0[22]), .Q(n31799) );
  hi1s1 U24128 ( .DIN1(n31055), .Q(n32254) );
  and2s1 U24129 ( .DIN1(n31553), .DIN2(n32254), .Q(n31798) );
  or2s1 U24130 ( .DIN1(n31798), .DIN2(n31799), .Q(n31797) );
  and2s1 U24131 ( .DIN1(n31561), .DIN2(u0_csc1[22]), .Q(n31803) );
  hi1s1 U24132 ( .DIN1(n31056), .Q(n32462) );
  and2s1 U24133 ( .DIN1(n31564), .DIN2(n32462), .Q(n31802) );
  or2s1 U24134 ( .DIN1(n31802), .DIN2(n31803), .Q(n31801) );
  and2s1 U24135 ( .DIN1(n31560), .DIN2(poc_o[22]), .Q(n31800) );
  or2s1 U24136 ( .DIN1(n31800), .DIN2(n31801), .Q(n31796) );
  or2s1 U24137 ( .DIN1(n31796), .DIN2(n31797), .Q(n5216) );
  hi1s1 U24138 ( .DIN1(n5216), .Q(n31795) );
  and2s1 U24139 ( .DIN1(n31545), .DIN2(n31795), .Q(n5215) );
  and2s1 U24140 ( .DIN1(n31555), .DIN2(u0_csc0[23]), .Q(n31808) );
  hi1s1 U24141 ( .DIN1(n31053), .Q(n32250) );
  and2s1 U24142 ( .DIN1(n31553), .DIN2(n32250), .Q(n31807) );
  or2s1 U24143 ( .DIN1(n31807), .DIN2(n31808), .Q(n31806) );
  and2s1 U24144 ( .DIN1(n31561), .DIN2(u0_csc1[23]), .Q(n31812) );
  hi1s1 U24145 ( .DIN1(n31054), .Q(n32459) );
  and2s1 U24146 ( .DIN1(n31564), .DIN2(n32459), .Q(n31811) );
  or2s1 U24147 ( .DIN1(n31811), .DIN2(n31812), .Q(n31810) );
  and2s1 U24148 ( .DIN1(n31560), .DIN2(poc_o[23]), .Q(n31809) );
  or2s1 U24149 ( .DIN1(n31809), .DIN2(n31810), .Q(n31805) );
  or2s1 U24150 ( .DIN1(n31805), .DIN2(n31806), .Q(n5212) );
  hi1s1 U24151 ( .DIN1(n5212), .Q(n31804) );
  and2s1 U24152 ( .DIN1(n31545), .DIN2(n31804), .Q(n5211) );
  hi1s1 U24153 ( .DIN1(n31049), .Q(n32246) );
  and2s1 U24154 ( .DIN1(n31553), .DIN2(n32246), .Q(n31819) );
  and2s1 U24155 ( .DIN1(n31554), .DIN2(u0_csr_r2[0]), .Q(n31818) );
  or2s1 U24156 ( .DIN1(n31818), .DIN2(n31819), .Q(n31817) );
  hi1s1 U24157 ( .DIN1(n31050), .Q(n32165) );
  and2s1 U24158 ( .DIN1(n31555), .DIN2(n32165), .Q(n31816) );
  or2s1 U24159 ( .DIN1(n31816), .DIN2(n31817), .Q(n31815) );
  hi1s1 U24160 ( .DIN1(n31051), .Q(n32368) );
  and2s1 U24161 ( .DIN1(n31561), .DIN2(n32368), .Q(n31823) );
  hi1s1 U24162 ( .DIN1(n31052), .Q(n32456) );
  and2s1 U24163 ( .DIN1(n31564), .DIN2(n32456), .Q(n31822) );
  or2s1 U24164 ( .DIN1(n31822), .DIN2(n31823), .Q(n31821) );
  and2s1 U24165 ( .DIN1(n31560), .DIN2(poc_o[24]), .Q(n31820) );
  or2s1 U24166 ( .DIN1(n31820), .DIN2(n31821), .Q(n31814) );
  or2s1 U24167 ( .DIN1(n31814), .DIN2(n31815), .Q(n5208) );
  hi1s1 U24168 ( .DIN1(n5208), .Q(n31813) );
  and2s1 U24169 ( .DIN1(n31545), .DIN2(n31813), .Q(n5207) );
  hi1s1 U24170 ( .DIN1(n31045), .Q(n32242) );
  and2s1 U24171 ( .DIN1(n31553), .DIN2(n32242), .Q(n31830) );
  and2s1 U24172 ( .DIN1(n31554), .DIN2(u0_csr_r2[1]), .Q(n31829) );
  or2s1 U24173 ( .DIN1(n31829), .DIN2(n31830), .Q(n31828) );
  hi1s1 U24174 ( .DIN1(n31046), .Q(n32162) );
  and2s1 U24175 ( .DIN1(n31555), .DIN2(n32162), .Q(n31827) );
  or2s1 U24176 ( .DIN1(n31827), .DIN2(n31828), .Q(n31826) );
  hi1s1 U24177 ( .DIN1(n31047), .Q(n32365) );
  and2s1 U24178 ( .DIN1(n31561), .DIN2(n32365), .Q(n31834) );
  hi1s1 U24179 ( .DIN1(n31048), .Q(n32453) );
  and2s1 U24180 ( .DIN1(n31564), .DIN2(n32453), .Q(n31833) );
  or2s1 U24181 ( .DIN1(n31833), .DIN2(n31834), .Q(n31832) );
  and2s1 U24182 ( .DIN1(n31560), .DIN2(poc_o[25]), .Q(n31831) );
  or2s1 U24183 ( .DIN1(n31831), .DIN2(n31832), .Q(n31825) );
  or2s1 U24184 ( .DIN1(n31825), .DIN2(n31826), .Q(n5204) );
  hi1s1 U24185 ( .DIN1(n5204), .Q(n31824) );
  and2s1 U24186 ( .DIN1(n31545), .DIN2(n31824), .Q(n5203) );
  hi1s1 U24187 ( .DIN1(n31041), .Q(n32238) );
  and2s1 U24188 ( .DIN1(n31553), .DIN2(n32238), .Q(n31841) );
  and2s1 U24189 ( .DIN1(n31554), .DIN2(u0_csr_r2[2]), .Q(n31840) );
  or2s1 U24190 ( .DIN1(n31840), .DIN2(n31841), .Q(n31839) );
  hi1s1 U24191 ( .DIN1(n31042), .Q(n32159) );
  and2s1 U24192 ( .DIN1(n31555), .DIN2(n32159), .Q(n31838) );
  or2s1 U24193 ( .DIN1(n31838), .DIN2(n31839), .Q(n31837) );
  hi1s1 U24194 ( .DIN1(n31043), .Q(n32362) );
  and2s1 U24195 ( .DIN1(n31561), .DIN2(n32362), .Q(n31845) );
  hi1s1 U24196 ( .DIN1(n31044), .Q(n32450) );
  and2s1 U24197 ( .DIN1(n31564), .DIN2(n32450), .Q(n31844) );
  or2s1 U24198 ( .DIN1(n31844), .DIN2(n31845), .Q(n31843) );
  and2s1 U24199 ( .DIN1(n31560), .DIN2(poc_o[26]), .Q(n31842) );
  or2s1 U24200 ( .DIN1(n31842), .DIN2(n31843), .Q(n31836) );
  or2s1 U24201 ( .DIN1(n31836), .DIN2(n31837), .Q(n5200) );
  hi1s1 U24202 ( .DIN1(n5200), .Q(n31835) );
  and2s1 U24203 ( .DIN1(n31545), .DIN2(n31835), .Q(n5199) );
  hi1s1 U24204 ( .DIN1(n31037), .Q(n32234) );
  and2s1 U24205 ( .DIN1(n31553), .DIN2(n32234), .Q(n31852) );
  and2s1 U24206 ( .DIN1(n31554), .DIN2(u0_csr_r2[3]), .Q(n31851) );
  or2s1 U24207 ( .DIN1(n31851), .DIN2(n31852), .Q(n31850) );
  hi1s1 U24208 ( .DIN1(n31038), .Q(n32156) );
  and2s1 U24209 ( .DIN1(n31555), .DIN2(n32156), .Q(n31849) );
  or2s1 U24210 ( .DIN1(n31849), .DIN2(n31850), .Q(n31848) );
  hi1s1 U24211 ( .DIN1(n31039), .Q(n32359) );
  and2s1 U24212 ( .DIN1(n31561), .DIN2(n32359), .Q(n31856) );
  hi1s1 U24213 ( .DIN1(n31040), .Q(n32447) );
  and2s1 U24214 ( .DIN1(n31564), .DIN2(n32447), .Q(n31855) );
  or2s1 U24215 ( .DIN1(n31855), .DIN2(n31856), .Q(n31854) );
  and2s1 U24216 ( .DIN1(n31560), .DIN2(poc_o[27]), .Q(n31853) );
  or2s1 U24217 ( .DIN1(n31853), .DIN2(n31854), .Q(n31847) );
  or2s1 U24218 ( .DIN1(n31847), .DIN2(n31848), .Q(n5196) );
  hi1s1 U24219 ( .DIN1(n5196), .Q(n31846) );
  and2s1 U24220 ( .DIN1(n31545), .DIN2(n31846), .Q(n5195) );
  hi1s1 U24221 ( .DIN1(n31033), .Q(n32230) );
  and2s1 U24222 ( .DIN1(n31553), .DIN2(n32230), .Q(n31863) );
  and2s1 U24223 ( .DIN1(n31554), .DIN2(u0_csr_r2[4]), .Q(n31862) );
  or2s1 U24224 ( .DIN1(n31862), .DIN2(n31863), .Q(n31861) );
  hi1s1 U24225 ( .DIN1(n31034), .Q(n32153) );
  and2s1 U24226 ( .DIN1(n31555), .DIN2(n32153), .Q(n31860) );
  or2s1 U24227 ( .DIN1(n31860), .DIN2(n31861), .Q(n31859) );
  hi1s1 U24228 ( .DIN1(n31035), .Q(n32356) );
  and2s1 U24229 ( .DIN1(n31561), .DIN2(n32356), .Q(n31867) );
  hi1s1 U24230 ( .DIN1(n31036), .Q(n32444) );
  and2s1 U24231 ( .DIN1(n31564), .DIN2(n32444), .Q(n31866) );
  or2s1 U24232 ( .DIN1(n31866), .DIN2(n31867), .Q(n31865) );
  and2s1 U24233 ( .DIN1(n31560), .DIN2(poc_o[28]), .Q(n31864) );
  or2s1 U24234 ( .DIN1(n31864), .DIN2(n31865), .Q(n31858) );
  or2s1 U24235 ( .DIN1(n31858), .DIN2(n31859), .Q(n5192) );
  hi1s1 U24236 ( .DIN1(n5192), .Q(n31857) );
  and2s1 U24237 ( .DIN1(n31545), .DIN2(n31857), .Q(n5191) );
  hi1s1 U24238 ( .DIN1(n31029), .Q(n32226) );
  and2s1 U24239 ( .DIN1(n31553), .DIN2(n32226), .Q(n31874) );
  and2s1 U24240 ( .DIN1(n31554), .DIN2(u0_csr_r2[5]), .Q(n31873) );
  or2s1 U24241 ( .DIN1(n31873), .DIN2(n31874), .Q(n31872) );
  hi1s1 U24242 ( .DIN1(n31030), .Q(n32150) );
  and2s1 U24243 ( .DIN1(n31555), .DIN2(n32150), .Q(n31871) );
  or2s1 U24244 ( .DIN1(n31871), .DIN2(n31872), .Q(n31870) );
  hi1s1 U24245 ( .DIN1(n31031), .Q(n32353) );
  and2s1 U24246 ( .DIN1(n31561), .DIN2(n32353), .Q(n31878) );
  hi1s1 U24247 ( .DIN1(n31032), .Q(n32441) );
  and2s1 U24248 ( .DIN1(n31564), .DIN2(n32441), .Q(n31877) );
  or2s1 U24249 ( .DIN1(n31877), .DIN2(n31878), .Q(n31876) );
  and2s1 U24250 ( .DIN1(n31560), .DIN2(poc_o[29]), .Q(n31875) );
  or2s1 U24251 ( .DIN1(n31875), .DIN2(n31876), .Q(n31869) );
  or2s1 U24252 ( .DIN1(n31869), .DIN2(n31870), .Q(n5188) );
  hi1s1 U24253 ( .DIN1(n5188), .Q(n31868) );
  and2s1 U24254 ( .DIN1(n31545), .DIN2(n31868), .Q(n5187) );
  hi1s1 U24255 ( .DIN1(n31025), .Q(n32222) );
  and2s1 U24256 ( .DIN1(n31553), .DIN2(n32222), .Q(n31885) );
  and2s1 U24257 ( .DIN1(n31554), .DIN2(u0_csr_r2[6]), .Q(n31884) );
  or2s1 U24258 ( .DIN1(n31884), .DIN2(n31885), .Q(n31883) );
  hi1s1 U24259 ( .DIN1(n31026), .Q(n32147) );
  and2s1 U24260 ( .DIN1(n31555), .DIN2(n32147), .Q(n31882) );
  or2s1 U24261 ( .DIN1(n31882), .DIN2(n31883), .Q(n31881) );
  hi1s1 U24262 ( .DIN1(n31027), .Q(n32350) );
  and2s1 U24263 ( .DIN1(n31561), .DIN2(n32350), .Q(n31889) );
  hi1s1 U24264 ( .DIN1(n31028), .Q(n32438) );
  and2s1 U24265 ( .DIN1(n31564), .DIN2(n32438), .Q(n31888) );
  or2s1 U24266 ( .DIN1(n31888), .DIN2(n31889), .Q(n31887) );
  and2s1 U24267 ( .DIN1(n31560), .DIN2(poc_o[30]), .Q(n31886) );
  or2s1 U24268 ( .DIN1(n31886), .DIN2(n31887), .Q(n31880) );
  or2s1 U24269 ( .DIN1(n31880), .DIN2(n31881), .Q(n5184) );
  hi1s1 U24270 ( .DIN1(n5184), .Q(n31879) );
  and2s1 U24271 ( .DIN1(n31545), .DIN2(n31879), .Q(n5183) );
  hi1s1 U24272 ( .DIN1(n31021), .Q(n32218) );
  and2s1 U24273 ( .DIN1(n31553), .DIN2(n32218), .Q(n31896) );
  and2s1 U24274 ( .DIN1(n31554), .DIN2(u0_csr_r2[7]), .Q(n31895) );
  or2s1 U24275 ( .DIN1(n31895), .DIN2(n31896), .Q(n31894) );
  hi1s1 U24276 ( .DIN1(n31022), .Q(n32144) );
  and2s1 U24277 ( .DIN1(n31555), .DIN2(n32144), .Q(n31893) );
  or2s1 U24278 ( .DIN1(n31893), .DIN2(n31894), .Q(n31892) );
  hi1s1 U24279 ( .DIN1(n31023), .Q(n32347) );
  and2s1 U24280 ( .DIN1(n31561), .DIN2(n32347), .Q(n31900) );
  hi1s1 U24281 ( .DIN1(n31024), .Q(n32435) );
  and2s1 U24282 ( .DIN1(n31564), .DIN2(n32435), .Q(n31899) );
  or2s1 U24283 ( .DIN1(n31899), .DIN2(n31900), .Q(n31898) );
  and2s1 U24284 ( .DIN1(n31560), .DIN2(poc_o[31]), .Q(n31897) );
  or2s1 U24285 ( .DIN1(n31897), .DIN2(n31898), .Q(n31891) );
  or2s1 U24286 ( .DIN1(n31891), .DIN2(n31892), .Q(n5180) );
  hi1s1 U24287 ( .DIN1(n5180), .Q(n31890) );
  and2s1 U24288 ( .DIN1(wb_addr_i[5]), .DIN2(n31907), .Q(n31906) );
  hi1s1 U24289 ( .DIN1(wb_addr_i[6]), .Q(n31907) );
  or2s1 U24290 ( .DIN1(wb_addr_i[4]), .DIN2(wb_addr_i[5]), .Q(n31909) );
  or2s1 U24291 ( .DIN1(n31909), .DIN2(n31907), .Q(n31908) );
  hi1s1 U24292 ( .DIN1(n31908), .Q(n31905) );
  or2s1 U24293 ( .DIN1(n31905), .DIN2(n31906), .Q(n31904) );
  or2s1 U24294 ( .DIN1(n31911), .DIN2(n31912), .Q(n31910) );
  hi1s1 U24295 ( .DIN1(n31910), .Q(n31565) );
  or2s1 U24296 ( .DIN1(n31916), .DIN2(n31917), .Q(n31915) );
  or2s1 U24297 ( .DIN1(n31914), .DIN2(n31915), .Q(n31913) );
  hi1s1 U24298 ( .DIN1(n31913), .Q(n31564) );
  or2s1 U24299 ( .DIN1(n31564), .DIN2(n31565), .Q(n31903) );
  or2s1 U24300 ( .DIN1(n31903), .DIN2(n31904), .Q(n31902) );
  hi1s1 U24301 ( .DIN1(wb_addr_i[3]), .Q(n31916) );
  or2s1 U24302 ( .DIN1(wb_addr_i[2]), .DIN2(n31916), .Q(n31912) );
  or2s1 U24303 ( .DIN1(n31914), .DIN2(n31912), .Q(n31920) );
  hi1s1 U24304 ( .DIN1(n31920), .Q(n31561) );
  or2s1 U24305 ( .DIN1(n31911), .DIN2(n31922), .Q(n31921) );
  hi1s1 U24306 ( .DIN1(n31921), .Q(n31560) );
  or2s1 U24307 ( .DIN1(n31560), .DIN2(n31561), .Q(n31919) );
  hi1s1 U24308 ( .DIN1(wb_addr_i[2]), .Q(n31917) );
  or2s1 U24309 ( .DIN1(wb_addr_i[3]), .DIN2(n31917), .Q(n31922) );
  or2s1 U24310 ( .DIN1(n31914), .DIN2(n31922), .Q(n31924) );
  hi1s1 U24311 ( .DIN1(n31924), .Q(n31553) );
  hi1s1 U24312 ( .DIN1(wb_addr_i[4]), .Q(n31927) );
  or2s1 U24313 ( .DIN1(n31927), .DIN2(n31928), .Q(n31914) );
  or2s1 U24314 ( .DIN1(n31914), .DIN2(n31926), .Q(n31925) );
  hi1s1 U24315 ( .DIN1(n31925), .Q(n31555) );
  or2s1 U24316 ( .DIN1(n31555), .DIN2(n31553), .Q(n31923) );
  or2s1 U24317 ( .DIN1(wb_addr_i[3]), .DIN2(wb_addr_i[2]), .Q(n31926) );
  or2s1 U24318 ( .DIN1(wb_addr_i[6]), .DIN2(wb_addr_i[5]), .Q(n31928) );
  or2s1 U24319 ( .DIN1(wb_addr_i[4]), .DIN2(n31928), .Q(n31911) );
  or2s1 U24320 ( .DIN1(n31911), .DIN2(n31926), .Q(n31929) );
  hi1s1 U24321 ( .DIN1(n31929), .Q(n31554) );
  or2s1 U24322 ( .DIN1(n31554), .DIN2(n31923), .Q(n31918) );
  or2s1 U24323 ( .DIN1(n31918), .DIN2(n31919), .Q(n31901) );
  or2s1 U24324 ( .DIN1(n31901), .DIN2(n31902), .Q(n31545) );
  and2s1 U24325 ( .DIN1(n31545), .DIN2(n31890), .Q(n5179) );
  and2s1 U24326 ( .DIN1(n32029), .DIN2(n32030), .Q(n9963) );
  and2s1 U24327 ( .DIN1(n32031), .DIN2(n32032), .Q(n32030) );
  and2s1 U24328 ( .DIN1(n32033), .DIN2(n32034), .Q(n32031) );
  or2s1 U24329 ( .DIN1(n32035), .DIN2(n32036), .Q(n9962) );
  and2s1 U24330 ( .DIN1(u0_csr_r2[7]), .DIN2(n32037), .Q(n32036) );
  and2s1 U24331 ( .DIN1(wb_data_i[31]), .DIN2(n32038), .Q(n32035) );
  or2s1 U24332 ( .DIN1(n32039), .DIN2(n32040), .Q(n9961) );
  and2s1 U24333 ( .DIN1(u0_csr_r2[6]), .DIN2(n32037), .Q(n32040) );
  and2s1 U24334 ( .DIN1(wb_data_i[30]), .DIN2(n32038), .Q(n32039) );
  or2s1 U24335 ( .DIN1(n32041), .DIN2(n32042), .Q(n9960) );
  and2s1 U24336 ( .DIN1(u0_csr_r2[5]), .DIN2(n32037), .Q(n32042) );
  and2s1 U24337 ( .DIN1(wb_data_i[29]), .DIN2(n32038), .Q(n32041) );
  or2s1 U24338 ( .DIN1(n32043), .DIN2(n32044), .Q(n9959) );
  and2s1 U24339 ( .DIN1(u0_csr_r2[4]), .DIN2(n32037), .Q(n32044) );
  and2s1 U24340 ( .DIN1(wb_data_i[28]), .DIN2(n32038), .Q(n32043) );
  or2s1 U24341 ( .DIN1(n32045), .DIN2(n32046), .Q(n9958) );
  and2s1 U24342 ( .DIN1(u0_csr_r2[3]), .DIN2(n32037), .Q(n32046) );
  and2s1 U24343 ( .DIN1(wb_data_i[27]), .DIN2(n32038), .Q(n32045) );
  or2s1 U24344 ( .DIN1(n32047), .DIN2(n32048), .Q(n9957) );
  and2s1 U24345 ( .DIN1(u0_csr_r2[2]), .DIN2(n32037), .Q(n32048) );
  and2s1 U24346 ( .DIN1(wb_data_i[26]), .DIN2(n32038), .Q(n32047) );
  or2s1 U24347 ( .DIN1(n32049), .DIN2(n32050), .Q(n9956) );
  and2s1 U24348 ( .DIN1(u0_csr_r2[1]), .DIN2(n32037), .Q(n32050) );
  and2s1 U24349 ( .DIN1(wb_data_i[25]), .DIN2(n32038), .Q(n32049) );
  or2s1 U24350 ( .DIN1(n32051), .DIN2(n32052), .Q(n9955) );
  and2s1 U24351 ( .DIN1(u0_csr_r2[0]), .DIN2(n32037), .Q(n32052) );
  and2s1 U24352 ( .DIN1(wb_data_i[24]), .DIN2(n32038), .Q(n32051) );
  or2s1 U24353 ( .DIN1(n32053), .DIN2(n32054), .Q(n9954) );
  and2s1 U24354 ( .DIN1(u0_csr_tj_val[7]), .DIN2(n32037), .Q(n32054) );
  and2s1 U24355 ( .DIN1(wb_data_i[23]), .DIN2(n32038), .Q(n32053) );
  or2s1 U24356 ( .DIN1(n32055), .DIN2(n32056), .Q(n9953) );
  and2s1 U24357 ( .DIN1(n32037), .DIN2(n32057), .Q(n32056) );
  and2s1 U24358 ( .DIN1(wb_data_i[22]), .DIN2(n32038), .Q(n32055) );
  or2s1 U24359 ( .DIN1(n32058), .DIN2(n32059), .Q(n9952) );
  and2s1 U24360 ( .DIN1(n32037), .DIN2(n32060), .Q(n32059) );
  and2s1 U24361 ( .DIN1(wb_data_i[21]), .DIN2(n32038), .Q(n32058) );
  or2s1 U24362 ( .DIN1(n32061), .DIN2(n32062), .Q(n9951) );
  and2s1 U24363 ( .DIN1(n32037), .DIN2(n32063), .Q(n32062) );
  and2s1 U24364 ( .DIN1(wb_data_i[20]), .DIN2(n32038), .Q(n32061) );
  or2s1 U24365 ( .DIN1(n32064), .DIN2(n32065), .Q(n9950) );
  and2s1 U24366 ( .DIN1(u0_csr_tj_val[3]), .DIN2(n32037), .Q(n32065) );
  and2s1 U24367 ( .DIN1(wb_data_i[19]), .DIN2(n32038), .Q(n32064) );
  or2s1 U24368 ( .DIN1(n32066), .DIN2(n32067), .Q(n9949) );
  and2s1 U24369 ( .DIN1(n32037), .DIN2(n32068), .Q(n32067) );
  and2s1 U24370 ( .DIN1(wb_data_i[18]), .DIN2(n32038), .Q(n32066) );
  or2s1 U24371 ( .DIN1(n32069), .DIN2(n32070), .Q(n9948) );
  and2s1 U24372 ( .DIN1(n32037), .DIN2(n32071), .Q(n32070) );
  and2s1 U24373 ( .DIN1(wb_data_i[17]), .DIN2(n32038), .Q(n32069) );
  or2s1 U24374 ( .DIN1(n32072), .DIN2(n32073), .Q(n9947) );
  and2s1 U24375 ( .DIN1(n32037), .DIN2(n32074), .Q(n32073) );
  and2s1 U24376 ( .DIN1(wb_data_i[16]), .DIN2(n32038), .Q(n32072) );
  or2s1 U24377 ( .DIN1(n32075), .DIN2(n32076), .Q(n9946) );
  and2s1 U24378 ( .DIN1(u0_csr_r[10]), .DIN2(n32037), .Q(n32076) );
  and2s1 U24379 ( .DIN1(wb_data_i[10]), .DIN2(n32038), .Q(n32075) );
  or2s1 U24380 ( .DIN1(n32077), .DIN2(n32078), .Q(n9945) );
  and2s1 U24381 ( .DIN1(u0_csr_r[9]), .DIN2(n32037), .Q(n32078) );
  and2s1 U24382 ( .DIN1(wb_data_i[9]), .DIN2(n32038), .Q(n32077) );
  or2s1 U24383 ( .DIN1(n32079), .DIN2(n32080), .Q(n9944) );
  and2s1 U24384 ( .DIN1(u0_csr_r[8]), .DIN2(n32037), .Q(n32080) );
  and2s1 U24385 ( .DIN1(wb_data_i[8]), .DIN2(n32038), .Q(n32079) );
  or2s1 U24386 ( .DIN1(n32081), .DIN2(n32082), .Q(n9943) );
  and2s1 U24387 ( .DIN1(n32037), .DIN2(n32083), .Q(n32082) );
  and2s1 U24388 ( .DIN1(wb_data_i[7]), .DIN2(n32038), .Q(n32081) );
  or2s1 U24389 ( .DIN1(n32084), .DIN2(n32085), .Q(n9942) );
  and2s1 U24390 ( .DIN1(n32037), .DIN2(n32086), .Q(n32085) );
  and2s1 U24391 ( .DIN1(wb_data_i[6]), .DIN2(n32038), .Q(n32084) );
  or2s1 U24392 ( .DIN1(n32087), .DIN2(n32088), .Q(n9941) );
  and2s1 U24393 ( .DIN1(n32037), .DIN2(n32089), .Q(n32088) );
  and2s1 U24394 ( .DIN1(wb_data_i[5]), .DIN2(n32038), .Q(n32087) );
  or2s1 U24395 ( .DIN1(n32090), .DIN2(n32091), .Q(n9940) );
  and2s1 U24396 ( .DIN1(n32037), .DIN2(n32092), .Q(n32091) );
  and2s1 U24397 ( .DIN1(wb_data_i[4]), .DIN2(n32038), .Q(n32090) );
  or2s1 U24398 ( .DIN1(n32093), .DIN2(n32094), .Q(n9939) );
  and2s1 U24399 ( .DIN1(n32037), .DIN2(n32095), .Q(n32094) );
  and2s1 U24400 ( .DIN1(wb_data_i[3]), .DIN2(n32038), .Q(n32093) );
  or2s1 U24401 ( .DIN1(n32096), .DIN2(n32097), .Q(n9938) );
  and2s1 U24402 ( .DIN1(n32037), .DIN2(n32098), .Q(n32097) );
  and2s1 U24403 ( .DIN1(wb_data_i[2]), .DIN2(n32038), .Q(n32096) );
  or2s1 U24404 ( .DIN1(n32099), .DIN2(n32100), .Q(n9937) );
  and2s1 U24405 ( .DIN1(n32037), .DIN2(n32101), .Q(n32100) );
  and2s1 U24406 ( .DIN1(wb_data_i[1]), .DIN2(n32038), .Q(n32099) );
  or2s1 U24407 ( .DIN1(n32102), .DIN2(n32103), .Q(n9936) );
  hi1s1 U24408 ( .DIN1(n15488), .Q(n32103) );
  and2s1 U24409 ( .DIN1(n32104), .DIN2(n32105), .Q(n32102) );
  and2s1 U24410 ( .DIN1(n32106), .DIN2(n32107), .Q(n32105) );
  hi1s1 U24411 ( .DIN1(n32108), .Q(n32107) );
  or2s1 U24412 ( .DIN1(u0_csr_tj_val[3]), .DIN2(u0_csr_tj_val[7]), .Q(n32108) );
  and2s1 U24413 ( .DIN1(n32060), .DIN2(n32057), .Q(n32106) );
  hi1s1 U24414 ( .DIN1(n36579), .Q(n32057) );
  hi1s1 U24415 ( .DIN1(n36580), .Q(n32060) );
  and2s1 U24416 ( .DIN1(n32109), .DIN2(n32110), .Q(n32104) );
  and2s1 U24417 ( .DIN1(n32068), .DIN2(n32063), .Q(n32110) );
  hi1s1 U24418 ( .DIN1(n36581), .Q(n32063) );
  hi1s1 U24419 ( .DIN1(n36582), .Q(n32068) );
  and2s1 U24420 ( .DIN1(n32074), .DIN2(n32071), .Q(n32109) );
  hi1s1 U24421 ( .DIN1(n36583), .Q(n32071) );
  hi1s1 U24422 ( .DIN1(n36584), .Q(n32074) );
  or2s1 U24423 ( .DIN1(n32111), .DIN2(n32112), .Q(n9935) );
  and2s1 U24424 ( .DIN1(n32113), .DIN2(n32114), .Q(n32112) );
  and2s1 U24425 ( .DIN1(n32115), .DIN2(wb_data_i[10]), .Q(n32111) );
  or2s1 U24426 ( .DIN1(n32116), .DIN2(n32117), .Q(n9934) );
  and2s1 U24427 ( .DIN1(n32113), .DIN2(n32118), .Q(n32117) );
  and2s1 U24428 ( .DIN1(n32115), .DIN2(wb_data_i[9]), .Q(n32116) );
  or2s1 U24429 ( .DIN1(n32119), .DIN2(n32120), .Q(n9933) );
  and2s1 U24430 ( .DIN1(n32113), .DIN2(n32121), .Q(n32120) );
  and2s1 U24431 ( .DIN1(n32115), .DIN2(wb_data_i[8]), .Q(n32119) );
  or2s1 U24432 ( .DIN1(n32122), .DIN2(n32123), .Q(n9932) );
  and2s1 U24433 ( .DIN1(u0_csc_mask_r[7]), .DIN2(n32113), .Q(n32123) );
  and2s1 U24434 ( .DIN1(n32115), .DIN2(wb_data_i[7]), .Q(n32122) );
  or2s1 U24435 ( .DIN1(n32124), .DIN2(n32125), .Q(n9931) );
  and2s1 U24436 ( .DIN1(u0_csc_mask_r[6]), .DIN2(n32113), .Q(n32125) );
  and2s1 U24437 ( .DIN1(n32115), .DIN2(wb_data_i[6]), .Q(n32124) );
  or2s1 U24438 ( .DIN1(n32126), .DIN2(n32127), .Q(n9930) );
  and2s1 U24439 ( .DIN1(u0_csc_mask_r[5]), .DIN2(n32113), .Q(n32127) );
  and2s1 U24440 ( .DIN1(n32115), .DIN2(wb_data_i[5]), .Q(n32126) );
  or2s1 U24441 ( .DIN1(n32128), .DIN2(n32129), .Q(n9929) );
  and2s1 U24442 ( .DIN1(u0_csc_mask_r[4]), .DIN2(n32113), .Q(n32129) );
  and2s1 U24443 ( .DIN1(n32115), .DIN2(wb_data_i[4]), .Q(n32128) );
  or2s1 U24444 ( .DIN1(n32130), .DIN2(n32131), .Q(n9928) );
  and2s1 U24445 ( .DIN1(u0_csc_mask_r[3]), .DIN2(n32113), .Q(n32131) );
  and2s1 U24446 ( .DIN1(n32115), .DIN2(wb_data_i[3]), .Q(n32130) );
  or2s1 U24447 ( .DIN1(n32132), .DIN2(n32133), .Q(n9927) );
  and2s1 U24448 ( .DIN1(u0_csc_mask_r[2]), .DIN2(n32113), .Q(n32133) );
  and2s1 U24449 ( .DIN1(n32115), .DIN2(wb_data_i[2]), .Q(n32132) );
  or2s1 U24450 ( .DIN1(n32134), .DIN2(n32135), .Q(n9926) );
  and2s1 U24451 ( .DIN1(u0_csc_mask_r[1]), .DIN2(n32113), .Q(n32135) );
  and2s1 U24452 ( .DIN1(n32115), .DIN2(wb_data_i[1]), .Q(n32134) );
  or2s1 U24453 ( .DIN1(n32136), .DIN2(n32137), .Q(n9925) );
  and2s1 U24454 ( .DIN1(u0_csc_mask_r[0]), .DIN2(n32113), .Q(n32137) );
  hi1s1 U24455 ( .DIN1(n32115), .Q(n32113) );
  and2s1 U24456 ( .DIN1(wb_data_i[0]), .DIN2(n32115), .Q(n32136) );
  and2s1 U24457 ( .DIN1(n32138), .DIN2(u0_wb_addr_r[3]), .Q(n32115) );
  hi1s1 U24458 ( .DIN1(n32139), .Q(n32138) );
  or2s1 U24459 ( .DIN1(n32140), .DIN2(n32141), .Q(n9921) );
  and2s1 U24460 ( .DIN1(n32142), .DIN2(wb_data_i[31]), .Q(n32141) );
  and2s1 U24461 ( .DIN1(n32143), .DIN2(n32144), .Q(n32140) );
  or2s1 U24462 ( .DIN1(n32145), .DIN2(n32146), .Q(n9920) );
  and2s1 U24463 ( .DIN1(n32142), .DIN2(wb_data_i[30]), .Q(n32146) );
  and2s1 U24464 ( .DIN1(n32143), .DIN2(n32147), .Q(n32145) );
  or2s1 U24465 ( .DIN1(n32148), .DIN2(n32149), .Q(n9919) );
  and2s1 U24466 ( .DIN1(n32142), .DIN2(wb_data_i[29]), .Q(n32149) );
  and2s1 U24467 ( .DIN1(n32143), .DIN2(n32150), .Q(n32148) );
  or2s1 U24468 ( .DIN1(n32151), .DIN2(n32152), .Q(n9918) );
  and2s1 U24469 ( .DIN1(n32142), .DIN2(wb_data_i[28]), .Q(n32152) );
  and2s1 U24470 ( .DIN1(n32143), .DIN2(n32153), .Q(n32151) );
  or2s1 U24471 ( .DIN1(n32154), .DIN2(n32155), .Q(n9917) );
  and2s1 U24472 ( .DIN1(n32142), .DIN2(wb_data_i[27]), .Q(n32155) );
  and2s1 U24473 ( .DIN1(n32143), .DIN2(n32156), .Q(n32154) );
  or2s1 U24474 ( .DIN1(n32157), .DIN2(n32158), .Q(n9916) );
  and2s1 U24475 ( .DIN1(n32142), .DIN2(wb_data_i[26]), .Q(n32158) );
  and2s1 U24476 ( .DIN1(n32143), .DIN2(n32159), .Q(n32157) );
  or2s1 U24477 ( .DIN1(n32160), .DIN2(n32161), .Q(n9915) );
  and2s1 U24478 ( .DIN1(n32142), .DIN2(wb_data_i[25]), .Q(n32161) );
  and2s1 U24479 ( .DIN1(n32143), .DIN2(n32162), .Q(n32160) );
  or2s1 U24480 ( .DIN1(n32163), .DIN2(n32164), .Q(n9914) );
  and2s1 U24481 ( .DIN1(n32142), .DIN2(wb_data_i[24]), .Q(n32164) );
  and2s1 U24482 ( .DIN1(n32143), .DIN2(n32165), .Q(n32163) );
  or2s1 U24483 ( .DIN1(n32166), .DIN2(n32167), .Q(n9913) );
  and2s1 U24484 ( .DIN1(n32142), .DIN2(wb_data_i[23]), .Q(n32167) );
  and2s1 U24485 ( .DIN1(u0_csc0[23]), .DIN2(n32143), .Q(n32166) );
  or2s1 U24486 ( .DIN1(n32168), .DIN2(n32169), .Q(n9912) );
  and2s1 U24487 ( .DIN1(n32142), .DIN2(wb_data_i[22]), .Q(n32169) );
  and2s1 U24488 ( .DIN1(u0_csc0[22]), .DIN2(n32143), .Q(n32168) );
  or2s1 U24489 ( .DIN1(n32170), .DIN2(n32171), .Q(n9911) );
  and2s1 U24490 ( .DIN1(n32142), .DIN2(wb_data_i[21]), .Q(n32171) );
  and2s1 U24491 ( .DIN1(u0_csc0[21]), .DIN2(n32143), .Q(n32170) );
  or2s1 U24492 ( .DIN1(n32172), .DIN2(n32173), .Q(n9910) );
  and2s1 U24493 ( .DIN1(n32142), .DIN2(wb_data_i[20]), .Q(n32173) );
  and2s1 U24494 ( .DIN1(u0_csc0[20]), .DIN2(n32143), .Q(n32172) );
  or2s1 U24495 ( .DIN1(n32174), .DIN2(n32175), .Q(n9909) );
  and2s1 U24496 ( .DIN1(n32142), .DIN2(wb_data_i[19]), .Q(n32175) );
  and2s1 U24497 ( .DIN1(u0_csc0[19]), .DIN2(n32143), .Q(n32174) );
  or2s1 U24498 ( .DIN1(n32176), .DIN2(n32177), .Q(n9908) );
  and2s1 U24499 ( .DIN1(n32142), .DIN2(wb_data_i[18]), .Q(n32177) );
  and2s1 U24500 ( .DIN1(u0_csc0[18]), .DIN2(n32143), .Q(n32176) );
  or2s1 U24501 ( .DIN1(n32178), .DIN2(n32179), .Q(n9907) );
  and2s1 U24502 ( .DIN1(n32142), .DIN2(wb_data_i[17]), .Q(n32179) );
  and2s1 U24503 ( .DIN1(u0_csc0[17]), .DIN2(n32143), .Q(n32178) );
  or2s1 U24504 ( .DIN1(n32180), .DIN2(n32181), .Q(n9906) );
  and2s1 U24505 ( .DIN1(n32142), .DIN2(wb_data_i[16]), .Q(n32181) );
  and2s1 U24506 ( .DIN1(u0_csc0[16]), .DIN2(n32143), .Q(n32180) );
  or2s1 U24507 ( .DIN1(n32182), .DIN2(n32183), .Q(n9905) );
  and2s1 U24508 ( .DIN1(wb_data_i[15]), .DIN2(n32142), .Q(n32183) );
  and2s1 U24509 ( .DIN1(n32143), .DIN2(n32184), .Q(n32182) );
  or2s1 U24510 ( .DIN1(n32185), .DIN2(n32186), .Q(n9904) );
  and2s1 U24511 ( .DIN1(wb_data_i[14]), .DIN2(n32142), .Q(n32186) );
  and2s1 U24512 ( .DIN1(n32143), .DIN2(n32187), .Q(n32185) );
  or2s1 U24513 ( .DIN1(n32188), .DIN2(n32189), .Q(n9903) );
  and2s1 U24514 ( .DIN1(wb_data_i[13]), .DIN2(n32142), .Q(n32189) );
  and2s1 U24515 ( .DIN1(n32143), .DIN2(n32190), .Q(n32188) );
  or2s1 U24516 ( .DIN1(n32191), .DIN2(n32192), .Q(n9902) );
  and2s1 U24517 ( .DIN1(wb_data_i[12]), .DIN2(n32142), .Q(n32192) );
  and2s1 U24518 ( .DIN1(n32143), .DIN2(n32193), .Q(n32191) );
  or2s1 U24519 ( .DIN1(n32194), .DIN2(n32195), .Q(n9901) );
  and2s1 U24520 ( .DIN1(wb_data_i[11]), .DIN2(n32142), .Q(n32195) );
  and2s1 U24521 ( .DIN1(n32143), .DIN2(n32196), .Q(n32194) );
  or2s1 U24522 ( .DIN1(n32197), .DIN2(n32198), .Q(n9900) );
  and2s1 U24523 ( .DIN1(n32142), .DIN2(wb_data_i[10]), .Q(n32198) );
  and2s1 U24524 ( .DIN1(n32143), .DIN2(n32199), .Q(n32197) );
  or2s1 U24525 ( .DIN1(n32200), .DIN2(n32201), .Q(n9899) );
  and2s1 U24526 ( .DIN1(n32142), .DIN2(wb_data_i[9]), .Q(n32201) );
  and2s1 U24527 ( .DIN1(n32143), .DIN2(n32202), .Q(n32200) );
  or2s1 U24528 ( .DIN1(n32203), .DIN2(n32204), .Q(n9898) );
  and2s1 U24529 ( .DIN1(n32142), .DIN2(wb_data_i[8]), .Q(n32204) );
  and2s1 U24530 ( .DIN1(u0_csc0[8]), .DIN2(n32143), .Q(n32203) );
  or2s1 U24531 ( .DIN1(n32205), .DIN2(n32206), .Q(n9897) );
  and2s1 U24532 ( .DIN1(n32142), .DIN2(wb_data_i[7]), .Q(n32206) );
  and2s1 U24533 ( .DIN1(n32143), .DIN2(n32207), .Q(n32205) );
  or2s1 U24534 ( .DIN1(n32208), .DIN2(n32209), .Q(n9896) );
  and2s1 U24535 ( .DIN1(n32142), .DIN2(wb_data_i[6]), .Q(n32209) );
  and2s1 U24536 ( .DIN1(n32143), .DIN2(n32210), .Q(n32208) );
  or2s1 U24537 ( .DIN1(n32211), .DIN2(n32212), .Q(n9895) );
  and2s1 U24538 ( .DIN1(n32142), .DIN2(wb_data_i[3]), .Q(n32212) );
  and2s1 U24539 ( .DIN1(u0_csc0[3]), .DIN2(n32143), .Q(n32211) );
  or2s1 U24540 ( .DIN1(n32213), .DIN2(n32214), .Q(n9894) );
  or2s1 U24541 ( .DIN1(n32215), .DIN2(n32216), .Q(n32214) );
  and2s1 U24542 ( .DIN1(n32217), .DIN2(n32218), .Q(n32216) );
  and2s1 U24543 ( .DIN1(n19406), .DIN2(wb_data_i[31]), .Q(n32215) );
  or2s1 U24544 ( .DIN1(n32213), .DIN2(n32219), .Q(n9893) );
  or2s1 U24545 ( .DIN1(n32220), .DIN2(n32221), .Q(n32219) );
  and2s1 U24546 ( .DIN1(n32217), .DIN2(n32222), .Q(n32221) );
  and2s1 U24547 ( .DIN1(n19406), .DIN2(wb_data_i[30]), .Q(n32220) );
  or2s1 U24548 ( .DIN1(n32213), .DIN2(n32223), .Q(n9892) );
  or2s1 U24549 ( .DIN1(n32224), .DIN2(n32225), .Q(n32223) );
  and2s1 U24550 ( .DIN1(n32217), .DIN2(n32226), .Q(n32225) );
  and2s1 U24551 ( .DIN1(n19406), .DIN2(wb_data_i[29]), .Q(n32224) );
  or2s1 U24552 ( .DIN1(n32213), .DIN2(n32227), .Q(n9891) );
  or2s1 U24553 ( .DIN1(n32228), .DIN2(n32229), .Q(n32227) );
  and2s1 U24554 ( .DIN1(n32217), .DIN2(n32230), .Q(n32229) );
  and2s1 U24555 ( .DIN1(n19406), .DIN2(wb_data_i[28]), .Q(n32228) );
  or2s1 U24556 ( .DIN1(n32213), .DIN2(n32231), .Q(n9890) );
  or2s1 U24557 ( .DIN1(n32232), .DIN2(n32233), .Q(n32231) );
  and2s1 U24558 ( .DIN1(n32217), .DIN2(n32234), .Q(n32233) );
  and2s1 U24559 ( .DIN1(n19406), .DIN2(wb_data_i[27]), .Q(n32232) );
  or2s1 U24560 ( .DIN1(n32213), .DIN2(n32235), .Q(n9889) );
  or2s1 U24561 ( .DIN1(n32236), .DIN2(n32237), .Q(n32235) );
  and2s1 U24562 ( .DIN1(n32217), .DIN2(n32238), .Q(n32237) );
  and2s1 U24563 ( .DIN1(n19406), .DIN2(wb_data_i[26]), .Q(n32236) );
  or2s1 U24564 ( .DIN1(n32213), .DIN2(n32239), .Q(n9888) );
  or2s1 U24565 ( .DIN1(n32240), .DIN2(n32241), .Q(n32239) );
  and2s1 U24566 ( .DIN1(n32217), .DIN2(n32242), .Q(n32241) );
  and2s1 U24567 ( .DIN1(n19406), .DIN2(wb_data_i[25]), .Q(n32240) );
  or2s1 U24568 ( .DIN1(n32213), .DIN2(n32243), .Q(n9887) );
  or2s1 U24569 ( .DIN1(n32244), .DIN2(n32245), .Q(n32243) );
  and2s1 U24570 ( .DIN1(n32217), .DIN2(n32246), .Q(n32245) );
  and2s1 U24571 ( .DIN1(n19406), .DIN2(wb_data_i[24]), .Q(n32244) );
  or2s1 U24572 ( .DIN1(n32213), .DIN2(n32247), .Q(n9886) );
  or2s1 U24573 ( .DIN1(n32248), .DIN2(n32249), .Q(n32247) );
  and2s1 U24574 ( .DIN1(n32217), .DIN2(n32250), .Q(n32249) );
  and2s1 U24575 ( .DIN1(n19406), .DIN2(wb_data_i[23]), .Q(n32248) );
  or2s1 U24576 ( .DIN1(n32213), .DIN2(n32251), .Q(n9885) );
  or2s1 U24577 ( .DIN1(n32252), .DIN2(n32253), .Q(n32251) );
  and2s1 U24578 ( .DIN1(n32217), .DIN2(n32254), .Q(n32253) );
  and2s1 U24579 ( .DIN1(n19406), .DIN2(wb_data_i[22]), .Q(n32252) );
  or2s1 U24580 ( .DIN1(n32213), .DIN2(n32255), .Q(n9884) );
  or2s1 U24581 ( .DIN1(n32256), .DIN2(n32257), .Q(n32255) );
  and2s1 U24582 ( .DIN1(n32217), .DIN2(n32258), .Q(n32257) );
  and2s1 U24583 ( .DIN1(n19406), .DIN2(wb_data_i[21]), .Q(n32256) );
  or2s1 U24584 ( .DIN1(n32213), .DIN2(n32259), .Q(n9883) );
  or2s1 U24585 ( .DIN1(n32260), .DIN2(n32261), .Q(n32259) );
  and2s1 U24586 ( .DIN1(n32217), .DIN2(n32262), .Q(n32261) );
  and2s1 U24587 ( .DIN1(n19406), .DIN2(wb_data_i[20]), .Q(n32260) );
  or2s1 U24588 ( .DIN1(n32213), .DIN2(n32263), .Q(n9882) );
  or2s1 U24589 ( .DIN1(n32264), .DIN2(n32265), .Q(n32263) );
  and2s1 U24590 ( .DIN1(n32217), .DIN2(n32266), .Q(n32265) );
  and2s1 U24591 ( .DIN1(n19406), .DIN2(wb_data_i[19]), .Q(n32264) );
  or2s1 U24592 ( .DIN1(n32213), .DIN2(n32267), .Q(n9881) );
  or2s1 U24593 ( .DIN1(n32268), .DIN2(n32269), .Q(n32267) );
  and2s1 U24594 ( .DIN1(n32217), .DIN2(n32270), .Q(n32269) );
  and2s1 U24595 ( .DIN1(n19406), .DIN2(wb_data_i[18]), .Q(n32268) );
  or2s1 U24596 ( .DIN1(n32213), .DIN2(n32271), .Q(n9880) );
  or2s1 U24597 ( .DIN1(n32272), .DIN2(n32273), .Q(n32271) );
  and2s1 U24598 ( .DIN1(n32217), .DIN2(n32274), .Q(n32273) );
  and2s1 U24599 ( .DIN1(n19406), .DIN2(wb_data_i[17]), .Q(n32272) );
  or2s1 U24600 ( .DIN1(n32213), .DIN2(n32275), .Q(n9879) );
  or2s1 U24601 ( .DIN1(n32276), .DIN2(n32277), .Q(n32275) );
  and2s1 U24602 ( .DIN1(n32217), .DIN2(n32278), .Q(n32277) );
  and2s1 U24603 ( .DIN1(n19406), .DIN2(wb_data_i[16]), .Q(n32276) );
  or2s1 U24604 ( .DIN1(n32213), .DIN2(n32279), .Q(n9878) );
  or2s1 U24605 ( .DIN1(n32280), .DIN2(n32281), .Q(n32279) );
  and2s1 U24606 ( .DIN1(n32217), .DIN2(n32282), .Q(n32281) );
  and2s1 U24607 ( .DIN1(n19406), .DIN2(wb_data_i[15]), .Q(n32280) );
  or2s1 U24608 ( .DIN1(n32213), .DIN2(n32283), .Q(n9877) );
  or2s1 U24609 ( .DIN1(n32284), .DIN2(n32285), .Q(n32283) );
  and2s1 U24610 ( .DIN1(n32217), .DIN2(n32286), .Q(n32285) );
  and2s1 U24611 ( .DIN1(n19406), .DIN2(wb_data_i[14]), .Q(n32284) );
  or2s1 U24612 ( .DIN1(n32213), .DIN2(n32287), .Q(n9876) );
  or2s1 U24613 ( .DIN1(n32288), .DIN2(n32289), .Q(n32287) );
  and2s1 U24614 ( .DIN1(n32217), .DIN2(n32290), .Q(n32289) );
  and2s1 U24615 ( .DIN1(n19406), .DIN2(wb_data_i[13]), .Q(n32288) );
  or2s1 U24616 ( .DIN1(n32213), .DIN2(n32291), .Q(n9875) );
  or2s1 U24617 ( .DIN1(n32292), .DIN2(n32293), .Q(n32291) );
  and2s1 U24618 ( .DIN1(n32217), .DIN2(n32294), .Q(n32293) );
  and2s1 U24619 ( .DIN1(n19406), .DIN2(wb_data_i[12]), .Q(n32292) );
  or2s1 U24620 ( .DIN1(n32213), .DIN2(n32295), .Q(n9874) );
  or2s1 U24621 ( .DIN1(n32296), .DIN2(n32297), .Q(n32295) );
  and2s1 U24622 ( .DIN1(n32217), .DIN2(n32298), .Q(n32297) );
  and2s1 U24623 ( .DIN1(n19406), .DIN2(wb_data_i[11]), .Q(n32296) );
  or2s1 U24624 ( .DIN1(n32213), .DIN2(n32299), .Q(n9873) );
  or2s1 U24625 ( .DIN1(n32300), .DIN2(n32301), .Q(n32299) );
  and2s1 U24626 ( .DIN1(n32217), .DIN2(n32302), .Q(n32301) );
  and2s1 U24627 ( .DIN1(n19406), .DIN2(wb_data_i[10]), .Q(n32300) );
  or2s1 U24628 ( .DIN1(n32213), .DIN2(n32303), .Q(n9872) );
  or2s1 U24629 ( .DIN1(n32304), .DIN2(n32305), .Q(n32303) );
  and2s1 U24630 ( .DIN1(n32217), .DIN2(n32306), .Q(n32305) );
  and2s1 U24631 ( .DIN1(n19406), .DIN2(wb_data_i[9]), .Q(n32304) );
  or2s1 U24632 ( .DIN1(n32213), .DIN2(n32307), .Q(n9871) );
  or2s1 U24633 ( .DIN1(n32308), .DIN2(n32309), .Q(n32307) );
  and2s1 U24634 ( .DIN1(n32217), .DIN2(n32310), .Q(n32309) );
  and2s1 U24635 ( .DIN1(n19406), .DIN2(wb_data_i[8]), .Q(n32308) );
  or2s1 U24636 ( .DIN1(n32213), .DIN2(n32311), .Q(n9870) );
  or2s1 U24637 ( .DIN1(n32312), .DIN2(n32313), .Q(n32311) );
  and2s1 U24638 ( .DIN1(n32217), .DIN2(n32314), .Q(n32313) );
  and2s1 U24639 ( .DIN1(n19406), .DIN2(wb_data_i[7]), .Q(n32312) );
  or2s1 U24640 ( .DIN1(n32213), .DIN2(n32315), .Q(n9869) );
  or2s1 U24641 ( .DIN1(n32316), .DIN2(n32317), .Q(n32315) );
  and2s1 U24642 ( .DIN1(n32217), .DIN2(n32318), .Q(n32317) );
  and2s1 U24643 ( .DIN1(n19406), .DIN2(wb_data_i[6]), .Q(n32316) );
  or2s1 U24644 ( .DIN1(n32213), .DIN2(n32319), .Q(n9868) );
  or2s1 U24645 ( .DIN1(n32320), .DIN2(n32321), .Q(n32319) );
  and2s1 U24646 ( .DIN1(n32217), .DIN2(n32322), .Q(n32321) );
  and2s1 U24647 ( .DIN1(n19406), .DIN2(wb_data_i[5]), .Q(n32320) );
  or2s1 U24648 ( .DIN1(n32213), .DIN2(n32323), .Q(n9867) );
  or2s1 U24649 ( .DIN1(n32324), .DIN2(n32325), .Q(n32323) );
  and2s1 U24650 ( .DIN1(n32217), .DIN2(n32326), .Q(n32325) );
  and2s1 U24651 ( .DIN1(n19406), .DIN2(wb_data_i[4]), .Q(n32324) );
  or2s1 U24652 ( .DIN1(n32213), .DIN2(n32327), .Q(n9866) );
  or2s1 U24653 ( .DIN1(n32328), .DIN2(n32329), .Q(n32327) );
  and2s1 U24654 ( .DIN1(n32217), .DIN2(n32330), .Q(n32329) );
  and2s1 U24655 ( .DIN1(n19406), .DIN2(wb_data_i[3]), .Q(n32328) );
  or2s1 U24656 ( .DIN1(n32213), .DIN2(n32331), .Q(n9865) );
  or2s1 U24657 ( .DIN1(n32332), .DIN2(n32333), .Q(n32331) );
  and2s1 U24658 ( .DIN1(n32217), .DIN2(n32334), .Q(n32333) );
  and2s1 U24659 ( .DIN1(n19406), .DIN2(wb_data_i[2]), .Q(n32332) );
  or2s1 U24660 ( .DIN1(n32213), .DIN2(n32335), .Q(n9864) );
  or2s1 U24661 ( .DIN1(n32336), .DIN2(n32337), .Q(n32335) );
  and2s1 U24662 ( .DIN1(n32217), .DIN2(n32338), .Q(n32337) );
  and2s1 U24663 ( .DIN1(n19406), .DIN2(wb_data_i[1]), .Q(n32336) );
  or2s1 U24664 ( .DIN1(n32213), .DIN2(n32339), .Q(n9863) );
  or2s1 U24665 ( .DIN1(n32340), .DIN2(n32341), .Q(n32339) );
  and2s1 U24666 ( .DIN1(n32217), .DIN2(n32342), .Q(n32341) );
  and2s1 U24667 ( .DIN1(n19406), .DIN2(wb_data_i[0]), .Q(n32340) );
  or2s1 U24668 ( .DIN1(n32343), .DIN2(n32344), .Q(n9859) );
  and2s1 U24669 ( .DIN1(n32345), .DIN2(wb_data_i[31]), .Q(n32344) );
  and2s1 U24670 ( .DIN1(n32346), .DIN2(n32347), .Q(n32343) );
  or2s1 U24671 ( .DIN1(n32348), .DIN2(n32349), .Q(n9858) );
  and2s1 U24672 ( .DIN1(n32345), .DIN2(wb_data_i[30]), .Q(n32349) );
  and2s1 U24673 ( .DIN1(n32346), .DIN2(n32350), .Q(n32348) );
  or2s1 U24674 ( .DIN1(n32351), .DIN2(n32352), .Q(n9857) );
  and2s1 U24675 ( .DIN1(n32345), .DIN2(wb_data_i[29]), .Q(n32352) );
  and2s1 U24676 ( .DIN1(n32346), .DIN2(n32353), .Q(n32351) );
  or2s1 U24677 ( .DIN1(n32354), .DIN2(n32355), .Q(n9856) );
  and2s1 U24678 ( .DIN1(n32345), .DIN2(wb_data_i[28]), .Q(n32355) );
  and2s1 U24679 ( .DIN1(n32346), .DIN2(n32356), .Q(n32354) );
  or2s1 U24680 ( .DIN1(n32357), .DIN2(n32358), .Q(n9855) );
  and2s1 U24681 ( .DIN1(n32345), .DIN2(wb_data_i[27]), .Q(n32358) );
  and2s1 U24682 ( .DIN1(n32346), .DIN2(n32359), .Q(n32357) );
  or2s1 U24683 ( .DIN1(n32360), .DIN2(n32361), .Q(n9854) );
  and2s1 U24684 ( .DIN1(n32345), .DIN2(wb_data_i[26]), .Q(n32361) );
  and2s1 U24685 ( .DIN1(n32346), .DIN2(n32362), .Q(n32360) );
  or2s1 U24686 ( .DIN1(n32363), .DIN2(n32364), .Q(n9853) );
  and2s1 U24687 ( .DIN1(n32345), .DIN2(wb_data_i[25]), .Q(n32364) );
  and2s1 U24688 ( .DIN1(n32346), .DIN2(n32365), .Q(n32363) );
  or2s1 U24689 ( .DIN1(n32366), .DIN2(n32367), .Q(n9852) );
  and2s1 U24690 ( .DIN1(n32345), .DIN2(wb_data_i[24]), .Q(n32367) );
  and2s1 U24691 ( .DIN1(n32346), .DIN2(n32368), .Q(n32366) );
  or2s1 U24692 ( .DIN1(n32369), .DIN2(n32370), .Q(n9851) );
  and2s1 U24693 ( .DIN1(n32345), .DIN2(wb_data_i[23]), .Q(n32370) );
  and2s1 U24694 ( .DIN1(u0_csc1[23]), .DIN2(n32346), .Q(n32369) );
  or2s1 U24695 ( .DIN1(n32371), .DIN2(n32372), .Q(n9850) );
  and2s1 U24696 ( .DIN1(n32345), .DIN2(wb_data_i[22]), .Q(n32372) );
  and2s1 U24697 ( .DIN1(u0_csc1[22]), .DIN2(n32346), .Q(n32371) );
  or2s1 U24698 ( .DIN1(n32373), .DIN2(n32374), .Q(n9849) );
  and2s1 U24699 ( .DIN1(n32345), .DIN2(wb_data_i[21]), .Q(n32374) );
  and2s1 U24700 ( .DIN1(u0_csc1[21]), .DIN2(n32346), .Q(n32373) );
  or2s1 U24701 ( .DIN1(n32375), .DIN2(n32376), .Q(n9848) );
  and2s1 U24702 ( .DIN1(n32345), .DIN2(wb_data_i[20]), .Q(n32376) );
  and2s1 U24703 ( .DIN1(u0_csc1[20]), .DIN2(n32346), .Q(n32375) );
  or2s1 U24704 ( .DIN1(n32377), .DIN2(n32378), .Q(n9847) );
  and2s1 U24705 ( .DIN1(n32345), .DIN2(wb_data_i[19]), .Q(n32378) );
  and2s1 U24706 ( .DIN1(u0_csc1[19]), .DIN2(n32346), .Q(n32377) );
  or2s1 U24707 ( .DIN1(n32379), .DIN2(n32380), .Q(n9846) );
  and2s1 U24708 ( .DIN1(n32345), .DIN2(wb_data_i[18]), .Q(n32380) );
  and2s1 U24709 ( .DIN1(u0_csc1[18]), .DIN2(n32346), .Q(n32379) );
  or2s1 U24710 ( .DIN1(n32381), .DIN2(n32382), .Q(n9845) );
  and2s1 U24711 ( .DIN1(n32345), .DIN2(wb_data_i[17]), .Q(n32382) );
  and2s1 U24712 ( .DIN1(u0_csc1[17]), .DIN2(n32346), .Q(n32381) );
  or2s1 U24713 ( .DIN1(n32383), .DIN2(n32384), .Q(n9844) );
  and2s1 U24714 ( .DIN1(n32345), .DIN2(wb_data_i[16]), .Q(n32384) );
  and2s1 U24715 ( .DIN1(u0_csc1[16]), .DIN2(n32346), .Q(n32383) );
  or2s1 U24716 ( .DIN1(n32385), .DIN2(n32386), .Q(n9843) );
  and2s1 U24717 ( .DIN1(n32345), .DIN2(wb_data_i[15]), .Q(n32386) );
  and2s1 U24718 ( .DIN1(n32346), .DIN2(n32387), .Q(n32385) );
  or2s1 U24719 ( .DIN1(n32388), .DIN2(n32389), .Q(n9842) );
  and2s1 U24720 ( .DIN1(n32345), .DIN2(wb_data_i[14]), .Q(n32389) );
  and2s1 U24721 ( .DIN1(n32346), .DIN2(n32390), .Q(n32388) );
  or2s1 U24722 ( .DIN1(n32391), .DIN2(n32392), .Q(n9841) );
  and2s1 U24723 ( .DIN1(n32345), .DIN2(wb_data_i[13]), .Q(n32392) );
  and2s1 U24724 ( .DIN1(n32346), .DIN2(n32393), .Q(n32391) );
  or2s1 U24725 ( .DIN1(n32394), .DIN2(n32395), .Q(n9840) );
  and2s1 U24726 ( .DIN1(n32345), .DIN2(wb_data_i[12]), .Q(n32395) );
  and2s1 U24727 ( .DIN1(n32346), .DIN2(n32396), .Q(n32394) );
  or2s1 U24728 ( .DIN1(n32397), .DIN2(n32398), .Q(n9839) );
  and2s1 U24729 ( .DIN1(n32345), .DIN2(wb_data_i[11]), .Q(n32398) );
  and2s1 U24730 ( .DIN1(n32346), .DIN2(n32399), .Q(n32397) );
  or2s1 U24731 ( .DIN1(n32400), .DIN2(n32401), .Q(n9838) );
  and2s1 U24732 ( .DIN1(n32345), .DIN2(wb_data_i[10]), .Q(n32401) );
  and2s1 U24733 ( .DIN1(n32346), .DIN2(n32402), .Q(n32400) );
  or2s1 U24734 ( .DIN1(n32403), .DIN2(n32404), .Q(n9837) );
  and2s1 U24735 ( .DIN1(n32345), .DIN2(wb_data_i[9]), .Q(n32404) );
  and2s1 U24736 ( .DIN1(n32346), .DIN2(n32405), .Q(n32403) );
  or2s1 U24737 ( .DIN1(n32406), .DIN2(n32407), .Q(n9836) );
  and2s1 U24738 ( .DIN1(n32345), .DIN2(wb_data_i[8]), .Q(n32407) );
  and2s1 U24739 ( .DIN1(u0_csc1[8]), .DIN2(n32346), .Q(n32406) );
  or2s1 U24740 ( .DIN1(n32408), .DIN2(n32409), .Q(n9835) );
  and2s1 U24741 ( .DIN1(n32345), .DIN2(wb_data_i[7]), .Q(n32409) );
  and2s1 U24742 ( .DIN1(n32346), .DIN2(n32410), .Q(n32408) );
  or2s1 U24743 ( .DIN1(n32411), .DIN2(n32412), .Q(n9834) );
  and2s1 U24744 ( .DIN1(n32345), .DIN2(wb_data_i[6]), .Q(n32412) );
  and2s1 U24745 ( .DIN1(n32346), .DIN2(n32413), .Q(n32411) );
  or2s1 U24746 ( .DIN1(n32414), .DIN2(n32415), .Q(n9833) );
  and2s1 U24747 ( .DIN1(n32345), .DIN2(wb_data_i[5]), .Q(n32415) );
  and2s1 U24748 ( .DIN1(n32346), .DIN2(n32416), .Q(n32414) );
  or2s1 U24749 ( .DIN1(n32417), .DIN2(n32418), .Q(n9832) );
  and2s1 U24750 ( .DIN1(n32345), .DIN2(wb_data_i[4]), .Q(n32418) );
  and2s1 U24751 ( .DIN1(n32346), .DIN2(n32419), .Q(n32417) );
  or2s1 U24752 ( .DIN1(n32420), .DIN2(n32421), .Q(n9831) );
  and2s1 U24753 ( .DIN1(n32345), .DIN2(wb_data_i[3]), .Q(n32421) );
  and2s1 U24754 ( .DIN1(u0_csc1[3]), .DIN2(n32346), .Q(n32420) );
  or2s1 U24755 ( .DIN1(n32422), .DIN2(n32423), .Q(n9830) );
  and2s1 U24756 ( .DIN1(n32345), .DIN2(wb_data_i[2]), .Q(n32423) );
  and2s1 U24757 ( .DIN1(u0_csc1[2]), .DIN2(n32346), .Q(n32422) );
  or2s1 U24758 ( .DIN1(n32424), .DIN2(n32425), .Q(n9829) );
  and2s1 U24759 ( .DIN1(n32345), .DIN2(wb_data_i[1]), .Q(n32425) );
  and2s1 U24760 ( .DIN1(n32346), .DIN2(n32426), .Q(n32424) );
  or2s1 U24761 ( .DIN1(n32427), .DIN2(n32428), .Q(n9828) );
  and2s1 U24762 ( .DIN1(n32345), .DIN2(wb_data_i[0]), .Q(n32428) );
  and2s1 U24763 ( .DIN1(u0_csc1[0]), .DIN2(n32346), .Q(n32427) );
  and2s1 U24764 ( .DIN1(n32429), .DIN2(n32430), .Q(n32346) );
  hi1s1 U24765 ( .DIN1(n32345), .Q(n32430) );
  and2s1 U24766 ( .DIN1(n32429), .DIN2(n9794), .Q(n32345) );
  or2s1 U24767 ( .DIN1(n32431), .DIN2(n32432), .Q(n9827) );
  and2s1 U24768 ( .DIN1(n32433), .DIN2(wb_data_i[31]), .Q(n32432) );
  and2s1 U24769 ( .DIN1(n32434), .DIN2(n32435), .Q(n32431) );
  or2s1 U24770 ( .DIN1(n32436), .DIN2(n32437), .Q(n9826) );
  and2s1 U24771 ( .DIN1(n32433), .DIN2(wb_data_i[30]), .Q(n32437) );
  and2s1 U24772 ( .DIN1(n32434), .DIN2(n32438), .Q(n32436) );
  or2s1 U24773 ( .DIN1(n32439), .DIN2(n32440), .Q(n9825) );
  and2s1 U24774 ( .DIN1(n32433), .DIN2(wb_data_i[29]), .Q(n32440) );
  and2s1 U24775 ( .DIN1(n32434), .DIN2(n32441), .Q(n32439) );
  or2s1 U24776 ( .DIN1(n32442), .DIN2(n32443), .Q(n9824) );
  and2s1 U24777 ( .DIN1(n32433), .DIN2(wb_data_i[28]), .Q(n32443) );
  and2s1 U24778 ( .DIN1(n32434), .DIN2(n32444), .Q(n32442) );
  or2s1 U24779 ( .DIN1(n32445), .DIN2(n32446), .Q(n9823) );
  and2s1 U24780 ( .DIN1(n32433), .DIN2(wb_data_i[27]), .Q(n32446) );
  and2s1 U24781 ( .DIN1(n32434), .DIN2(n32447), .Q(n32445) );
  or2s1 U24782 ( .DIN1(n32448), .DIN2(n32449), .Q(n9822) );
  and2s1 U24783 ( .DIN1(n32433), .DIN2(wb_data_i[26]), .Q(n32449) );
  and2s1 U24784 ( .DIN1(n32434), .DIN2(n32450), .Q(n32448) );
  or2s1 U24785 ( .DIN1(n32451), .DIN2(n32452), .Q(n9821) );
  and2s1 U24786 ( .DIN1(n32433), .DIN2(wb_data_i[25]), .Q(n32452) );
  and2s1 U24787 ( .DIN1(n32434), .DIN2(n32453), .Q(n32451) );
  or2s1 U24788 ( .DIN1(n32454), .DIN2(n32455), .Q(n9820) );
  and2s1 U24789 ( .DIN1(n32433), .DIN2(wb_data_i[24]), .Q(n32455) );
  and2s1 U24790 ( .DIN1(n32434), .DIN2(n32456), .Q(n32454) );
  or2s1 U24791 ( .DIN1(n32457), .DIN2(n32458), .Q(n9819) );
  and2s1 U24792 ( .DIN1(n32433), .DIN2(wb_data_i[23]), .Q(n32458) );
  and2s1 U24793 ( .DIN1(n32434), .DIN2(n32459), .Q(n32457) );
  or2s1 U24794 ( .DIN1(n32460), .DIN2(n32461), .Q(n9818) );
  and2s1 U24795 ( .DIN1(n32433), .DIN2(wb_data_i[22]), .Q(n32461) );
  and2s1 U24796 ( .DIN1(n32434), .DIN2(n32462), .Q(n32460) );
  or2s1 U24797 ( .DIN1(n32463), .DIN2(n32464), .Q(n9817) );
  and2s1 U24798 ( .DIN1(n32433), .DIN2(wb_data_i[21]), .Q(n32464) );
  and2s1 U24799 ( .DIN1(n32434), .DIN2(n32465), .Q(n32463) );
  or2s1 U24800 ( .DIN1(n32466), .DIN2(n32467), .Q(n9816) );
  and2s1 U24801 ( .DIN1(n32433), .DIN2(wb_data_i[20]), .Q(n32467) );
  and2s1 U24802 ( .DIN1(n32434), .DIN2(n32468), .Q(n32466) );
  or2s1 U24803 ( .DIN1(n32469), .DIN2(n32470), .Q(n9815) );
  and2s1 U24804 ( .DIN1(n32433), .DIN2(wb_data_i[19]), .Q(n32470) );
  and2s1 U24805 ( .DIN1(n32434), .DIN2(n32471), .Q(n32469) );
  or2s1 U24806 ( .DIN1(n32472), .DIN2(n32473), .Q(n9814) );
  and2s1 U24807 ( .DIN1(n32433), .DIN2(wb_data_i[18]), .Q(n32473) );
  and2s1 U24808 ( .DIN1(n32434), .DIN2(n32474), .Q(n32472) );
  or2s1 U24809 ( .DIN1(n32475), .DIN2(n32476), .Q(n9813) );
  and2s1 U24810 ( .DIN1(n32433), .DIN2(wb_data_i[17]), .Q(n32476) );
  and2s1 U24811 ( .DIN1(n32434), .DIN2(n32477), .Q(n32475) );
  or2s1 U24812 ( .DIN1(n32478), .DIN2(n32479), .Q(n9812) );
  and2s1 U24813 ( .DIN1(n32433), .DIN2(wb_data_i[16]), .Q(n32479) );
  and2s1 U24814 ( .DIN1(n32434), .DIN2(n32480), .Q(n32478) );
  or2s1 U24815 ( .DIN1(n32481), .DIN2(n32482), .Q(n9811) );
  and2s1 U24816 ( .DIN1(n32433), .DIN2(wb_data_i[15]), .Q(n32482) );
  and2s1 U24817 ( .DIN1(n32434), .DIN2(n32483), .Q(n32481) );
  or2s1 U24818 ( .DIN1(n32484), .DIN2(n32485), .Q(n9810) );
  and2s1 U24819 ( .DIN1(n32433), .DIN2(wb_data_i[14]), .Q(n32485) );
  and2s1 U24820 ( .DIN1(n32434), .DIN2(n32486), .Q(n32484) );
  or2s1 U24821 ( .DIN1(n32487), .DIN2(n32488), .Q(n9809) );
  and2s1 U24822 ( .DIN1(n32433), .DIN2(wb_data_i[13]), .Q(n32488) );
  and2s1 U24823 ( .DIN1(n32434), .DIN2(n32489), .Q(n32487) );
  or2s1 U24824 ( .DIN1(n32490), .DIN2(n32491), .Q(n9808) );
  and2s1 U24825 ( .DIN1(n32433), .DIN2(wb_data_i[12]), .Q(n32491) );
  and2s1 U24826 ( .DIN1(n32434), .DIN2(n32492), .Q(n32490) );
  or2s1 U24827 ( .DIN1(n32493), .DIN2(n32494), .Q(n9807) );
  and2s1 U24828 ( .DIN1(n32433), .DIN2(wb_data_i[11]), .Q(n32494) );
  and2s1 U24829 ( .DIN1(n32434), .DIN2(n32495), .Q(n32493) );
  or2s1 U24830 ( .DIN1(n32496), .DIN2(n32497), .Q(n9806) );
  and2s1 U24831 ( .DIN1(n32433), .DIN2(wb_data_i[10]), .Q(n32497) );
  and2s1 U24832 ( .DIN1(n32434), .DIN2(n32498), .Q(n32496) );
  or2s1 U24833 ( .DIN1(n32499), .DIN2(n32500), .Q(n9805) );
  and2s1 U24834 ( .DIN1(n32433), .DIN2(wb_data_i[9]), .Q(n32500) );
  and2s1 U24835 ( .DIN1(n32434), .DIN2(n32501), .Q(n32499) );
  or2s1 U24836 ( .DIN1(n32502), .DIN2(n32503), .Q(n9804) );
  and2s1 U24837 ( .DIN1(n32433), .DIN2(wb_data_i[8]), .Q(n32503) );
  and2s1 U24838 ( .DIN1(n32434), .DIN2(n32504), .Q(n32502) );
  or2s1 U24839 ( .DIN1(n32505), .DIN2(n32506), .Q(n9803) );
  and2s1 U24840 ( .DIN1(n32433), .DIN2(wb_data_i[7]), .Q(n32506) );
  and2s1 U24841 ( .DIN1(n32434), .DIN2(n32507), .Q(n32505) );
  or2s1 U24842 ( .DIN1(n32508), .DIN2(n32509), .Q(n9802) );
  and2s1 U24843 ( .DIN1(n32433), .DIN2(wb_data_i[6]), .Q(n32509) );
  and2s1 U24844 ( .DIN1(n32434), .DIN2(n32510), .Q(n32508) );
  or2s1 U24845 ( .DIN1(n32511), .DIN2(n32512), .Q(n9801) );
  and2s1 U24846 ( .DIN1(n32433), .DIN2(wb_data_i[5]), .Q(n32512) );
  and2s1 U24847 ( .DIN1(n32434), .DIN2(n32513), .Q(n32511) );
  or2s1 U24848 ( .DIN1(n32514), .DIN2(n32515), .Q(n9800) );
  and2s1 U24849 ( .DIN1(n32433), .DIN2(wb_data_i[4]), .Q(n32515) );
  and2s1 U24850 ( .DIN1(n32434), .DIN2(n32516), .Q(n32514) );
  or2s1 U24851 ( .DIN1(n32517), .DIN2(n32518), .Q(n9799) );
  and2s1 U24852 ( .DIN1(n32433), .DIN2(wb_data_i[3]), .Q(n32518) );
  and2s1 U24853 ( .DIN1(n32434), .DIN2(n32519), .Q(n32517) );
  or2s1 U24854 ( .DIN1(n32520), .DIN2(n32521), .Q(n9798) );
  and2s1 U24855 ( .DIN1(n32433), .DIN2(wb_data_i[2]), .Q(n32521) );
  and2s1 U24856 ( .DIN1(n32434), .DIN2(n32522), .Q(n32520) );
  or2s1 U24857 ( .DIN1(n32523), .DIN2(n32524), .Q(n9797) );
  and2s1 U24858 ( .DIN1(n32433), .DIN2(wb_data_i[1]), .Q(n32524) );
  and2s1 U24859 ( .DIN1(n32434), .DIN2(n32525), .Q(n32523) );
  or2s1 U24860 ( .DIN1(n32526), .DIN2(n32527), .Q(n9796) );
  and2s1 U24861 ( .DIN1(n32433), .DIN2(wb_data_i[0]), .Q(n32527) );
  and2s1 U24862 ( .DIN1(n32434), .DIN2(n32528), .Q(n32526) );
  hi1s1 U24863 ( .DIN1(n32529), .Q(n32434) );
  or2s1 U24864 ( .DIN1(n36585), .DIN2(n32433), .Q(n32529) );
  and2s1 U24865 ( .DIN1(n32429), .DIN2(n9795), .Q(n32433) );
  hi1s1 U24866 ( .DIN1(n36585), .Q(n32429) );
  and2s1 U24867 ( .DIN1(n32530), .DIN2(n32531), .Q(n9795) );
  and2s1 U24868 ( .DIN1(n36589), .DIN2(n32532), .Q(n32530) );
  and2s1 U24869 ( .DIN1(n32533), .DIN2(n36609), .Q(n32532) );
  hi1s1 U24870 ( .DIN1(n15486), .Q(n32533) );
  and2s1 U24871 ( .DIN1(n32534), .DIN2(n32531), .Q(n9794) );
  and2s1 U24872 ( .DIN1(n36586), .DIN2(n32535), .Q(n32531) );
  and2s1 U24873 ( .DIN1(n36588), .DIN2(n36587), .Q(n32535) );
  and2s1 U24874 ( .DIN1(n36589), .DIN2(n32536), .Q(n32534) );
  and2s1 U24875 ( .DIN1(n36609), .DIN2(n15486), .Q(n32536) );
  or2s1 U24876 ( .DIN1(n32537), .DIN2(n32538), .Q(n9793) );
  and2s1 U24877 ( .DIN1(wb_addr_i[25]), .DIN2(wb_stb_i), .Q(n32538) );
  and2s1 U24878 ( .DIN1(n32539), .DIN2(n32540), .Q(n32537) );
  or2s1 U24879 ( .DIN1(n32541), .DIN2(n32542), .Q(n9792) );
  and2s1 U24880 ( .DIN1(wb_addr_i[24]), .DIN2(wb_stb_i), .Q(n32542) );
  and2s1 U24881 ( .DIN1(n32543), .DIN2(n32540), .Q(n32541) );
  or2s1 U24882 ( .DIN1(n32544), .DIN2(n32545), .Q(n9791) );
  and2s1 U24883 ( .DIN1(wb_addr_i[23]), .DIN2(wb_stb_i), .Q(n32545) );
  and2s1 U24884 ( .DIN1(n32546), .DIN2(n32540), .Q(n32544) );
  or2s1 U24885 ( .DIN1(n32547), .DIN2(n32548), .Q(n9790) );
  and2s1 U24886 ( .DIN1(wb_addr_i[22]), .DIN2(wb_stb_i), .Q(n32548) );
  and2s1 U24887 ( .DIN1(n32549), .DIN2(n32540), .Q(n32547) );
  or2s1 U24888 ( .DIN1(n32550), .DIN2(n32551), .Q(n9789) );
  and2s1 U24889 ( .DIN1(wb_addr_i[21]), .DIN2(wb_stb_i), .Q(n32551) );
  and2s1 U24890 ( .DIN1(n32552), .DIN2(n32540), .Q(n32550) );
  or2s1 U24891 ( .DIN1(n32553), .DIN2(n32554), .Q(n9788) );
  and2s1 U24892 ( .DIN1(wb_addr_i[20]), .DIN2(wb_stb_i), .Q(n32554) );
  and2s1 U24893 ( .DIN1(n32555), .DIN2(n32540), .Q(n32553) );
  or2s1 U24894 ( .DIN1(n32556), .DIN2(n32557), .Q(n9787) );
  and2s1 U24895 ( .DIN1(wb_addr_i[19]), .DIN2(wb_stb_i), .Q(n32557) );
  and2s1 U24896 ( .DIN1(n32558), .DIN2(n32540), .Q(n32556) );
  or2s1 U24897 ( .DIN1(n32559), .DIN2(n32560), .Q(n9786) );
  and2s1 U24898 ( .DIN1(wb_addr_i[18]), .DIN2(wb_stb_i), .Q(n32560) );
  and2s1 U24899 ( .DIN1(n32561), .DIN2(n32540), .Q(n32559) );
  or2s1 U24900 ( .DIN1(n32562), .DIN2(n32563), .Q(n9785) );
  and2s1 U24901 ( .DIN1(wb_addr_i[17]), .DIN2(wb_stb_i), .Q(n32563) );
  and2s1 U24902 ( .DIN1(n32564), .DIN2(n32540), .Q(n32562) );
  or2s1 U24903 ( .DIN1(n32565), .DIN2(n32566), .Q(n9784) );
  and2s1 U24904 ( .DIN1(wb_addr_i[16]), .DIN2(wb_stb_i), .Q(n32566) );
  and2s1 U24905 ( .DIN1(n32567), .DIN2(n32540), .Q(n32565) );
  or2s1 U24906 ( .DIN1(n32568), .DIN2(n32569), .Q(n9783) );
  and2s1 U24907 ( .DIN1(wb_addr_i[15]), .DIN2(wb_stb_i), .Q(n32569) );
  and2s1 U24908 ( .DIN1(n32570), .DIN2(n32540), .Q(n32568) );
  or2s1 U24909 ( .DIN1(n32571), .DIN2(n32572), .Q(n9782) );
  and2s1 U24910 ( .DIN1(wb_addr_i[14]), .DIN2(wb_stb_i), .Q(n32572) );
  and2s1 U24911 ( .DIN1(n32573), .DIN2(n32540), .Q(n32571) );
  or2s1 U24912 ( .DIN1(n32574), .DIN2(n32575), .Q(n9781) );
  and2s1 U24913 ( .DIN1(wb_addr_i[13]), .DIN2(wb_stb_i), .Q(n32575) );
  and2s1 U24914 ( .DIN1(n32576), .DIN2(n32540), .Q(n32574) );
  or2s1 U24915 ( .DIN1(n32577), .DIN2(n32578), .Q(n9780) );
  and2s1 U24916 ( .DIN1(wb_addr_i[12]), .DIN2(wb_stb_i), .Q(n32578) );
  and2s1 U24917 ( .DIN1(n32579), .DIN2(n32540), .Q(n32577) );
  or2s1 U24918 ( .DIN1(n32580), .DIN2(n32581), .Q(n9779) );
  and2s1 U24919 ( .DIN1(wb_addr_i[11]), .DIN2(wb_stb_i), .Q(n32581) );
  and2s1 U24920 ( .DIN1(n32582), .DIN2(n32540), .Q(n32580) );
  or2s1 U24921 ( .DIN1(n32583), .DIN2(n32584), .Q(n9778) );
  and2s1 U24922 ( .DIN1(wb_addr_i[10]), .DIN2(wb_stb_i), .Q(n32584) );
  and2s1 U24923 ( .DIN1(n32585), .DIN2(n32540), .Q(n32583) );
  or2s1 U24924 ( .DIN1(n32586), .DIN2(n32587), .Q(n9777) );
  and2s1 U24925 ( .DIN1(wb_addr_i[9]), .DIN2(wb_stb_i), .Q(n32587) );
  and2s1 U24926 ( .DIN1(n32588), .DIN2(n32540), .Q(n32586) );
  or2s1 U24927 ( .DIN1(n32589), .DIN2(n32590), .Q(n9776) );
  and2s1 U24928 ( .DIN1(wb_addr_i[8]), .DIN2(wb_stb_i), .Q(n32590) );
  and2s1 U24929 ( .DIN1(n32591), .DIN2(n32540), .Q(n32589) );
  or2s1 U24930 ( .DIN1(n32592), .DIN2(n32593), .Q(n9775) );
  and2s1 U24931 ( .DIN1(wb_addr_i[7]), .DIN2(wb_stb_i), .Q(n32593) );
  and2s1 U24932 ( .DIN1(n32594), .DIN2(n32540), .Q(n32592) );
  or2s1 U24933 ( .DIN1(n32595), .DIN2(n32596), .Q(n9774) );
  and2s1 U24934 ( .DIN1(wb_addr_i[6]), .DIN2(wb_stb_i), .Q(n32596) );
  and2s1 U24935 ( .DIN1(n32597), .DIN2(n32540), .Q(n32595) );
  or2s1 U24936 ( .DIN1(n32598), .DIN2(n32599), .Q(n9773) );
  and2s1 U24937 ( .DIN1(wb_addr_i[5]), .DIN2(wb_stb_i), .Q(n32599) );
  and2s1 U24938 ( .DIN1(n32600), .DIN2(n32540), .Q(n32598) );
  or2s1 U24939 ( .DIN1(n32601), .DIN2(n32602), .Q(n9772) );
  and2s1 U24940 ( .DIN1(wb_addr_i[4]), .DIN2(wb_stb_i), .Q(n32602) );
  and2s1 U24941 ( .DIN1(n32603), .DIN2(n32540), .Q(n32601) );
  or2s1 U24942 ( .DIN1(n32604), .DIN2(n32605), .Q(n9771) );
  and2s1 U24943 ( .DIN1(wb_addr_i[3]), .DIN2(wb_stb_i), .Q(n32605) );
  and2s1 U24944 ( .DIN1(n32606), .DIN2(n32540), .Q(n32604) );
  or2s1 U24945 ( .DIN1(n32607), .DIN2(n32608), .Q(n9770) );
  and2s1 U24946 ( .DIN1(wb_addr_i[2]), .DIN2(wb_stb_i), .Q(n32608) );
  and2s1 U24947 ( .DIN1(n32609), .DIN2(n32540), .Q(n32607) );
  and2s1 U24948 ( .DIN1(u3_u0_rd_adr[3]), .DIN2(n32610), .Q(n9769) );
  and2s1 U24949 ( .DIN1(u3_u0_rd_adr[2]), .DIN2(n32610), .Q(n9768) );
  and2s1 U24950 ( .DIN1(u3_u0_rd_adr[1]), .DIN2(n32610), .Q(n9767) );
  or2s1 U24951 ( .DIN1(u3_u0_rd_adr[0]), .DIN2(n32611), .Q(n9766) );
  and2s1 U24952 ( .DIN1(n32612), .DIN2(wb_cyc_i), .Q(n9762) );
  and2s1 U24953 ( .DIN1(u5_wb_cycle), .DIN2(n32613), .Q(n32612) );
  or2s1 U24954 ( .DIN1(n32614), .DIN2(n32540), .Q(n32613) );
  and2s1 U24955 ( .DIN1(n32615), .DIN2(wb_cyc_i), .Q(n9761) );
  and2s1 U24956 ( .DIN1(n32616), .DIN2(n4820), .Q(n32615) );
  or2s1 U24957 ( .DIN1(wb_we_i), .DIN2(n32540), .Q(n32616) );
  or2s1 U24958 ( .DIN1(n32617), .DIN2(n32618), .Q(n9760) );
  and2s1 U24959 ( .DIN1(wb_cyc_i), .DIN2(n32619), .Q(n32618) );
  hi1s1 U24960 ( .DIN1(n15472), .Q(n32619) );
  and2s1 U24961 ( .DIN1(n32614), .DIN2(n32032), .Q(n32617) );
  or2s1 U24962 ( .DIN1(n32620), .DIN2(n32032), .Q(n9759) );
  and2s1 U24963 ( .DIN1(n32621), .DIN2(n32622), .Q(n32620) );
  and2s1 U24964 ( .DIN1(n32029), .DIN2(n32623), .Q(n9758) );
  and2s1 U24965 ( .DIN1(n32624), .DIN2(n32625), .Q(n32623) );
  and2s1 U24966 ( .DIN1(n32626), .DIN2(n32034), .Q(n32624) );
  hi1s1 U24967 ( .DIN1(wb_addr_i[31]), .Q(n32034) );
  and2s1 U24968 ( .DIN1(wb_addr_i[30]), .DIN2(wb_addr_i[29]), .Q(n32029) );
  or2s1 U24969 ( .DIN1(n32627), .DIN2(wb_ack_o), .Q(n9757) );
  and2s1 U24970 ( .DIN1(wb_cyc_i), .DIN2(n32628), .Q(n32627) );
  and2s1 U24971 ( .DIN1(n32629), .DIN2(n15514), .Q(n9756) );
  and2s1 U24972 ( .DIN1(n32032), .DIN2(n32628), .Q(n32629) );
  hi1s1 U24973 ( .DIN1(n15471), .Q(n32628) );
  and2s1 U24974 ( .DIN1(n32625), .DIN2(wb_we_i), .Q(n32032) );
  and2s1 U24975 ( .DIN1(n32630), .DIN2(n15475), .Q(n9755) );
  and2s1 U24976 ( .DIN1(n32631), .DIN2(n32632), .Q(n32630) );
  or2s1 U24977 ( .DIN1(n32633), .DIN2(n32634), .Q(n32632) );
  or2s1 U24978 ( .DIN1(n15471), .DIN2(n32622), .Q(n32634) );
  hi1s1 U24979 ( .DIN1(n15514), .Q(n32622) );
  or2s1 U24980 ( .DIN1(n32635), .DIN2(n32636), .Q(n32631) );
  and2s1 U24981 ( .DIN1(wb_cyc_i), .DIN2(n32637), .Q(n32636) );
  hi1s1 U24982 ( .DIN1(n15473), .Q(n32637) );
  and2s1 U24983 ( .DIN1(n32638), .DIN2(n32639), .Q(n32635) );
  or2s1 U24984 ( .DIN1(n32640), .DIN2(n32641), .Q(n9754) );
  and2s1 U24985 ( .DIN1(n32037), .DIN2(n32642), .Q(n32641) );
  and2s1 U24986 ( .DIN1(n32038), .DIN2(n4814), .Q(n32640) );
  hi1s1 U24987 ( .DIN1(n32037), .Q(n32038) );
  or2s1 U24988 ( .DIN1(u0_wb_addr_r[3]), .DIN2(n32139), .Q(n32037) );
  or2s1 U24989 ( .DIN1(n32643), .DIN2(n32644), .Q(n32139) );
  or2s1 U24990 ( .DIN1(n32033), .DIN2(n4975), .Q(n32644) );
  or2s1 U24991 ( .DIN1(u0_wb_addr_r[2]), .DIN2(n32645), .Q(n32643) );
  or2s1 U24992 ( .DIN1(u0_wb_addr_r[6]), .DIN2(u0_wb_addr_r[5]), .Q(n32645) );
  or2s1 U24993 ( .DIN1(n32646), .DIN2(n32647), .Q(n9753) );
  and2s1 U24994 ( .DIN1(poc_o[31]), .DIN2(n15521), .Q(n32647) );
  and2s1 U24995 ( .DIN1(n32648), .DIN2(n32649), .Q(n32646) );
  or2s1 U24996 ( .DIN1(n32650), .DIN2(n32651), .Q(n9752) );
  and2s1 U24997 ( .DIN1(poc_o[30]), .DIN2(n15521), .Q(n32651) );
  and2s1 U24998 ( .DIN1(n32648), .DIN2(n32652), .Q(n32650) );
  or2s1 U24999 ( .DIN1(n32653), .DIN2(n32654), .Q(n9751) );
  and2s1 U25000 ( .DIN1(poc_o[29]), .DIN2(n15521), .Q(n32654) );
  and2s1 U25001 ( .DIN1(n32648), .DIN2(n32655), .Q(n32653) );
  or2s1 U25002 ( .DIN1(n32656), .DIN2(n32657), .Q(n9750) );
  and2s1 U25003 ( .DIN1(poc_o[28]), .DIN2(n15521), .Q(n32657) );
  and2s1 U25004 ( .DIN1(n32648), .DIN2(n32658), .Q(n32656) );
  or2s1 U25005 ( .DIN1(n32659), .DIN2(n32660), .Q(n9749) );
  and2s1 U25006 ( .DIN1(poc_o[27]), .DIN2(n15521), .Q(n32660) );
  and2s1 U25007 ( .DIN1(n32648), .DIN2(n32661), .Q(n32659) );
  or2s1 U25008 ( .DIN1(n32662), .DIN2(n32663), .Q(n9748) );
  and2s1 U25009 ( .DIN1(poc_o[26]), .DIN2(n15521), .Q(n32663) );
  and2s1 U25010 ( .DIN1(n32648), .DIN2(n32664), .Q(n32662) );
  or2s1 U25011 ( .DIN1(n32665), .DIN2(n32666), .Q(n9747) );
  and2s1 U25012 ( .DIN1(poc_o[25]), .DIN2(n15521), .Q(n32666) );
  and2s1 U25013 ( .DIN1(n32648), .DIN2(n32667), .Q(n32665) );
  or2s1 U25014 ( .DIN1(n32668), .DIN2(n32669), .Q(n9746) );
  and2s1 U25015 ( .DIN1(poc_o[24]), .DIN2(n15521), .Q(n32669) );
  and2s1 U25016 ( .DIN1(n32648), .DIN2(n32670), .Q(n32668) );
  or2s1 U25017 ( .DIN1(n32671), .DIN2(n32672), .Q(n9745) );
  and2s1 U25018 ( .DIN1(poc_o[23]), .DIN2(n15521), .Q(n32672) );
  and2s1 U25019 ( .DIN1(n32648), .DIN2(n32673), .Q(n32671) );
  or2s1 U25020 ( .DIN1(n32674), .DIN2(n32675), .Q(n9744) );
  and2s1 U25021 ( .DIN1(poc_o[22]), .DIN2(n15521), .Q(n32675) );
  and2s1 U25022 ( .DIN1(n32648), .DIN2(n32676), .Q(n32674) );
  or2s1 U25023 ( .DIN1(n32677), .DIN2(n32678), .Q(n9743) );
  and2s1 U25024 ( .DIN1(poc_o[21]), .DIN2(n15521), .Q(n32678) );
  and2s1 U25025 ( .DIN1(n32648), .DIN2(n32679), .Q(n32677) );
  or2s1 U25026 ( .DIN1(n32680), .DIN2(n32681), .Q(n9742) );
  and2s1 U25027 ( .DIN1(poc_o[20]), .DIN2(n15521), .Q(n32681) );
  and2s1 U25028 ( .DIN1(n32648), .DIN2(n32682), .Q(n32680) );
  or2s1 U25029 ( .DIN1(n32683), .DIN2(n32684), .Q(n9741) );
  and2s1 U25030 ( .DIN1(poc_o[19]), .DIN2(n15521), .Q(n32684) );
  and2s1 U25031 ( .DIN1(n32648), .DIN2(n32685), .Q(n32683) );
  or2s1 U25032 ( .DIN1(n32686), .DIN2(n32687), .Q(n9740) );
  and2s1 U25033 ( .DIN1(poc_o[18]), .DIN2(n15521), .Q(n32687) );
  and2s1 U25034 ( .DIN1(n32648), .DIN2(n32688), .Q(n32686) );
  or2s1 U25035 ( .DIN1(n32689), .DIN2(n32690), .Q(n9739) );
  and2s1 U25036 ( .DIN1(poc_o[17]), .DIN2(n15521), .Q(n32690) );
  and2s1 U25037 ( .DIN1(n32648), .DIN2(n32691), .Q(n32689) );
  or2s1 U25038 ( .DIN1(n32692), .DIN2(n32693), .Q(n9738) );
  and2s1 U25039 ( .DIN1(poc_o[16]), .DIN2(n15521), .Q(n32693) );
  and2s1 U25040 ( .DIN1(n32648), .DIN2(n32694), .Q(n32692) );
  or2s1 U25041 ( .DIN1(n32695), .DIN2(n32696), .Q(n9737) );
  and2s1 U25042 ( .DIN1(poc_o[15]), .DIN2(n15521), .Q(n32696) );
  and2s1 U25043 ( .DIN1(n32648), .DIN2(n32697), .Q(n32695) );
  or2s1 U25044 ( .DIN1(n32698), .DIN2(n32699), .Q(n9736) );
  and2s1 U25045 ( .DIN1(poc_o[14]), .DIN2(n15521), .Q(n32699) );
  and2s1 U25046 ( .DIN1(n32648), .DIN2(n32700), .Q(n32698) );
  or2s1 U25047 ( .DIN1(n32701), .DIN2(n32702), .Q(n9735) );
  and2s1 U25048 ( .DIN1(poc_o[13]), .DIN2(n15521), .Q(n32702) );
  and2s1 U25049 ( .DIN1(n32648), .DIN2(n32703), .Q(n32701) );
  or2s1 U25050 ( .DIN1(n32704), .DIN2(n32705), .Q(n9734) );
  and2s1 U25051 ( .DIN1(poc_o[12]), .DIN2(n15521), .Q(n32705) );
  and2s1 U25052 ( .DIN1(n32648), .DIN2(n32706), .Q(n32704) );
  or2s1 U25053 ( .DIN1(n32707), .DIN2(n32708), .Q(n9733) );
  and2s1 U25054 ( .DIN1(poc_o[11]), .DIN2(n15521), .Q(n32708) );
  and2s1 U25055 ( .DIN1(n32648), .DIN2(n32709), .Q(n32707) );
  or2s1 U25056 ( .DIN1(n32710), .DIN2(n32711), .Q(n9732) );
  and2s1 U25057 ( .DIN1(poc_o[10]), .DIN2(n15521), .Q(n32711) );
  and2s1 U25058 ( .DIN1(n32648), .DIN2(n32712), .Q(n32710) );
  or2s1 U25059 ( .DIN1(n32713), .DIN2(n32714), .Q(n9731) );
  and2s1 U25060 ( .DIN1(poc_o[9]), .DIN2(n15521), .Q(n32714) );
  and2s1 U25061 ( .DIN1(n32648), .DIN2(n32715), .Q(n32713) );
  or2s1 U25062 ( .DIN1(n32716), .DIN2(n32717), .Q(n9730) );
  and2s1 U25063 ( .DIN1(poc_o[8]), .DIN2(n15521), .Q(n32717) );
  and2s1 U25064 ( .DIN1(n32648), .DIN2(n32718), .Q(n32716) );
  or2s1 U25065 ( .DIN1(n32719), .DIN2(n32720), .Q(n9729) );
  and2s1 U25066 ( .DIN1(poc_o[7]), .DIN2(n15521), .Q(n32720) );
  and2s1 U25067 ( .DIN1(n32648), .DIN2(n32721), .Q(n32719) );
  or2s1 U25068 ( .DIN1(n32722), .DIN2(n32723), .Q(n9728) );
  and2s1 U25069 ( .DIN1(poc_o[6]), .DIN2(n15521), .Q(n32723) );
  and2s1 U25070 ( .DIN1(n32648), .DIN2(n32724), .Q(n32722) );
  or2s1 U25071 ( .DIN1(n32725), .DIN2(n32726), .Q(n9727) );
  and2s1 U25072 ( .DIN1(poc_o[5]), .DIN2(n15521), .Q(n32726) );
  and2s1 U25073 ( .DIN1(n32648), .DIN2(n32727), .Q(n32725) );
  or2s1 U25074 ( .DIN1(n32728), .DIN2(n32729), .Q(n9726) );
  and2s1 U25075 ( .DIN1(poc_o[4]), .DIN2(n15521), .Q(n32729) );
  and2s1 U25076 ( .DIN1(n32648), .DIN2(n32730), .Q(n32728) );
  or2s1 U25077 ( .DIN1(n32731), .DIN2(n32732), .Q(n9725) );
  and2s1 U25078 ( .DIN1(poc_o[3]), .DIN2(n15521), .Q(n32732) );
  and2s1 U25079 ( .DIN1(n32648), .DIN2(n32733), .Q(n32731) );
  or2s1 U25080 ( .DIN1(n32734), .DIN2(n32735), .Q(n9724) );
  or2s1 U25081 ( .DIN1(n32736), .DIN2(n32737), .Q(n32735) );
  and2s1 U25082 ( .DIN1(n32142), .DIN2(wb_data_i[2]), .Q(n32737) );
  and2s1 U25083 ( .DIN1(u0_csc0[2]), .DIN2(n32143), .Q(n32736) );
  and2s1 U25084 ( .DIN1(poc_o[3]), .DIN2(n32213), .Q(n32734) );
  or2s1 U25085 ( .DIN1(n32738), .DIN2(n32739), .Q(n9723) );
  and2s1 U25086 ( .DIN1(poc_o[2]), .DIN2(n15521), .Q(n32739) );
  and2s1 U25087 ( .DIN1(n32648), .DIN2(n32740), .Q(n32738) );
  or2s1 U25088 ( .DIN1(n32741), .DIN2(n32742), .Q(n9722) );
  or2s1 U25089 ( .DIN1(n32743), .DIN2(n32744), .Q(n32742) );
  and2s1 U25090 ( .DIN1(u0_csc0[0]), .DIN2(n32143), .Q(n32744) );
  and2s1 U25091 ( .DIN1(n32745), .DIN2(n32213), .Q(n32743) );
  or2s1 U25092 ( .DIN1(poc_o[2]), .DIN2(poc_o[3]), .Q(n32745) );
  and2s1 U25093 ( .DIN1(n32142), .DIN2(wb_data_i[0]), .Q(n32741) );
  or2s1 U25094 ( .DIN1(n32746), .DIN2(n32747), .Q(n9721) );
  or2s1 U25095 ( .DIN1(n32748), .DIN2(n32749), .Q(n32747) );
  and2s1 U25096 ( .DIN1(n32142), .DIN2(wb_data_i[1]), .Q(n32749) );
  and2s1 U25097 ( .DIN1(n32143), .DIN2(n32750), .Q(n32748) );
  and2s1 U25098 ( .DIN1(poc_o[2]), .DIN2(n32213), .Q(n32746) );
  or2s1 U25099 ( .DIN1(n32751), .DIN2(n32752), .Q(n9720) );
  or2s1 U25100 ( .DIN1(n32753), .DIN2(n32754), .Q(n9719) );
  and2s1 U25101 ( .DIN1(u4_ps_cnt[7]), .DIN2(n32755), .Q(n32754) );
  or2s1 U25102 ( .DIN1(n32756), .DIN2(n32757), .Q(n32755) );
  and2s1 U25103 ( .DIN1(n32758), .DIN2(n32759), .Q(n32756) );
  and2s1 U25104 ( .DIN1(n32760), .DIN2(n32761), .Q(n32753) );
  and2s1 U25105 ( .DIN1(u4_ps_cnt[6]), .DIN2(n32762), .Q(n32760) );
  or2s1 U25106 ( .DIN1(n32763), .DIN2(n32764), .Q(n9718) );
  and2s1 U25107 ( .DIN1(n32765), .DIN2(u4_ps_cnt[0]), .Q(n32763) );
  or2s1 U25108 ( .DIN1(n32766), .DIN2(n32767), .Q(n9717) );
  and2s1 U25109 ( .DIN1(u4_ps_cnt[1]), .DIN2(n32768), .Q(n32767) );
  and2s1 U25110 ( .DIN1(n32769), .DIN2(n32758), .Q(n32766) );
  and2s1 U25111 ( .DIN1(u4_ps_cnt[0]), .DIN2(n32770), .Q(n32769) );
  or2s1 U25112 ( .DIN1(n32771), .DIN2(n32772), .Q(n9716) );
  and2s1 U25113 ( .DIN1(u4_ps_cnt[2]), .DIN2(n32773), .Q(n32772) );
  or2s1 U25114 ( .DIN1(n32774), .DIN2(n32768), .Q(n32773) );
  or2s1 U25115 ( .DIN1(n32764), .DIN2(n32765), .Q(n32768) );
  and2s1 U25116 ( .DIN1(n32758), .DIN2(n32775), .Q(n32764) );
  and2s1 U25117 ( .DIN1(n32758), .DIN2(n32770), .Q(n32774) );
  and2s1 U25118 ( .DIN1(n32776), .DIN2(n32777), .Q(n32771) );
  and2s1 U25119 ( .DIN1(u4_ps_cnt[0]), .DIN2(n32778), .Q(n32777) );
  and2s1 U25120 ( .DIN1(n32758), .DIN2(u4_ps_cnt[1]), .Q(n32776) );
  or2s1 U25121 ( .DIN1(n32779), .DIN2(n32780), .Q(n9715) );
  and2s1 U25122 ( .DIN1(u4_ps_cnt[3]), .DIN2(n32781), .Q(n32780) );
  and2s1 U25123 ( .DIN1(n32782), .DIN2(n32758), .Q(n32779) );
  and2s1 U25124 ( .DIN1(n32783), .DIN2(n32784), .Q(n32782) );
  or2s1 U25125 ( .DIN1(n32785), .DIN2(n32786), .Q(n9714) );
  and2s1 U25126 ( .DIN1(u4_ps_cnt[4]), .DIN2(n32787), .Q(n32786) );
  or2s1 U25127 ( .DIN1(n32788), .DIN2(n32781), .Q(n32787) );
  or2s1 U25128 ( .DIN1(n32789), .DIN2(n32765), .Q(n32781) );
  and2s1 U25129 ( .DIN1(n32758), .DIN2(n32790), .Q(n32789) );
  and2s1 U25130 ( .DIN1(n32758), .DIN2(n32784), .Q(n32788) );
  and2s1 U25131 ( .DIN1(n32791), .DIN2(n32792), .Q(n32785) );
  and2s1 U25132 ( .DIN1(u4_ps_cnt[3]), .DIN2(n32793), .Q(n32792) );
  and2s1 U25133 ( .DIN1(n32758), .DIN2(n32783), .Q(n32791) );
  hi1s1 U25134 ( .DIN1(n32790), .Q(n32783) );
  or2s1 U25135 ( .DIN1(n32794), .DIN2(n32795), .Q(n9713) );
  and2s1 U25136 ( .DIN1(u4_ps_cnt[5]), .DIN2(n32796), .Q(n32795) );
  and2s1 U25137 ( .DIN1(n32797), .DIN2(n32758), .Q(n32794) );
  and2s1 U25138 ( .DIN1(n32798), .DIN2(n32799), .Q(n32797) );
  hi1s1 U25139 ( .DIN1(n32800), .Q(n32798) );
  or2s1 U25140 ( .DIN1(n32801), .DIN2(n32802), .Q(n9712) );
  and2s1 U25141 ( .DIN1(u4_ps_cnt[6]), .DIN2(n32757), .Q(n32802) );
  or2s1 U25142 ( .DIN1(n32803), .DIN2(n32796), .Q(n32757) );
  or2s1 U25143 ( .DIN1(n32804), .DIN2(n32765), .Q(n32796) );
  and2s1 U25144 ( .DIN1(n32805), .DIN2(n32806), .Q(n32765) );
  and2s1 U25145 ( .DIN1(n32758), .DIN2(n32800), .Q(n32804) );
  and2s1 U25146 ( .DIN1(n32758), .DIN2(n32799), .Q(n32803) );
  hi1s1 U25147 ( .DIN1(n32806), .Q(n32758) );
  and2s1 U25148 ( .DIN1(n32761), .DIN2(n32759), .Q(n32801) );
  hi1s1 U25149 ( .DIN1(n32807), .Q(n32761) );
  or2s1 U25150 ( .DIN1(n32806), .DIN2(n32808), .Q(n32807) );
  or2s1 U25151 ( .DIN1(n32799), .DIN2(n32800), .Q(n32808) );
  or2s1 U25152 ( .DIN1(n32790), .DIN2(n32809), .Q(n32800) );
  or2s1 U25153 ( .DIN1(n32793), .DIN2(n32784), .Q(n32809) );
  or2s1 U25154 ( .DIN1(n32770), .DIN2(n32810), .Q(n32790) );
  or2s1 U25155 ( .DIN1(n32778), .DIN2(n32775), .Q(n32810) );
  or2s1 U25156 ( .DIN1(n9711), .DIN2(n4986), .Q(n32806) );
  hi1s1 U25157 ( .DIN1(n32805), .Q(n9711) );
  or2s1 U25158 ( .DIN1(n32811), .DIN2(n32812), .Q(n32805) );
  and2s1 U25159 ( .DIN1(n32813), .DIN2(n32814), .Q(n32811) );
  and2s1 U25160 ( .DIN1(n32815), .DIN2(n32816), .Q(n32814) );
  and2s1 U25161 ( .DIN1(n32817), .DIN2(n32818), .Q(n32816) );
  and2s1 U25162 ( .DIN1(n32819), .DIN2(n32820), .Q(n32815) );
  and2s1 U25163 ( .DIN1(n32821), .DIN2(n32822), .Q(n32813) );
  and2s1 U25164 ( .DIN1(n32823), .DIN2(n32824), .Q(n32822) );
  and2s1 U25165 ( .DIN1(n32825), .DIN2(n32826), .Q(n32821) );
  or2s1 U25166 ( .DIN1(n32827), .DIN2(n32828), .Q(n9710) );
  and2s1 U25167 ( .DIN1(poc_o[1]), .DIN2(n15521), .Q(n32828) );
  and2s1 U25168 ( .DIN1(n32648), .DIN2(n32829), .Q(n32827) );
  or2s1 U25169 ( .DIN1(n32830), .DIN2(n32831), .Q(n9709) );
  or2s1 U25170 ( .DIN1(n32832), .DIN2(n32833), .Q(n32831) );
  and2s1 U25171 ( .DIN1(n32142), .DIN2(wb_data_i[5]), .Q(n32833) );
  and2s1 U25172 ( .DIN1(n32143), .DIN2(n32834), .Q(n32832) );
  and2s1 U25173 ( .DIN1(poc_o[1]), .DIN2(n32213), .Q(n32830) );
  or2s1 U25174 ( .DIN1(n32835), .DIN2(n32836), .Q(n9708) );
  and2s1 U25175 ( .DIN1(poc_o[0]), .DIN2(n15521), .Q(n32836) );
  and2s1 U25176 ( .DIN1(n32648), .DIN2(n32837), .Q(n32835) );
  hi1s1 U25177 ( .DIN1(n15521), .Q(n32648) );
  or2s1 U25178 ( .DIN1(n32838), .DIN2(n32839), .Q(n9707) );
  or2s1 U25179 ( .DIN1(n32840), .DIN2(n32841), .Q(n32839) );
  and2s1 U25180 ( .DIN1(n32142), .DIN2(wb_data_i[4]), .Q(n32841) );
  and2s1 U25181 ( .DIN1(n32143), .DIN2(n32842), .Q(n32840) );
  hi1s1 U25182 ( .DIN1(n32843), .Q(n32143) );
  or2s1 U25183 ( .DIN1(n32142), .DIN2(n32213), .Q(n32843) );
  and2s1 U25184 ( .DIN1(n19405), .DIN2(n15487), .Q(n32142) );
  and2s1 U25185 ( .DIN1(poc_o[0]), .DIN2(n32213), .Q(n32838) );
  hi1s1 U25186 ( .DIN1(n15487), .Q(n32213) );
  and2s1 U25187 ( .DIN1(u5_state[8]), .DIN2(n32844), .Q(n9706) );
  and2s1 U25188 ( .DIN1(u5_state[63]), .DIN2(n32844), .Q(n9705) );
  and2s1 U25189 ( .DIN1(u5_state[60]), .DIN2(n32844), .Q(n9704) );
  and2s1 U25190 ( .DIN1(u5_state[59]), .DIN2(n32844), .Q(n9703) );
  and2s1 U25191 ( .DIN1(u5_state[58]), .DIN2(n32844), .Q(n9702) );
  and2s1 U25192 ( .DIN1(u5_state[56]), .DIN2(n32844), .Q(n9701) );
  and2s1 U25193 ( .DIN1(u5_state[52]), .DIN2(n32844), .Q(n9700) );
  and2s1 U25194 ( .DIN1(u5_state[47]), .DIN2(n32844), .Q(n9699) );
  and2s1 U25195 ( .DIN1(u5_state[36]), .DIN2(n32844), .Q(n9698) );
  and2s1 U25196 ( .DIN1(u5_state[14]), .DIN2(n32844), .Q(n9697) );
  and2s1 U25197 ( .DIN1(u5_state[13]), .DIN2(n32844), .Q(n9696) );
  and2s1 U25198 ( .DIN1(u5_state[0]), .DIN2(n32844), .Q(n9695) );
  or2s1 U25199 ( .DIN1(n32845), .DIN2(n32846), .Q(n9694) );
  and2s1 U25200 ( .DIN1(u5_state[37]), .DIN2(n32844), .Q(n32845) );
  or2s1 U25201 ( .DIN1(n32847), .DIN2(n32848), .Q(n9693) );
  and2s1 U25202 ( .DIN1(u5_state[38]), .DIN2(n32844), .Q(n32848) );
  and2s1 U25203 ( .DIN1(n32849), .DIN2(n32850), .Q(n32847) );
  or2s1 U25204 ( .DIN1(n32851), .DIN2(n32852), .Q(n9692) );
  or2s1 U25205 ( .DIN1(n32853), .DIN2(n32854), .Q(n32852) );
  and2s1 U25206 ( .DIN1(u5_state[39]), .DIN2(n32855), .Q(n32854) );
  and2s1 U25207 ( .DIN1(n32856), .DIN2(u5_tmr2_done), .Q(n32851) );
  or2s1 U25208 ( .DIN1(n32857), .DIN2(n32858), .Q(n9691) );
  and2s1 U25209 ( .DIN1(u5_state[40]), .DIN2(n32844), .Q(n32857) );
  or2s1 U25210 ( .DIN1(n32859), .DIN2(n32860), .Q(n9690) );
  or2s1 U25211 ( .DIN1(n32861), .DIN2(n32862), .Q(n32860) );
  or2s1 U25212 ( .DIN1(n32863), .DIN2(n32864), .Q(n32862) );
  and2s1 U25213 ( .DIN1(n32865), .DIN2(u7_mc_br_r), .Q(n32863) );
  or2s1 U25214 ( .DIN1(n32866), .DIN2(n32867), .Q(n32859) );
  or2s1 U25215 ( .DIN1(n32868), .DIN2(n32869), .Q(n32867) );
  and2s1 U25216 ( .DIN1(n32870), .DIN2(n32871), .Q(n32866) );
  or2s1 U25217 ( .DIN1(n32872), .DIN2(n32873), .Q(n9688) );
  or2s1 U25218 ( .DIN1(n32874), .DIN2(n32875), .Q(n32873) );
  or2s1 U25219 ( .DIN1(n32876), .DIN2(n32877), .Q(n32875) );
  and2s1 U25220 ( .DIN1(n32878), .DIN2(n32879), .Q(n32876) );
  or2s1 U25221 ( .DIN1(n32880), .DIN2(n32881), .Q(n32874) );
  or2s1 U25222 ( .DIN1(n32882), .DIN2(n32883), .Q(n32881) );
  and2s1 U25223 ( .DIN1(n32884), .DIN2(n32885), .Q(n32883) );
  and2s1 U25224 ( .DIN1(n32886), .DIN2(n32887), .Q(n32882) );
  and2s1 U25225 ( .DIN1(n32888), .DIN2(n32889), .Q(n32880) );
  or2s1 U25226 ( .DIN1(n32890), .DIN2(n32891), .Q(n32872) );
  or2s1 U25227 ( .DIN1(n32892), .DIN2(n32893), .Q(n32891) );
  or2s1 U25228 ( .DIN1(n32894), .DIN2(n32895), .Q(n32893) );
  and2s1 U25229 ( .DIN1(n32896), .DIN2(n32897), .Q(n32895) );
  and2s1 U25230 ( .DIN1(n32898), .DIN2(n32899), .Q(n32894) );
  and2s1 U25231 ( .DIN1(n32900), .DIN2(n32901), .Q(n32892) );
  or2s1 U25232 ( .DIN1(n32902), .DIN2(n32903), .Q(n32890) );
  or2s1 U25233 ( .DIN1(n32904), .DIN2(n32905), .Q(n32903) );
  and2s1 U25234 ( .DIN1(n32906), .DIN2(n32907), .Q(n32905) );
  or2s1 U25235 ( .DIN1(n32908), .DIN2(n32909), .Q(n32906) );
  and2s1 U25236 ( .DIN1(n32910), .DIN2(n32911), .Q(n32909) );
  hi1s1 U25237 ( .DIN1(n32912), .Q(n32908) );
  or2s1 U25238 ( .DIN1(n32911), .DIN2(n32910), .Q(n32912) );
  or2s1 U25239 ( .DIN1(n32913), .DIN2(n32914), .Q(n32911) );
  and2s1 U25240 ( .DIN1(n32915), .DIN2(n32916), .Q(n32904) );
  hi1s1 U25241 ( .DIN1(n32917), .Q(n32915) );
  or2s1 U25242 ( .DIN1(u5_timer[0]), .DIN2(u5_timer[1]), .Q(n32917) );
  and2s1 U25243 ( .DIN1(u5_timer[1]), .DIN2(n32918), .Q(n32902) );
  or2s1 U25244 ( .DIN1(n32919), .DIN2(n32920), .Q(n9686) );
  and2s1 U25245 ( .DIN1(n32884), .DIN2(n32921), .Q(n32920) );
  and2s1 U25246 ( .DIN1(u5_state[10]), .DIN2(n32922), .Q(n32919) );
  or2s1 U25247 ( .DIN1(n32923), .DIN2(n32924), .Q(n9685) );
  and2s1 U25248 ( .DIN1(u5_state[11]), .DIN2(n32925), .Q(n32924) );
  and2s1 U25249 ( .DIN1(n32926), .DIN2(n32927), .Q(n32923) );
  and2s1 U25250 ( .DIN1(n32928), .DIN2(n32929), .Q(n32927) );
  and2s1 U25251 ( .DIN1(u5_state[10]), .DIN2(u5_tmr_done), .Q(n32926) );
  or2s1 U25252 ( .DIN1(n32930), .DIN2(n32931), .Q(n9684) );
  or2s1 U25253 ( .DIN1(n32932), .DIN2(n32933), .Q(n32931) );
  and2s1 U25254 ( .DIN1(u5_state[15]), .DIN2(n32844), .Q(n32933) );
  and2s1 U25255 ( .DIN1(n32934), .DIN2(n32935), .Q(n32932) );
  or2s1 U25256 ( .DIN1(n32936), .DIN2(n32937), .Q(n32935) );
  and2s1 U25257 ( .DIN1(n32869), .DIN2(n32938), .Q(n32937) );
  and2s1 U25258 ( .DIN1(n32939), .DIN2(n32940), .Q(n32936) );
  and2s1 U25259 ( .DIN1(n32941), .DIN2(n32921), .Q(n32939) );
  and2s1 U25260 ( .DIN1(n32942), .DIN2(n32943), .Q(n32930) );
  or2s1 U25261 ( .DIN1(n32944), .DIN2(n32945), .Q(n9683) );
  or2s1 U25262 ( .DIN1(n32946), .DIN2(n32947), .Q(n32945) );
  and2s1 U25263 ( .DIN1(n32948), .DIN2(n32949), .Q(n32947) );
  hi1s1 U25264 ( .DIN1(u5_ap_en), .Q(n32949) );
  or2s1 U25265 ( .DIN1(n32950), .DIN2(n32951), .Q(n32948) );
  or2s1 U25266 ( .DIN1(n32952), .DIN2(n32953), .Q(n32951) );
  and2s1 U25267 ( .DIN1(n32954), .DIN2(n32955), .Q(n32953) );
  and2s1 U25268 ( .DIN1(n32956), .DIN2(n32957), .Q(n32955) );
  and2s1 U25269 ( .DIN1(n32958), .DIN2(n32943), .Q(n32954) );
  and2s1 U25270 ( .DIN1(n32959), .DIN2(n32960), .Q(n32950) );
  and2s1 U25271 ( .DIN1(n32961), .DIN2(n32962), .Q(n32959) );
  and2s1 U25272 ( .DIN1(u5_state[16]), .DIN2(n32963), .Q(n32946) );
  or2s1 U25273 ( .DIN1(n32964), .DIN2(n32965), .Q(n32963) );
  and2s1 U25274 ( .DIN1(n15512), .DIN2(n32966), .Q(n32964) );
  and2s1 U25275 ( .DIN1(n32967), .DIN2(n32921), .Q(n32944) );
  or2s1 U25276 ( .DIN1(n32968), .DIN2(n32969), .Q(n9680) );
  and2s1 U25277 ( .DIN1(n32921), .DIN2(n32970), .Q(n32969) );
  and2s1 U25278 ( .DIN1(n9764), .DIN2(n9682), .Q(n32968) );
  or2s1 U25279 ( .DIN1(n32971), .DIN2(n32972), .Q(n9679) );
  and2s1 U25280 ( .DIN1(u5_cmd_asserted2), .DIN2(n32970), .Q(n32972) );
  and2s1 U25281 ( .DIN1(n9764), .DIN2(n32921), .Q(n32971) );
  or2s1 U25282 ( .DIN1(n32973), .DIN2(n32974), .Q(n9678) );
  or2s1 U25283 ( .DIN1(n32975), .DIN2(n32976), .Q(n32974) );
  or2s1 U25284 ( .DIN1(n32977), .DIN2(n32978), .Q(n32976) );
  and2s1 U25285 ( .DIN1(n32865), .DIN2(n32979), .Q(n32978) );
  and2s1 U25286 ( .DIN1(n32952), .DIN2(u5_ap_en), .Q(n32977) );
  hi1s1 U25287 ( .DIN1(n32980), .Q(n32952) );
  or2s1 U25288 ( .DIN1(n32981), .DIN2(n32982), .Q(n32980) );
  or2s1 U25289 ( .DIN1(n32983), .DIN2(n32984), .Q(n32982) );
  or2s1 U25290 ( .DIN1(n15512), .DIN2(n32985), .Q(n32981) );
  and2s1 U25291 ( .DIN1(n32941), .DIN2(n32934), .Q(n32985) );
  or2s1 U25292 ( .DIN1(n32986), .DIN2(n32987), .Q(n32975) );
  and2s1 U25293 ( .DIN1(u5_state[2]), .DIN2(n32988), .Q(n32987) );
  and2s1 U25294 ( .DIN1(n32989), .DIN2(n32921), .Q(n32986) );
  or2s1 U25295 ( .DIN1(n32990), .DIN2(n32991), .Q(n32989) );
  or2s1 U25296 ( .DIN1(n32992), .DIN2(n32993), .Q(n32991) );
  and2s1 U25297 ( .DIN1(n32983), .DIN2(n32940), .Q(n32993) );
  and2s1 U25298 ( .DIN1(u5_wb_cycle), .DIN2(n32957), .Q(n32983) );
  or2s1 U25299 ( .DIN1(n32994), .DIN2(n32995), .Q(n32973) );
  or2s1 U25300 ( .DIN1(n32996), .DIN2(n32997), .Q(n32995) );
  and2s1 U25301 ( .DIN1(n32998), .DIN2(n32943), .Q(n32997) );
  and2s1 U25302 ( .DIN1(n32999), .DIN2(n32956), .Q(n32998) );
  or2s1 U25303 ( .DIN1(n33000), .DIN2(n33001), .Q(n32999) );
  and2s1 U25304 ( .DIN1(u5_ap_en), .DIN2(n32957), .Q(n33000) );
  and2s1 U25305 ( .DIN1(n33002), .DIN2(n33003), .Q(n32996) );
  and2s1 U25306 ( .DIN1(n33004), .DIN2(n33005), .Q(n33003) );
  hi1s1 U25307 ( .DIN1(u5_mem_ack_r), .Q(n33005) );
  and2s1 U25308 ( .DIN1(n32960), .DIN2(n32961), .Q(n33002) );
  or2s1 U25309 ( .DIN1(n33006), .DIN2(n33007), .Q(n32994) );
  and2s1 U25310 ( .DIN1(u5_cke_r), .DIN2(n33008), .Q(n9677) );
  or2s1 U25311 ( .DIN1(n33009), .DIN2(n33010), .Q(n33008) );
  or2s1 U25312 ( .DIN1(n33011), .DIN2(n33012), .Q(n33010) );
  or2s1 U25313 ( .DIN1(n33013), .DIN2(n33014), .Q(n33009) );
  and2s1 U25314 ( .DIN1(n32869), .DIN2(n33015), .Q(n33014) );
  or2s1 U25315 ( .DIN1(n33016), .DIN2(mc_cke_pad_o_), .Q(n33015) );
  and2s1 U25316 ( .DIN1(u5_cnt), .DIN2(n33017), .Q(n33016) );
  or2s1 U25317 ( .DIN1(n33018), .DIN2(n33019), .Q(n9674) );
  and2s1 U25318 ( .DIN1(n33020), .DIN2(n32610), .Q(n33019) );
  and2s1 U25319 ( .DIN1(n33021), .DIN2(n33022), .Q(n33018) );
  or2s1 U25320 ( .DIN1(n32611), .DIN2(n33023), .Q(n9673) );
  or2s1 U25321 ( .DIN1(n33024), .DIN2(n33025), .Q(n33023) );
  and2s1 U25322 ( .DIN1(n36595), .DIN2(n33026), .Q(n33025) );
  hi1s1 U25323 ( .DIN1(n32610), .Q(n32611) );
  or2s1 U25324 ( .DIN1(n33027), .DIN2(n33028), .Q(n9672) );
  and2s1 U25325 ( .DIN1(n33029), .DIN2(n32610), .Q(n33028) );
  and2s1 U25326 ( .DIN1(n33021), .DIN2(n33030), .Q(n33027) );
  or2s1 U25327 ( .DIN1(n33031), .DIN2(n33032), .Q(n9671) );
  and2s1 U25328 ( .DIN1(n33033), .DIN2(n32610), .Q(n33032) );
  and2s1 U25329 ( .DIN1(n33021), .DIN2(n33034), .Q(n33031) );
  and2s1 U25330 ( .DIN1(n33026), .DIN2(n32610), .Q(n33021) );
  and2s1 U25331 ( .DIN1(n32633), .DIN2(wb_cyc_i), .Q(n32610) );
  hi1s1 U25332 ( .DIN1(n33035), .Q(n32633) );
  hi1s1 U25333 ( .DIN1(u5_dv), .Q(n33026) );
  or2s1 U25334 ( .DIN1(n33036), .DIN2(n33037), .Q(n9670) );
  and2s1 U25335 ( .DIN1(n33038), .DIN2(n33039), .Q(n33037) );
  and2s1 U25336 ( .DIN1(n33029), .DIN2(n32837), .Q(n33036) );
  or2s1 U25337 ( .DIN1(n33040), .DIN2(n33041), .Q(n9669) );
  and2s1 U25338 ( .DIN1(n33038), .DIN2(n33042), .Q(n33041) );
  and2s1 U25339 ( .DIN1(n33029), .DIN2(n32829), .Q(n33040) );
  or2s1 U25340 ( .DIN1(n33043), .DIN2(n33044), .Q(n9668) );
  and2s1 U25341 ( .DIN1(n33038), .DIN2(n33045), .Q(n33044) );
  and2s1 U25342 ( .DIN1(n33029), .DIN2(n32740), .Q(n33043) );
  or2s1 U25343 ( .DIN1(n33046), .DIN2(n33047), .Q(n9667) );
  and2s1 U25344 ( .DIN1(n33038), .DIN2(n33048), .Q(n33047) );
  and2s1 U25345 ( .DIN1(n33029), .DIN2(n32733), .Q(n33046) );
  or2s1 U25346 ( .DIN1(n33049), .DIN2(n33050), .Q(n9666) );
  and2s1 U25347 ( .DIN1(n33038), .DIN2(n33051), .Q(n33050) );
  and2s1 U25348 ( .DIN1(n33029), .DIN2(n32730), .Q(n33049) );
  or2s1 U25349 ( .DIN1(n33052), .DIN2(n33053), .Q(n9665) );
  and2s1 U25350 ( .DIN1(n33038), .DIN2(n33054), .Q(n33053) );
  and2s1 U25351 ( .DIN1(n33029), .DIN2(n32727), .Q(n33052) );
  or2s1 U25352 ( .DIN1(n33055), .DIN2(n33056), .Q(n9664) );
  and2s1 U25353 ( .DIN1(n33038), .DIN2(n33057), .Q(n33056) );
  and2s1 U25354 ( .DIN1(n33029), .DIN2(n32724), .Q(n33055) );
  or2s1 U25355 ( .DIN1(n33058), .DIN2(n33059), .Q(n9663) );
  and2s1 U25356 ( .DIN1(n33038), .DIN2(n33060), .Q(n33059) );
  and2s1 U25357 ( .DIN1(n33029), .DIN2(n32721), .Q(n33058) );
  or2s1 U25358 ( .DIN1(n33061), .DIN2(n33062), .Q(n9662) );
  and2s1 U25359 ( .DIN1(n33038), .DIN2(n33063), .Q(n33062) );
  and2s1 U25360 ( .DIN1(n33029), .DIN2(n32718), .Q(n33061) );
  or2s1 U25361 ( .DIN1(n33064), .DIN2(n33065), .Q(n9661) );
  and2s1 U25362 ( .DIN1(n33038), .DIN2(n33066), .Q(n33065) );
  and2s1 U25363 ( .DIN1(n33029), .DIN2(n32715), .Q(n33064) );
  or2s1 U25364 ( .DIN1(n33067), .DIN2(n33068), .Q(n9660) );
  and2s1 U25365 ( .DIN1(n33038), .DIN2(n33069), .Q(n33068) );
  and2s1 U25366 ( .DIN1(n33029), .DIN2(n32712), .Q(n33067) );
  or2s1 U25367 ( .DIN1(n33070), .DIN2(n33071), .Q(n9659) );
  and2s1 U25368 ( .DIN1(n33038), .DIN2(n33072), .Q(n33071) );
  and2s1 U25369 ( .DIN1(n33029), .DIN2(n32709), .Q(n33070) );
  or2s1 U25370 ( .DIN1(n33073), .DIN2(n33074), .Q(n9658) );
  and2s1 U25371 ( .DIN1(n33038), .DIN2(n33075), .Q(n33074) );
  and2s1 U25372 ( .DIN1(n33029), .DIN2(n32706), .Q(n33073) );
  or2s1 U25373 ( .DIN1(n33076), .DIN2(n33077), .Q(n9657) );
  and2s1 U25374 ( .DIN1(n33038), .DIN2(n33078), .Q(n33077) );
  and2s1 U25375 ( .DIN1(n33029), .DIN2(n32703), .Q(n33076) );
  or2s1 U25376 ( .DIN1(n33079), .DIN2(n33080), .Q(n9656) );
  and2s1 U25377 ( .DIN1(n33038), .DIN2(n33081), .Q(n33080) );
  and2s1 U25378 ( .DIN1(n33029), .DIN2(n32700), .Q(n33079) );
  or2s1 U25379 ( .DIN1(n33082), .DIN2(n33083), .Q(n9655) );
  and2s1 U25380 ( .DIN1(n33038), .DIN2(n33084), .Q(n33083) );
  and2s1 U25381 ( .DIN1(n33029), .DIN2(n32697), .Q(n33082) );
  or2s1 U25382 ( .DIN1(n33085), .DIN2(n33086), .Q(n9654) );
  and2s1 U25383 ( .DIN1(n33038), .DIN2(n33087), .Q(n33086) );
  and2s1 U25384 ( .DIN1(n33029), .DIN2(n32694), .Q(n33085) );
  or2s1 U25385 ( .DIN1(n33088), .DIN2(n33089), .Q(n9653) );
  and2s1 U25386 ( .DIN1(n33038), .DIN2(n33090), .Q(n33089) );
  and2s1 U25387 ( .DIN1(n33029), .DIN2(n32691), .Q(n33088) );
  or2s1 U25388 ( .DIN1(n33091), .DIN2(n33092), .Q(n9652) );
  and2s1 U25389 ( .DIN1(n33038), .DIN2(n33093), .Q(n33092) );
  and2s1 U25390 ( .DIN1(n33029), .DIN2(n32688), .Q(n33091) );
  or2s1 U25391 ( .DIN1(n33094), .DIN2(n33095), .Q(n9651) );
  and2s1 U25392 ( .DIN1(n33038), .DIN2(n33096), .Q(n33095) );
  and2s1 U25393 ( .DIN1(n33029), .DIN2(n32685), .Q(n33094) );
  or2s1 U25394 ( .DIN1(n33097), .DIN2(n33098), .Q(n9650) );
  and2s1 U25395 ( .DIN1(n33038), .DIN2(n33099), .Q(n33098) );
  and2s1 U25396 ( .DIN1(n33029), .DIN2(n32682), .Q(n33097) );
  or2s1 U25397 ( .DIN1(n33100), .DIN2(n33101), .Q(n9649) );
  and2s1 U25398 ( .DIN1(n33038), .DIN2(n33102), .Q(n33101) );
  and2s1 U25399 ( .DIN1(n33029), .DIN2(n32679), .Q(n33100) );
  or2s1 U25400 ( .DIN1(n33103), .DIN2(n33104), .Q(n9648) );
  and2s1 U25401 ( .DIN1(n33038), .DIN2(n33105), .Q(n33104) );
  and2s1 U25402 ( .DIN1(n33029), .DIN2(n32676), .Q(n33103) );
  or2s1 U25403 ( .DIN1(n33106), .DIN2(n33107), .Q(n9647) );
  and2s1 U25404 ( .DIN1(n33038), .DIN2(n33108), .Q(n33107) );
  and2s1 U25405 ( .DIN1(n33029), .DIN2(n32673), .Q(n33106) );
  or2s1 U25406 ( .DIN1(n33109), .DIN2(n33110), .Q(n9646) );
  and2s1 U25407 ( .DIN1(n33038), .DIN2(n33111), .Q(n33110) );
  and2s1 U25408 ( .DIN1(n33029), .DIN2(n32670), .Q(n33109) );
  or2s1 U25409 ( .DIN1(n33112), .DIN2(n33113), .Q(n9645) );
  and2s1 U25410 ( .DIN1(n33038), .DIN2(n33114), .Q(n33113) );
  and2s1 U25411 ( .DIN1(n33029), .DIN2(n32667), .Q(n33112) );
  or2s1 U25412 ( .DIN1(n33115), .DIN2(n33116), .Q(n9644) );
  and2s1 U25413 ( .DIN1(n33038), .DIN2(n33117), .Q(n33116) );
  and2s1 U25414 ( .DIN1(n33029), .DIN2(n32664), .Q(n33115) );
  or2s1 U25415 ( .DIN1(n33118), .DIN2(n33119), .Q(n9643) );
  and2s1 U25416 ( .DIN1(n33038), .DIN2(n33120), .Q(n33119) );
  and2s1 U25417 ( .DIN1(n33029), .DIN2(n32661), .Q(n33118) );
  or2s1 U25418 ( .DIN1(n33121), .DIN2(n33122), .Q(n9642) );
  and2s1 U25419 ( .DIN1(n33038), .DIN2(n33123), .Q(n33122) );
  and2s1 U25420 ( .DIN1(n33029), .DIN2(n32658), .Q(n33121) );
  or2s1 U25421 ( .DIN1(n33124), .DIN2(n33125), .Q(n9641) );
  and2s1 U25422 ( .DIN1(n33038), .DIN2(n33126), .Q(n33125) );
  and2s1 U25423 ( .DIN1(n33029), .DIN2(n32655), .Q(n33124) );
  or2s1 U25424 ( .DIN1(n33127), .DIN2(n33128), .Q(n9640) );
  and2s1 U25425 ( .DIN1(n33038), .DIN2(n33129), .Q(n33128) );
  and2s1 U25426 ( .DIN1(n33029), .DIN2(n32652), .Q(n33127) );
  or2s1 U25427 ( .DIN1(n33130), .DIN2(n33131), .Q(n9639) );
  and2s1 U25428 ( .DIN1(n33038), .DIN2(n33132), .Q(n33131) );
  hi1s1 U25429 ( .DIN1(n33029), .Q(n33038) );
  and2s1 U25430 ( .DIN1(n33029), .DIN2(n32649), .Q(n33130) );
  and2s1 U25431 ( .DIN1(u5_dv), .DIN2(n36595), .Q(n33029) );
  or2s1 U25432 ( .DIN1(n33133), .DIN2(n33134), .Q(n9638) );
  and2s1 U25433 ( .DIN1(n33135), .DIN2(n33136), .Q(n33134) );
  and2s1 U25434 ( .DIN1(n33033), .DIN2(n32837), .Q(n33133) );
  or2s1 U25435 ( .DIN1(n33137), .DIN2(n33138), .Q(n9637) );
  and2s1 U25436 ( .DIN1(n33135), .DIN2(n33139), .Q(n33138) );
  and2s1 U25437 ( .DIN1(n33033), .DIN2(n32829), .Q(n33137) );
  or2s1 U25438 ( .DIN1(n33140), .DIN2(n33141), .Q(n9636) );
  and2s1 U25439 ( .DIN1(n33135), .DIN2(n33142), .Q(n33141) );
  and2s1 U25440 ( .DIN1(n33033), .DIN2(n32740), .Q(n33140) );
  or2s1 U25441 ( .DIN1(n33143), .DIN2(n33144), .Q(n9635) );
  and2s1 U25442 ( .DIN1(n33135), .DIN2(n33145), .Q(n33144) );
  and2s1 U25443 ( .DIN1(n33033), .DIN2(n32733), .Q(n33143) );
  or2s1 U25444 ( .DIN1(n33146), .DIN2(n33147), .Q(n9634) );
  and2s1 U25445 ( .DIN1(n33135), .DIN2(n33148), .Q(n33147) );
  and2s1 U25446 ( .DIN1(n33033), .DIN2(n32730), .Q(n33146) );
  or2s1 U25447 ( .DIN1(n33149), .DIN2(n33150), .Q(n9633) );
  and2s1 U25448 ( .DIN1(n33135), .DIN2(n33151), .Q(n33150) );
  and2s1 U25449 ( .DIN1(n33033), .DIN2(n32727), .Q(n33149) );
  or2s1 U25450 ( .DIN1(n33152), .DIN2(n33153), .Q(n9632) );
  and2s1 U25451 ( .DIN1(n33135), .DIN2(n33154), .Q(n33153) );
  and2s1 U25452 ( .DIN1(n33033), .DIN2(n32724), .Q(n33152) );
  or2s1 U25453 ( .DIN1(n33155), .DIN2(n33156), .Q(n9631) );
  and2s1 U25454 ( .DIN1(n33135), .DIN2(n33157), .Q(n33156) );
  and2s1 U25455 ( .DIN1(n33033), .DIN2(n32721), .Q(n33155) );
  or2s1 U25456 ( .DIN1(n33158), .DIN2(n33159), .Q(n9630) );
  and2s1 U25457 ( .DIN1(n33135), .DIN2(n33160), .Q(n33159) );
  and2s1 U25458 ( .DIN1(n33033), .DIN2(n32718), .Q(n33158) );
  or2s1 U25459 ( .DIN1(n33161), .DIN2(n33162), .Q(n9629) );
  and2s1 U25460 ( .DIN1(n33135), .DIN2(n33163), .Q(n33162) );
  and2s1 U25461 ( .DIN1(n33033), .DIN2(n32715), .Q(n33161) );
  or2s1 U25462 ( .DIN1(n33164), .DIN2(n33165), .Q(n9628) );
  and2s1 U25463 ( .DIN1(n33135), .DIN2(n33166), .Q(n33165) );
  and2s1 U25464 ( .DIN1(n33033), .DIN2(n32712), .Q(n33164) );
  or2s1 U25465 ( .DIN1(n33167), .DIN2(n33168), .Q(n9627) );
  and2s1 U25466 ( .DIN1(n33135), .DIN2(n33169), .Q(n33168) );
  and2s1 U25467 ( .DIN1(n33033), .DIN2(n32709), .Q(n33167) );
  or2s1 U25468 ( .DIN1(n33170), .DIN2(n33171), .Q(n9626) );
  and2s1 U25469 ( .DIN1(n33135), .DIN2(n33172), .Q(n33171) );
  and2s1 U25470 ( .DIN1(n33033), .DIN2(n32706), .Q(n33170) );
  or2s1 U25471 ( .DIN1(n33173), .DIN2(n33174), .Q(n9625) );
  and2s1 U25472 ( .DIN1(n33135), .DIN2(n33175), .Q(n33174) );
  and2s1 U25473 ( .DIN1(n33033), .DIN2(n32703), .Q(n33173) );
  or2s1 U25474 ( .DIN1(n33176), .DIN2(n33177), .Q(n9624) );
  and2s1 U25475 ( .DIN1(n33135), .DIN2(n33178), .Q(n33177) );
  and2s1 U25476 ( .DIN1(n33033), .DIN2(n32700), .Q(n33176) );
  or2s1 U25477 ( .DIN1(n33179), .DIN2(n33180), .Q(n9623) );
  and2s1 U25478 ( .DIN1(n33135), .DIN2(n33181), .Q(n33180) );
  and2s1 U25479 ( .DIN1(n33033), .DIN2(n32697), .Q(n33179) );
  or2s1 U25480 ( .DIN1(n33182), .DIN2(n33183), .Q(n9622) );
  and2s1 U25481 ( .DIN1(n33135), .DIN2(n33184), .Q(n33183) );
  and2s1 U25482 ( .DIN1(n33033), .DIN2(n32694), .Q(n33182) );
  or2s1 U25483 ( .DIN1(n33185), .DIN2(n33186), .Q(n9621) );
  and2s1 U25484 ( .DIN1(n33135), .DIN2(n33187), .Q(n33186) );
  and2s1 U25485 ( .DIN1(n33033), .DIN2(n32691), .Q(n33185) );
  or2s1 U25486 ( .DIN1(n33188), .DIN2(n33189), .Q(n9620) );
  and2s1 U25487 ( .DIN1(n33135), .DIN2(n33190), .Q(n33189) );
  and2s1 U25488 ( .DIN1(n33033), .DIN2(n32688), .Q(n33188) );
  or2s1 U25489 ( .DIN1(n33191), .DIN2(n33192), .Q(n9619) );
  and2s1 U25490 ( .DIN1(n33135), .DIN2(n33193), .Q(n33192) );
  and2s1 U25491 ( .DIN1(n33033), .DIN2(n32685), .Q(n33191) );
  or2s1 U25492 ( .DIN1(n33194), .DIN2(n33195), .Q(n9618) );
  and2s1 U25493 ( .DIN1(n33135), .DIN2(n33196), .Q(n33195) );
  and2s1 U25494 ( .DIN1(n33033), .DIN2(n32682), .Q(n33194) );
  or2s1 U25495 ( .DIN1(n33197), .DIN2(n33198), .Q(n9617) );
  and2s1 U25496 ( .DIN1(n33135), .DIN2(n33199), .Q(n33198) );
  and2s1 U25497 ( .DIN1(n33033), .DIN2(n32679), .Q(n33197) );
  or2s1 U25498 ( .DIN1(n33200), .DIN2(n33201), .Q(n9616) );
  and2s1 U25499 ( .DIN1(n33135), .DIN2(n33202), .Q(n33201) );
  and2s1 U25500 ( .DIN1(n33033), .DIN2(n32676), .Q(n33200) );
  or2s1 U25501 ( .DIN1(n33203), .DIN2(n33204), .Q(n9615) );
  and2s1 U25502 ( .DIN1(n33135), .DIN2(n33205), .Q(n33204) );
  and2s1 U25503 ( .DIN1(n33033), .DIN2(n32673), .Q(n33203) );
  or2s1 U25504 ( .DIN1(n33206), .DIN2(n33207), .Q(n9614) );
  and2s1 U25505 ( .DIN1(n33135), .DIN2(n33208), .Q(n33207) );
  and2s1 U25506 ( .DIN1(n33033), .DIN2(n32670), .Q(n33206) );
  or2s1 U25507 ( .DIN1(n33209), .DIN2(n33210), .Q(n9613) );
  and2s1 U25508 ( .DIN1(n33135), .DIN2(n33211), .Q(n33210) );
  and2s1 U25509 ( .DIN1(n33033), .DIN2(n32667), .Q(n33209) );
  or2s1 U25510 ( .DIN1(n33212), .DIN2(n33213), .Q(n9612) );
  and2s1 U25511 ( .DIN1(n33135), .DIN2(n33214), .Q(n33213) );
  and2s1 U25512 ( .DIN1(n33033), .DIN2(n32664), .Q(n33212) );
  or2s1 U25513 ( .DIN1(n33215), .DIN2(n33216), .Q(n9611) );
  and2s1 U25514 ( .DIN1(n33135), .DIN2(n33217), .Q(n33216) );
  and2s1 U25515 ( .DIN1(n33033), .DIN2(n32661), .Q(n33215) );
  or2s1 U25516 ( .DIN1(n33218), .DIN2(n33219), .Q(n9610) );
  and2s1 U25517 ( .DIN1(n33135), .DIN2(n33220), .Q(n33219) );
  and2s1 U25518 ( .DIN1(n33033), .DIN2(n32658), .Q(n33218) );
  or2s1 U25519 ( .DIN1(n33221), .DIN2(n33222), .Q(n9609) );
  and2s1 U25520 ( .DIN1(n33135), .DIN2(n33223), .Q(n33222) );
  and2s1 U25521 ( .DIN1(n33033), .DIN2(n32655), .Q(n33221) );
  or2s1 U25522 ( .DIN1(n33224), .DIN2(n33225), .Q(n9608) );
  and2s1 U25523 ( .DIN1(n33135), .DIN2(n33226), .Q(n33225) );
  and2s1 U25524 ( .DIN1(n33033), .DIN2(n32652), .Q(n33224) );
  or2s1 U25525 ( .DIN1(n33227), .DIN2(n33228), .Q(n9607) );
  and2s1 U25526 ( .DIN1(n33135), .DIN2(n33229), .Q(n33228) );
  hi1s1 U25527 ( .DIN1(n33033), .Q(n33135) );
  and2s1 U25528 ( .DIN1(n33033), .DIN2(n32649), .Q(n33227) );
  and2s1 U25529 ( .DIN1(u5_dv), .DIN2(n33030), .Q(n33033) );
  hi1s1 U25530 ( .DIN1(n15479), .Q(n33030) );
  or2s1 U25531 ( .DIN1(n33230), .DIN2(n33231), .Q(n9606) );
  and2s1 U25532 ( .DIN1(n33232), .DIN2(n33233), .Q(n33231) );
  and2s1 U25533 ( .DIN1(n33020), .DIN2(n32837), .Q(n33230) );
  or2s1 U25534 ( .DIN1(n33234), .DIN2(n33235), .Q(n9605) );
  and2s1 U25535 ( .DIN1(n33232), .DIN2(n33236), .Q(n33235) );
  and2s1 U25536 ( .DIN1(n33020), .DIN2(n32829), .Q(n33234) );
  or2s1 U25537 ( .DIN1(n33237), .DIN2(n33238), .Q(n9604) );
  and2s1 U25538 ( .DIN1(n33232), .DIN2(n33239), .Q(n33238) );
  and2s1 U25539 ( .DIN1(n33020), .DIN2(n32740), .Q(n33237) );
  or2s1 U25540 ( .DIN1(n33240), .DIN2(n33241), .Q(n9603) );
  and2s1 U25541 ( .DIN1(n33232), .DIN2(n33242), .Q(n33241) );
  and2s1 U25542 ( .DIN1(n33020), .DIN2(n32733), .Q(n33240) );
  or2s1 U25543 ( .DIN1(n33243), .DIN2(n33244), .Q(n9602) );
  and2s1 U25544 ( .DIN1(n33232), .DIN2(n33245), .Q(n33244) );
  and2s1 U25545 ( .DIN1(n33020), .DIN2(n32730), .Q(n33243) );
  or2s1 U25546 ( .DIN1(n33246), .DIN2(n33247), .Q(n9601) );
  and2s1 U25547 ( .DIN1(n33232), .DIN2(n33248), .Q(n33247) );
  and2s1 U25548 ( .DIN1(n33020), .DIN2(n32727), .Q(n33246) );
  or2s1 U25549 ( .DIN1(n33249), .DIN2(n33250), .Q(n9600) );
  and2s1 U25550 ( .DIN1(n33232), .DIN2(n33251), .Q(n33250) );
  and2s1 U25551 ( .DIN1(n33020), .DIN2(n32724), .Q(n33249) );
  or2s1 U25552 ( .DIN1(n33252), .DIN2(n33253), .Q(n9599) );
  and2s1 U25553 ( .DIN1(n33232), .DIN2(n33254), .Q(n33253) );
  and2s1 U25554 ( .DIN1(n33020), .DIN2(n32721), .Q(n33252) );
  or2s1 U25555 ( .DIN1(n33255), .DIN2(n33256), .Q(n9598) );
  and2s1 U25556 ( .DIN1(n33232), .DIN2(n33257), .Q(n33256) );
  and2s1 U25557 ( .DIN1(n33020), .DIN2(n32718), .Q(n33255) );
  or2s1 U25558 ( .DIN1(n33258), .DIN2(n33259), .Q(n9597) );
  and2s1 U25559 ( .DIN1(n33232), .DIN2(n33260), .Q(n33259) );
  and2s1 U25560 ( .DIN1(n33020), .DIN2(n32715), .Q(n33258) );
  or2s1 U25561 ( .DIN1(n33261), .DIN2(n33262), .Q(n9596) );
  and2s1 U25562 ( .DIN1(n33232), .DIN2(n33263), .Q(n33262) );
  and2s1 U25563 ( .DIN1(n33020), .DIN2(n32712), .Q(n33261) );
  or2s1 U25564 ( .DIN1(n33264), .DIN2(n33265), .Q(n9595) );
  and2s1 U25565 ( .DIN1(n33232), .DIN2(n33266), .Q(n33265) );
  and2s1 U25566 ( .DIN1(n33020), .DIN2(n32709), .Q(n33264) );
  or2s1 U25567 ( .DIN1(n33267), .DIN2(n33268), .Q(n9594) );
  and2s1 U25568 ( .DIN1(n33232), .DIN2(n33269), .Q(n33268) );
  and2s1 U25569 ( .DIN1(n33020), .DIN2(n32706), .Q(n33267) );
  or2s1 U25570 ( .DIN1(n33270), .DIN2(n33271), .Q(n9593) );
  and2s1 U25571 ( .DIN1(n33232), .DIN2(n33272), .Q(n33271) );
  and2s1 U25572 ( .DIN1(n33020), .DIN2(n32703), .Q(n33270) );
  or2s1 U25573 ( .DIN1(n33273), .DIN2(n33274), .Q(n9592) );
  and2s1 U25574 ( .DIN1(n33232), .DIN2(n33275), .Q(n33274) );
  and2s1 U25575 ( .DIN1(n33020), .DIN2(n32700), .Q(n33273) );
  or2s1 U25576 ( .DIN1(n33276), .DIN2(n33277), .Q(n9591) );
  and2s1 U25577 ( .DIN1(n33232), .DIN2(n33278), .Q(n33277) );
  and2s1 U25578 ( .DIN1(n33020), .DIN2(n32697), .Q(n33276) );
  or2s1 U25579 ( .DIN1(n33279), .DIN2(n33280), .Q(n9590) );
  and2s1 U25580 ( .DIN1(n33232), .DIN2(n33281), .Q(n33280) );
  and2s1 U25581 ( .DIN1(n33020), .DIN2(n32694), .Q(n33279) );
  or2s1 U25582 ( .DIN1(n33282), .DIN2(n33283), .Q(n9589) );
  and2s1 U25583 ( .DIN1(n33232), .DIN2(n33284), .Q(n33283) );
  and2s1 U25584 ( .DIN1(n33020), .DIN2(n32691), .Q(n33282) );
  or2s1 U25585 ( .DIN1(n33285), .DIN2(n33286), .Q(n9588) );
  and2s1 U25586 ( .DIN1(n33232), .DIN2(n33287), .Q(n33286) );
  and2s1 U25587 ( .DIN1(n33020), .DIN2(n32688), .Q(n33285) );
  or2s1 U25588 ( .DIN1(n33288), .DIN2(n33289), .Q(n9587) );
  and2s1 U25589 ( .DIN1(n33232), .DIN2(n33290), .Q(n33289) );
  and2s1 U25590 ( .DIN1(n33020), .DIN2(n32685), .Q(n33288) );
  or2s1 U25591 ( .DIN1(n33291), .DIN2(n33292), .Q(n9586) );
  and2s1 U25592 ( .DIN1(n33232), .DIN2(n33293), .Q(n33292) );
  and2s1 U25593 ( .DIN1(n33020), .DIN2(n32682), .Q(n33291) );
  or2s1 U25594 ( .DIN1(n33294), .DIN2(n33295), .Q(n9585) );
  and2s1 U25595 ( .DIN1(n33232), .DIN2(n33296), .Q(n33295) );
  and2s1 U25596 ( .DIN1(n33020), .DIN2(n32679), .Q(n33294) );
  or2s1 U25597 ( .DIN1(n33297), .DIN2(n33298), .Q(n9584) );
  and2s1 U25598 ( .DIN1(n33232), .DIN2(n33299), .Q(n33298) );
  and2s1 U25599 ( .DIN1(n33020), .DIN2(n32676), .Q(n33297) );
  or2s1 U25600 ( .DIN1(n33300), .DIN2(n33301), .Q(n9583) );
  and2s1 U25601 ( .DIN1(n33232), .DIN2(n33302), .Q(n33301) );
  and2s1 U25602 ( .DIN1(n33020), .DIN2(n32673), .Q(n33300) );
  or2s1 U25603 ( .DIN1(n33303), .DIN2(n33304), .Q(n9582) );
  and2s1 U25604 ( .DIN1(n33232), .DIN2(n33305), .Q(n33304) );
  and2s1 U25605 ( .DIN1(n33020), .DIN2(n32670), .Q(n33303) );
  or2s1 U25606 ( .DIN1(n33306), .DIN2(n33307), .Q(n9581) );
  and2s1 U25607 ( .DIN1(n33232), .DIN2(n33308), .Q(n33307) );
  and2s1 U25608 ( .DIN1(n33020), .DIN2(n32667), .Q(n33306) );
  or2s1 U25609 ( .DIN1(n33309), .DIN2(n33310), .Q(n9580) );
  and2s1 U25610 ( .DIN1(n33232), .DIN2(n33311), .Q(n33310) );
  and2s1 U25611 ( .DIN1(n33020), .DIN2(n32664), .Q(n33309) );
  or2s1 U25612 ( .DIN1(n33312), .DIN2(n33313), .Q(n9579) );
  and2s1 U25613 ( .DIN1(n33232), .DIN2(n33314), .Q(n33313) );
  and2s1 U25614 ( .DIN1(n33020), .DIN2(n32661), .Q(n33312) );
  or2s1 U25615 ( .DIN1(n33315), .DIN2(n33316), .Q(n9578) );
  and2s1 U25616 ( .DIN1(n33232), .DIN2(n33317), .Q(n33316) );
  and2s1 U25617 ( .DIN1(n33020), .DIN2(n32658), .Q(n33315) );
  or2s1 U25618 ( .DIN1(n33318), .DIN2(n33319), .Q(n9577) );
  and2s1 U25619 ( .DIN1(n33232), .DIN2(n33320), .Q(n33319) );
  and2s1 U25620 ( .DIN1(n33020), .DIN2(n32655), .Q(n33318) );
  or2s1 U25621 ( .DIN1(n33321), .DIN2(n33322), .Q(n9576) );
  and2s1 U25622 ( .DIN1(n33232), .DIN2(n33323), .Q(n33322) );
  and2s1 U25623 ( .DIN1(n33020), .DIN2(n32652), .Q(n33321) );
  or2s1 U25624 ( .DIN1(n33324), .DIN2(n33325), .Q(n9575) );
  and2s1 U25625 ( .DIN1(n33232), .DIN2(n33326), .Q(n33325) );
  hi1s1 U25626 ( .DIN1(n33020), .Q(n33232) );
  and2s1 U25627 ( .DIN1(n33020), .DIN2(n32649), .Q(n33324) );
  and2s1 U25628 ( .DIN1(u5_dv), .DIN2(n33034), .Q(n33020) );
  hi1s1 U25629 ( .DIN1(n15478), .Q(n33034) );
  or2s1 U25630 ( .DIN1(n33327), .DIN2(n33328), .Q(n9574) );
  and2s1 U25631 ( .DIN1(n33329), .DIN2(n33330), .Q(n33328) );
  and2s1 U25632 ( .DIN1(n33024), .DIN2(n32837), .Q(n33327) );
  or2s1 U25633 ( .DIN1(n33331), .DIN2(n33332), .Q(n9573) );
  and2s1 U25634 ( .DIN1(n33329), .DIN2(n33333), .Q(n33332) );
  and2s1 U25635 ( .DIN1(n33024), .DIN2(n32829), .Q(n33331) );
  or2s1 U25636 ( .DIN1(n33334), .DIN2(n33335), .Q(n9572) );
  and2s1 U25637 ( .DIN1(n33329), .DIN2(n33336), .Q(n33335) );
  and2s1 U25638 ( .DIN1(n33024), .DIN2(n32740), .Q(n33334) );
  or2s1 U25639 ( .DIN1(n33337), .DIN2(n33338), .Q(n9571) );
  and2s1 U25640 ( .DIN1(n33329), .DIN2(n33339), .Q(n33338) );
  and2s1 U25641 ( .DIN1(n33024), .DIN2(n32733), .Q(n33337) );
  or2s1 U25642 ( .DIN1(n33340), .DIN2(n33341), .Q(n9570) );
  and2s1 U25643 ( .DIN1(n33329), .DIN2(n33342), .Q(n33341) );
  and2s1 U25644 ( .DIN1(n33024), .DIN2(n32730), .Q(n33340) );
  or2s1 U25645 ( .DIN1(n33343), .DIN2(n33344), .Q(n9569) );
  and2s1 U25646 ( .DIN1(n33329), .DIN2(n33345), .Q(n33344) );
  and2s1 U25647 ( .DIN1(n33024), .DIN2(n32727), .Q(n33343) );
  or2s1 U25648 ( .DIN1(n33346), .DIN2(n33347), .Q(n9568) );
  and2s1 U25649 ( .DIN1(n33329), .DIN2(n33348), .Q(n33347) );
  and2s1 U25650 ( .DIN1(n33024), .DIN2(n32724), .Q(n33346) );
  or2s1 U25651 ( .DIN1(n33349), .DIN2(n33350), .Q(n9567) );
  and2s1 U25652 ( .DIN1(n33329), .DIN2(n33351), .Q(n33350) );
  and2s1 U25653 ( .DIN1(n33024), .DIN2(n32721), .Q(n33349) );
  or2s1 U25654 ( .DIN1(n33352), .DIN2(n33353), .Q(n9566) );
  and2s1 U25655 ( .DIN1(n33329), .DIN2(n33354), .Q(n33353) );
  and2s1 U25656 ( .DIN1(n33024), .DIN2(n32718), .Q(n33352) );
  or2s1 U25657 ( .DIN1(n33355), .DIN2(n33356), .Q(n9565) );
  and2s1 U25658 ( .DIN1(n33329), .DIN2(n33357), .Q(n33356) );
  and2s1 U25659 ( .DIN1(n33024), .DIN2(n32715), .Q(n33355) );
  or2s1 U25660 ( .DIN1(n33358), .DIN2(n33359), .Q(n9564) );
  and2s1 U25661 ( .DIN1(n33329), .DIN2(n33360), .Q(n33359) );
  and2s1 U25662 ( .DIN1(n33024), .DIN2(n32712), .Q(n33358) );
  or2s1 U25663 ( .DIN1(n33361), .DIN2(n33362), .Q(n9563) );
  and2s1 U25664 ( .DIN1(n33329), .DIN2(n33363), .Q(n33362) );
  and2s1 U25665 ( .DIN1(n33024), .DIN2(n32709), .Q(n33361) );
  or2s1 U25666 ( .DIN1(n33364), .DIN2(n33365), .Q(n9562) );
  and2s1 U25667 ( .DIN1(n33329), .DIN2(n33366), .Q(n33365) );
  and2s1 U25668 ( .DIN1(n33024), .DIN2(n32706), .Q(n33364) );
  or2s1 U25669 ( .DIN1(n33367), .DIN2(n33368), .Q(n9561) );
  and2s1 U25670 ( .DIN1(n33329), .DIN2(n33369), .Q(n33368) );
  and2s1 U25671 ( .DIN1(n33024), .DIN2(n32703), .Q(n33367) );
  or2s1 U25672 ( .DIN1(n33370), .DIN2(n33371), .Q(n9560) );
  and2s1 U25673 ( .DIN1(n33329), .DIN2(n33372), .Q(n33371) );
  and2s1 U25674 ( .DIN1(n33024), .DIN2(n32700), .Q(n33370) );
  or2s1 U25675 ( .DIN1(n33373), .DIN2(n33374), .Q(n9559) );
  and2s1 U25676 ( .DIN1(n33329), .DIN2(n33375), .Q(n33374) );
  and2s1 U25677 ( .DIN1(n33024), .DIN2(n32697), .Q(n33373) );
  or2s1 U25678 ( .DIN1(n33376), .DIN2(n33377), .Q(n9558) );
  and2s1 U25679 ( .DIN1(n33329), .DIN2(n33378), .Q(n33377) );
  and2s1 U25680 ( .DIN1(n33024), .DIN2(n32694), .Q(n33376) );
  or2s1 U25681 ( .DIN1(n33379), .DIN2(n33380), .Q(n9557) );
  and2s1 U25682 ( .DIN1(n33329), .DIN2(n33381), .Q(n33380) );
  and2s1 U25683 ( .DIN1(n33024), .DIN2(n32691), .Q(n33379) );
  or2s1 U25684 ( .DIN1(n33382), .DIN2(n33383), .Q(n9556) );
  and2s1 U25685 ( .DIN1(n33329), .DIN2(n33384), .Q(n33383) );
  and2s1 U25686 ( .DIN1(n33024), .DIN2(n32688), .Q(n33382) );
  or2s1 U25687 ( .DIN1(n33385), .DIN2(n33386), .Q(n9555) );
  and2s1 U25688 ( .DIN1(n33329), .DIN2(n33387), .Q(n33386) );
  and2s1 U25689 ( .DIN1(n33024), .DIN2(n32685), .Q(n33385) );
  or2s1 U25690 ( .DIN1(n33388), .DIN2(n33389), .Q(n9554) );
  and2s1 U25691 ( .DIN1(n33329), .DIN2(n33390), .Q(n33389) );
  and2s1 U25692 ( .DIN1(n33024), .DIN2(n32682), .Q(n33388) );
  or2s1 U25693 ( .DIN1(n33391), .DIN2(n33392), .Q(n9553) );
  and2s1 U25694 ( .DIN1(n33329), .DIN2(n33393), .Q(n33392) );
  and2s1 U25695 ( .DIN1(n33024), .DIN2(n32679), .Q(n33391) );
  or2s1 U25696 ( .DIN1(n33394), .DIN2(n33395), .Q(n9552) );
  and2s1 U25697 ( .DIN1(n33329), .DIN2(n33396), .Q(n33395) );
  and2s1 U25698 ( .DIN1(n33024), .DIN2(n32676), .Q(n33394) );
  or2s1 U25699 ( .DIN1(n33397), .DIN2(n33398), .Q(n9551) );
  and2s1 U25700 ( .DIN1(n33329), .DIN2(n33399), .Q(n33398) );
  and2s1 U25701 ( .DIN1(n33024), .DIN2(n32673), .Q(n33397) );
  or2s1 U25702 ( .DIN1(n33400), .DIN2(n33401), .Q(n9550) );
  and2s1 U25703 ( .DIN1(n33329), .DIN2(n33402), .Q(n33401) );
  and2s1 U25704 ( .DIN1(n33024), .DIN2(n32670), .Q(n33400) );
  or2s1 U25705 ( .DIN1(n33403), .DIN2(n33404), .Q(n9549) );
  and2s1 U25706 ( .DIN1(n33329), .DIN2(n33405), .Q(n33404) );
  and2s1 U25707 ( .DIN1(n33024), .DIN2(n32667), .Q(n33403) );
  or2s1 U25708 ( .DIN1(n33406), .DIN2(n33407), .Q(n9548) );
  and2s1 U25709 ( .DIN1(n33329), .DIN2(n33408), .Q(n33407) );
  and2s1 U25710 ( .DIN1(n33024), .DIN2(n32664), .Q(n33406) );
  or2s1 U25711 ( .DIN1(n33409), .DIN2(n33410), .Q(n9547) );
  and2s1 U25712 ( .DIN1(n33329), .DIN2(n33411), .Q(n33410) );
  and2s1 U25713 ( .DIN1(n33024), .DIN2(n32661), .Q(n33409) );
  or2s1 U25714 ( .DIN1(n33412), .DIN2(n33413), .Q(n9546) );
  and2s1 U25715 ( .DIN1(n33329), .DIN2(n33414), .Q(n33413) );
  and2s1 U25716 ( .DIN1(n33024), .DIN2(n32658), .Q(n33412) );
  or2s1 U25717 ( .DIN1(n33415), .DIN2(n33416), .Q(n9545) );
  and2s1 U25718 ( .DIN1(n33329), .DIN2(n33417), .Q(n33416) );
  and2s1 U25719 ( .DIN1(n33024), .DIN2(n32655), .Q(n33415) );
  or2s1 U25720 ( .DIN1(n33418), .DIN2(n33419), .Q(n9544) );
  and2s1 U25721 ( .DIN1(n33329), .DIN2(n33420), .Q(n33419) );
  and2s1 U25722 ( .DIN1(n33024), .DIN2(n32652), .Q(n33418) );
  or2s1 U25723 ( .DIN1(n33421), .DIN2(n33422), .Q(n9543) );
  and2s1 U25724 ( .DIN1(n33329), .DIN2(n33423), .Q(n33422) );
  hi1s1 U25725 ( .DIN1(n33024), .Q(n33329) );
  and2s1 U25726 ( .DIN1(n33024), .DIN2(n32649), .Q(n33421) );
  and2s1 U25727 ( .DIN1(u5_dv), .DIN2(n33022), .Q(n33024) );
  hi1s1 U25728 ( .DIN1(n15477), .Q(n33022) );
  and2s1 U25729 ( .DIN1(n33424), .DIN2(n33425), .Q(n9542) );
  and2s1 U25730 ( .DIN1(n33426), .DIN2(n33427), .Q(n33424) );
  or2s1 U25731 ( .DIN1(n33428), .DIN2(n33429), .Q(n33427) );
  or2s1 U25732 ( .DIN1(u5_ack_cnt[0]), .DIN2(n33430), .Q(n33426) );
  and2s1 U25733 ( .DIN1(n33431), .DIN2(n33425), .Q(n9541) );
  or2s1 U25734 ( .DIN1(n33432), .DIN2(n33433), .Q(n33431) );
  hi1s1 U25735 ( .DIN1(n33434), .Q(n33433) );
  or2s1 U25736 ( .DIN1(n33435), .DIN2(u5_ack_cnt[3]), .Q(n33434) );
  and2s1 U25737 ( .DIN1(u5_ack_cnt[3]), .DIN2(n33435), .Q(n33432) );
  or2s1 U25738 ( .DIN1(n33436), .DIN2(n33428), .Q(n33435) );
  and2s1 U25739 ( .DIN1(n33437), .DIN2(n33438), .Q(n33436) );
  or2s1 U25740 ( .DIN1(n33439), .DIN2(n33440), .Q(n33438) );
  hi1s1 U25741 ( .DIN1(u5_ack_cnt[2]), .Q(n33439) );
  or2s1 U25742 ( .DIN1(n33441), .DIN2(n33442), .Q(n33437) );
  or2s1 U25743 ( .DIN1(u5_ack_cnt[2]), .DIN2(n33443), .Q(n33442) );
  and2s1 U25744 ( .DIN1(n33444), .DIN2(n33425), .Q(n9540) );
  or2s1 U25745 ( .DIN1(n33445), .DIN2(n33446), .Q(n33444) );
  and2s1 U25746 ( .DIN1(u5_ack_cnt[1]), .DIN2(n33428), .Q(n33446) );
  and2s1 U25747 ( .DIN1(n33447), .DIN2(n33448), .Q(n33445) );
  or2s1 U25748 ( .DIN1(n33449), .DIN2(n33450), .Q(n33448) );
  or2s1 U25749 ( .DIN1(n33451), .DIN2(n33452), .Q(n33450) );
  hi1s1 U25750 ( .DIN1(n33453), .Q(n33452) );
  or2s1 U25751 ( .DIN1(n33429), .DIN2(u5_ack_cnt[1]), .Q(n33453) );
  and2s1 U25752 ( .DIN1(u5_ack_cnt[1]), .DIN2(n33429), .Q(n33451) );
  hi1s1 U25753 ( .DIN1(u5_ack_cnt[0]), .Q(n33429) );
  or2s1 U25754 ( .DIN1(n33454), .DIN2(n33455), .Q(n33447) );
  and2s1 U25755 ( .DIN1(n33456), .DIN2(n33430), .Q(n33454) );
  hi1s1 U25756 ( .DIN1(n33428), .Q(n33430) );
  hi1s1 U25757 ( .DIN1(n33457), .Q(n33456) );
  and2s1 U25758 ( .DIN1(n33458), .DIN2(n33425), .Q(n9539) );
  hi1s1 U25759 ( .DIN1(n36596), .Q(n33425) );
  or2s1 U25760 ( .DIN1(n33459), .DIN2(n33460), .Q(n33458) );
  hi1s1 U25761 ( .DIN1(n33461), .Q(n33460) );
  or2s1 U25762 ( .DIN1(n33462), .DIN2(u5_ack_cnt[2]), .Q(n33461) );
  and2s1 U25763 ( .DIN1(u5_ack_cnt[2]), .DIN2(n33462), .Q(n33459) );
  or2s1 U25764 ( .DIN1(n33428), .DIN2(n33463), .Q(n33462) );
  and2s1 U25765 ( .DIN1(n33464), .DIN2(n33440), .Q(n33463) );
  or2s1 U25766 ( .DIN1(n33465), .DIN2(n33449), .Q(n33440) );
  hi1s1 U25767 ( .DIN1(n33441), .Q(n33465) );
  or2s1 U25768 ( .DIN1(n33443), .DIN2(n33441), .Q(n33464) );
  or2s1 U25769 ( .DIN1(n33457), .DIN2(n33455), .Q(n33441) );
  and2s1 U25770 ( .DIN1(u5_ack_cnt[1]), .DIN2(u5_ack_cnt[0]), .Q(n33455) );
  and2s1 U25771 ( .DIN1(n33466), .DIN2(n33449), .Q(n33457) );
  and2s1 U25772 ( .DIN1(n33449), .DIN2(n33467), .Q(n33428) );
  or2s1 U25773 ( .DIN1(n33468), .DIN2(u5_dv), .Q(n33467) );
  hi1s1 U25774 ( .DIN1(n33443), .Q(n33449) );
  and2s1 U25775 ( .DIN1(u5_dv), .DIN2(n33468), .Q(n33443) );
  or2s1 U25776 ( .DIN1(n33469), .DIN2(n33470), .Q(n33468) );
  or2s1 U25777 ( .DIN1(n33471), .DIN2(n33472), .Q(n33470) );
  or2s1 U25778 ( .DIN1(n32961), .DIN2(n32621), .Q(n33472) );
  hi1s1 U25779 ( .DIN1(n33473), .Q(n32961) );
  hi1s1 U25780 ( .DIN1(n15475), .Q(n33471) );
  or2s1 U25781 ( .DIN1(n36597), .DIN2(n33474), .Q(n33469) );
  or2s1 U25782 ( .DIN1(wb_we_i), .DIN2(u5_mem_ack_r), .Q(n33474) );
  or2s1 U25783 ( .DIN1(n33475), .DIN2(n33476), .Q(n9538) );
  or2s1 U25784 ( .DIN1(n33477), .DIN2(n33478), .Q(n33476) );
  and2s1 U25785 ( .DIN1(n33479), .DIN2(n33480), .Q(n33478) );
  and2s1 U25786 ( .DIN1(u5_burst_cnt[10]), .DIN2(n33481), .Q(n33477) );
  or2s1 U25787 ( .DIN1(n33482), .DIN2(n33483), .Q(n33481) );
  and2s1 U25788 ( .DIN1(u5_burst_cnt[9]), .DIN2(n33479), .Q(n33482) );
  and2s1 U25789 ( .DIN1(n32870), .DIN2(n9017), .Q(n33475) );
  or2s1 U25790 ( .DIN1(n33484), .DIN2(n33485), .Q(n9536) );
  and2s1 U25791 ( .DIN1(n32869), .DIN2(n32957), .Q(n33485) );
  and2s1 U25792 ( .DIN1(u5_state[12]), .DIN2(n32844), .Q(n33484) );
  or2s1 U25793 ( .DIN1(n33486), .DIN2(n33487), .Q(n9535) );
  and2s1 U25794 ( .DIN1(u5_state[50]), .DIN2(n32844), .Q(n33486) );
  or2s1 U25795 ( .DIN1(n33488), .DIN2(n33489), .Q(n9534) );
  and2s1 U25796 ( .DIN1(u5_state[17]), .DIN2(n32925), .Q(n33489) );
  and2s1 U25797 ( .DIN1(u5_tmr_done), .DIN2(n33490), .Q(n33488) );
  or2s1 U25798 ( .DIN1(n33491), .DIN2(n33492), .Q(n33490) );
  or2s1 U25799 ( .DIN1(n33493), .DIN2(n33494), .Q(n9531) );
  and2s1 U25800 ( .DIN1(u0_cs[0]), .DIN2(n33495), .Q(n33494) );
  and2s1 U25801 ( .DIN1(u5_cs_le), .DIN2(n33496), .Q(n33493) );
  or2s1 U25802 ( .DIN1(n33497), .DIN2(n33498), .Q(n9530) );
  and2s1 U25803 ( .DIN1(u0_cs[1]), .DIN2(n33495), .Q(n33498) );
  and2s1 U25804 ( .DIN1(n33499), .DIN2(n33500), .Q(n33497) );
  and2s1 U25805 ( .DIN1(u5_cs_le), .DIN2(n33501), .Q(n33499) );
  hi1s1 U25806 ( .DIN1(n33502), .Q(n9529) );
  or2s1 U25807 ( .DIN1(n15500), .DIN2(u5_cs_le), .Q(n33502) );
  hi1s1 U25808 ( .DIN1(n33503), .Q(n9528) );
  or2s1 U25809 ( .DIN1(n15499), .DIN2(u5_cs_le), .Q(n33503) );
  hi1s1 U25810 ( .DIN1(n33504), .Q(n9527) );
  or2s1 U25811 ( .DIN1(n15498), .DIN2(u5_cs_le), .Q(n33504) );
  hi1s1 U25812 ( .DIN1(n33505), .Q(n9526) );
  or2s1 U25813 ( .DIN1(n15497), .DIN2(u5_cs_le), .Q(n33505) );
  hi1s1 U25814 ( .DIN1(n33506), .Q(n9525) );
  or2s1 U25815 ( .DIN1(n15496), .DIN2(u5_cs_le), .Q(n33506) );
  hi1s1 U25816 ( .DIN1(n33507), .Q(n9524) );
  or2s1 U25817 ( .DIN1(n15495), .DIN2(u5_cs_le), .Q(n33507) );
  and2s1 U25818 ( .DIN1(n32625), .DIN2(n4629), .Q(n9522) );
  or2s1 U25819 ( .DIN1(n33508), .DIN2(n33509), .Q(n9521) );
  and2s1 U25820 ( .DIN1(n33510), .DIN2(wb_cyc_i), .Q(n33509) );
  and2s1 U25821 ( .DIN1(n33511), .DIN2(n33512), .Q(n33510) );
  or2s1 U25822 ( .DIN1(n32540), .DIN2(n33495), .Q(n33511) );
  and2s1 U25823 ( .DIN1(n33513), .DIN2(n9523), .Q(n33508) );
  and2s1 U25824 ( .DIN1(n32625), .DIN2(u5_cs_le), .Q(n9523) );
  and2s1 U25825 ( .DIN1(wb_we_i), .DIN2(n33514), .Q(n33513) );
  or2s1 U25826 ( .DIN1(n33515), .DIN2(n33516), .Q(n33514) );
  and2s1 U25827 ( .DIN1(n33517), .DIN2(u0_csc0[8]), .Q(n33516) );
  and2s1 U25828 ( .DIN1(n33500), .DIN2(u0_csc1[8]), .Q(n33515) );
  or2s1 U25829 ( .DIN1(n33518), .DIN2(n33519), .Q(n9520) );
  or2s1 U25830 ( .DIN1(n33520), .DIN2(n33521), .Q(n33519) );
  and2s1 U25831 ( .DIN1(n33522), .DIN2(n32234), .Q(n33521) );
  and2s1 U25832 ( .DIN1(n33523), .DIN2(n32447), .Q(n33520) );
  and2s1 U25833 ( .DIN1(u0_tms[27]), .DIN2(n33524), .Q(n33518) );
  or2s1 U25834 ( .DIN1(n33525), .DIN2(n33526), .Q(n9519) );
  or2s1 U25835 ( .DIN1(n33527), .DIN2(n33528), .Q(n33526) );
  and2s1 U25836 ( .DIN1(n33522), .DIN2(n32238), .Q(n33528) );
  and2s1 U25837 ( .DIN1(n33523), .DIN2(n32450), .Q(n33527) );
  and2s1 U25838 ( .DIN1(u0_tms[26]), .DIN2(n33524), .Q(n33525) );
  or2s1 U25839 ( .DIN1(n33529), .DIN2(n33530), .Q(n9518) );
  or2s1 U25840 ( .DIN1(n33531), .DIN2(n33532), .Q(n33530) );
  and2s1 U25841 ( .DIN1(n33522), .DIN2(n32242), .Q(n33532) );
  and2s1 U25842 ( .DIN1(n33523), .DIN2(n32453), .Q(n33531) );
  and2s1 U25843 ( .DIN1(n33524), .DIN2(u0_tms[25]), .Q(n33529) );
  or2s1 U25844 ( .DIN1(n33533), .DIN2(n33534), .Q(n9517) );
  or2s1 U25845 ( .DIN1(n33535), .DIN2(n33536), .Q(n33534) );
  and2s1 U25846 ( .DIN1(n33522), .DIN2(n32246), .Q(n33536) );
  and2s1 U25847 ( .DIN1(n33523), .DIN2(n32456), .Q(n33535) );
  and2s1 U25848 ( .DIN1(u0_tms[24]), .DIN2(n33524), .Q(n33533) );
  or2s1 U25849 ( .DIN1(n33537), .DIN2(n33538), .Q(n9516) );
  or2s1 U25850 ( .DIN1(n33539), .DIN2(n33540), .Q(n33538) );
  and2s1 U25851 ( .DIN1(n33522), .DIN2(n32250), .Q(n33540) );
  and2s1 U25852 ( .DIN1(n33523), .DIN2(n32459), .Q(n33539) );
  and2s1 U25853 ( .DIN1(u0_tms[23]), .DIN2(n33524), .Q(n33537) );
  or2s1 U25854 ( .DIN1(n33541), .DIN2(n33542), .Q(n9515) );
  or2s1 U25855 ( .DIN1(n33543), .DIN2(n33544), .Q(n33542) );
  and2s1 U25856 ( .DIN1(n33522), .DIN2(n32254), .Q(n33544) );
  and2s1 U25857 ( .DIN1(n33523), .DIN2(n32462), .Q(n33543) );
  and2s1 U25858 ( .DIN1(u0_tms[22]), .DIN2(n33524), .Q(n33541) );
  or2s1 U25859 ( .DIN1(n33545), .DIN2(n33546), .Q(n9514) );
  or2s1 U25860 ( .DIN1(n33547), .DIN2(n33548), .Q(n33546) );
  and2s1 U25861 ( .DIN1(n33522), .DIN2(n32258), .Q(n33548) );
  and2s1 U25862 ( .DIN1(n33523), .DIN2(n32465), .Q(n33547) );
  and2s1 U25863 ( .DIN1(n33524), .DIN2(u0_tms[21]), .Q(n33545) );
  or2s1 U25864 ( .DIN1(n33549), .DIN2(n33550), .Q(n9513) );
  or2s1 U25865 ( .DIN1(n33551), .DIN2(n33552), .Q(n33550) );
  and2s1 U25866 ( .DIN1(n33522), .DIN2(n32262), .Q(n33552) );
  and2s1 U25867 ( .DIN1(n33523), .DIN2(n32468), .Q(n33551) );
  and2s1 U25868 ( .DIN1(n33524), .DIN2(u0_tms[20]), .Q(n33549) );
  or2s1 U25869 ( .DIN1(n33553), .DIN2(n33554), .Q(n9512) );
  or2s1 U25870 ( .DIN1(n33555), .DIN2(n33556), .Q(n33554) );
  and2s1 U25871 ( .DIN1(n33522), .DIN2(n32266), .Q(n33556) );
  and2s1 U25872 ( .DIN1(n33523), .DIN2(n32471), .Q(n33555) );
  and2s1 U25873 ( .DIN1(n33524), .DIN2(u0_tms[19]), .Q(n33553) );
  or2s1 U25874 ( .DIN1(n33557), .DIN2(n33558), .Q(n9511) );
  or2s1 U25875 ( .DIN1(n33559), .DIN2(n33560), .Q(n33558) );
  and2s1 U25876 ( .DIN1(n33522), .DIN2(n32270), .Q(n33560) );
  and2s1 U25877 ( .DIN1(n33523), .DIN2(n32474), .Q(n33559) );
  and2s1 U25878 ( .DIN1(n33524), .DIN2(u0_tms[18]), .Q(n33557) );
  or2s1 U25879 ( .DIN1(n33561), .DIN2(n33562), .Q(n9510) );
  or2s1 U25880 ( .DIN1(n33563), .DIN2(n33564), .Q(n33562) );
  and2s1 U25881 ( .DIN1(n33522), .DIN2(n32274), .Q(n33564) );
  and2s1 U25882 ( .DIN1(n33523), .DIN2(n32477), .Q(n33563) );
  and2s1 U25883 ( .DIN1(n33524), .DIN2(u0_tms[17]), .Q(n33561) );
  or2s1 U25884 ( .DIN1(n33565), .DIN2(n33566), .Q(n9509) );
  or2s1 U25885 ( .DIN1(n33567), .DIN2(n33568), .Q(n33566) );
  and2s1 U25886 ( .DIN1(n33522), .DIN2(n32278), .Q(n33568) );
  and2s1 U25887 ( .DIN1(n33523), .DIN2(n32480), .Q(n33567) );
  and2s1 U25888 ( .DIN1(n33524), .DIN2(u0_tms[16]), .Q(n33565) );
  or2s1 U25889 ( .DIN1(n33569), .DIN2(n33570), .Q(n9508) );
  or2s1 U25890 ( .DIN1(n33571), .DIN2(n33572), .Q(n33570) );
  and2s1 U25891 ( .DIN1(n33522), .DIN2(n32282), .Q(n33572) );
  and2s1 U25892 ( .DIN1(n33523), .DIN2(n32483), .Q(n33571) );
  and2s1 U25893 ( .DIN1(n33524), .DIN2(u0_tms[15]), .Q(n33569) );
  or2s1 U25894 ( .DIN1(n33573), .DIN2(n33574), .Q(n9507) );
  or2s1 U25895 ( .DIN1(n33575), .DIN2(n33576), .Q(n33574) );
  and2s1 U25896 ( .DIN1(n33522), .DIN2(n32286), .Q(n33576) );
  and2s1 U25897 ( .DIN1(n33523), .DIN2(n32486), .Q(n33575) );
  and2s1 U25898 ( .DIN1(u0_tms[14]), .DIN2(n33524), .Q(n33573) );
  or2s1 U25899 ( .DIN1(n33577), .DIN2(n33578), .Q(n9506) );
  or2s1 U25900 ( .DIN1(n33579), .DIN2(n33580), .Q(n33578) );
  and2s1 U25901 ( .DIN1(n33522), .DIN2(n32290), .Q(n33580) );
  and2s1 U25902 ( .DIN1(n33523), .DIN2(n32489), .Q(n33579) );
  and2s1 U25903 ( .DIN1(n33524), .DIN2(u0_tms[13]), .Q(n33577) );
  or2s1 U25904 ( .DIN1(n33581), .DIN2(n33582), .Q(n9505) );
  or2s1 U25905 ( .DIN1(n33583), .DIN2(n33584), .Q(n33582) );
  and2s1 U25906 ( .DIN1(n33522), .DIN2(n32294), .Q(n33584) );
  and2s1 U25907 ( .DIN1(n33523), .DIN2(n32492), .Q(n33583) );
  and2s1 U25908 ( .DIN1(u0_tms[12]), .DIN2(n33524), .Q(n33581) );
  or2s1 U25909 ( .DIN1(n33585), .DIN2(n33586), .Q(n9504) );
  or2s1 U25910 ( .DIN1(n33587), .DIN2(n33588), .Q(n33586) );
  and2s1 U25911 ( .DIN1(n33522), .DIN2(n32298), .Q(n33588) );
  and2s1 U25912 ( .DIN1(n33523), .DIN2(n32495), .Q(n33587) );
  and2s1 U25913 ( .DIN1(u0_tms[11]), .DIN2(n33524), .Q(n33585) );
  or2s1 U25914 ( .DIN1(n33589), .DIN2(n33590), .Q(n9503) );
  or2s1 U25915 ( .DIN1(n33591), .DIN2(n33592), .Q(n33590) );
  and2s1 U25916 ( .DIN1(n33522), .DIN2(n32302), .Q(n33592) );
  and2s1 U25917 ( .DIN1(n33523), .DIN2(n32498), .Q(n33591) );
  and2s1 U25918 ( .DIN1(u0_tms[10]), .DIN2(n33524), .Q(n33589) );
  or2s1 U25919 ( .DIN1(n33593), .DIN2(n33594), .Q(n9502) );
  or2s1 U25920 ( .DIN1(n33595), .DIN2(n33596), .Q(n33594) );
  and2s1 U25921 ( .DIN1(n33522), .DIN2(n32306), .Q(n33596) );
  and2s1 U25922 ( .DIN1(n33523), .DIN2(n32501), .Q(n33595) );
  and2s1 U25923 ( .DIN1(n33524), .DIN2(u0_tms[9]), .Q(n33593) );
  or2s1 U25924 ( .DIN1(n33597), .DIN2(n33598), .Q(n9501) );
  or2s1 U25925 ( .DIN1(n33599), .DIN2(n33600), .Q(n33598) );
  and2s1 U25926 ( .DIN1(n33522), .DIN2(n32310), .Q(n33600) );
  and2s1 U25927 ( .DIN1(n33523), .DIN2(n32504), .Q(n33599) );
  and2s1 U25928 ( .DIN1(u0_tms[8]), .DIN2(n33524), .Q(n33597) );
  or2s1 U25929 ( .DIN1(n33601), .DIN2(n33602), .Q(n9500) );
  or2s1 U25930 ( .DIN1(n33603), .DIN2(n33604), .Q(n33602) );
  and2s1 U25931 ( .DIN1(n33522), .DIN2(n32314), .Q(n33604) );
  and2s1 U25932 ( .DIN1(n33523), .DIN2(n32507), .Q(n33603) );
  and2s1 U25933 ( .DIN1(u0_tms[7]), .DIN2(n33524), .Q(n33601) );
  or2s1 U25934 ( .DIN1(n33605), .DIN2(n33606), .Q(n9499) );
  or2s1 U25935 ( .DIN1(n33607), .DIN2(n33608), .Q(n33606) );
  and2s1 U25936 ( .DIN1(n33522), .DIN2(n32318), .Q(n33608) );
  and2s1 U25937 ( .DIN1(n33523), .DIN2(n32510), .Q(n33607) );
  and2s1 U25938 ( .DIN1(u0_tms[6]), .DIN2(n33524), .Q(n33605) );
  or2s1 U25939 ( .DIN1(n33609), .DIN2(n33610), .Q(n9498) );
  or2s1 U25940 ( .DIN1(n33611), .DIN2(n33612), .Q(n33610) );
  and2s1 U25941 ( .DIN1(n33522), .DIN2(n32322), .Q(n33612) );
  and2s1 U25942 ( .DIN1(n33523), .DIN2(n32513), .Q(n33611) );
  and2s1 U25943 ( .DIN1(n33524), .DIN2(u0_tms[5]), .Q(n33609) );
  or2s1 U25944 ( .DIN1(n33613), .DIN2(n33614), .Q(n9497) );
  or2s1 U25945 ( .DIN1(n33615), .DIN2(n33616), .Q(n33614) );
  and2s1 U25946 ( .DIN1(n33522), .DIN2(n32326), .Q(n33616) );
  and2s1 U25947 ( .DIN1(n33523), .DIN2(n32516), .Q(n33615) );
  and2s1 U25948 ( .DIN1(u0_tms[4]), .DIN2(n33524), .Q(n33613) );
  or2s1 U25949 ( .DIN1(n33617), .DIN2(n33618), .Q(n9496) );
  or2s1 U25950 ( .DIN1(n33619), .DIN2(n33620), .Q(n33618) );
  and2s1 U25951 ( .DIN1(n33522), .DIN2(n32330), .Q(n33620) );
  and2s1 U25952 ( .DIN1(n33523), .DIN2(n32519), .Q(n33619) );
  and2s1 U25953 ( .DIN1(u0_tms[3]), .DIN2(n33524), .Q(n33617) );
  or2s1 U25954 ( .DIN1(n33621), .DIN2(n33622), .Q(n9495) );
  or2s1 U25955 ( .DIN1(n33623), .DIN2(n33624), .Q(n33622) );
  and2s1 U25956 ( .DIN1(n33522), .DIN2(n32334), .Q(n33624) );
  and2s1 U25957 ( .DIN1(n33523), .DIN2(n32522), .Q(n33623) );
  and2s1 U25958 ( .DIN1(n33524), .DIN2(u0_tms[2]), .Q(n33621) );
  or2s1 U25959 ( .DIN1(n33625), .DIN2(n33626), .Q(n9494) );
  or2s1 U25960 ( .DIN1(n33627), .DIN2(n33628), .Q(n33626) );
  and2s1 U25961 ( .DIN1(n33522), .DIN2(n32338), .Q(n33628) );
  and2s1 U25962 ( .DIN1(n33523), .DIN2(n32525), .Q(n33627) );
  and2s1 U25963 ( .DIN1(n33524), .DIN2(u0_tms[1]), .Q(n33625) );
  or2s1 U25964 ( .DIN1(n33629), .DIN2(n33630), .Q(n9493) );
  or2s1 U25965 ( .DIN1(n33631), .DIN2(n33632), .Q(n33630) );
  and2s1 U25966 ( .DIN1(n33522), .DIN2(n32342), .Q(n33632) );
  and2s1 U25967 ( .DIN1(n33633), .DIN2(n33496), .Q(n33522) );
  and2s1 U25968 ( .DIN1(n33523), .DIN2(n32528), .Q(n33631) );
  and2s1 U25969 ( .DIN1(n33633), .DIN2(n33634), .Q(n33523) );
  and2s1 U25970 ( .DIN1(n33524), .DIN2(u0_tms[0]), .Q(n33629) );
  or2s1 U25971 ( .DIN1(n33635), .DIN2(n33636), .Q(n9492) );
  or2s1 U25972 ( .DIN1(n33637), .DIN2(n33638), .Q(n33636) );
  and2s1 U25973 ( .DIN1(n33639), .DIN2(n32199), .Q(n33638) );
  and2s1 U25974 ( .DIN1(n33640), .DIN2(n32402), .Q(n33637) );
  and2s1 U25975 ( .DIN1(u0_csc_10), .DIN2(n33641), .Q(n33635) );
  or2s1 U25976 ( .DIN1(n33642), .DIN2(n33643), .Q(n9491) );
  or2s1 U25977 ( .DIN1(n33644), .DIN2(n33645), .Q(n33643) );
  and2s1 U25978 ( .DIN1(n33639), .DIN2(n32202), .Q(n33645) );
  and2s1 U25979 ( .DIN1(n33640), .DIN2(n32405), .Q(n33644) );
  and2s1 U25980 ( .DIN1(u0_csc_9), .DIN2(n33641), .Q(n33642) );
  or2s1 U25981 ( .DIN1(n33646), .DIN2(n33647), .Q(n9490) );
  or2s1 U25982 ( .DIN1(n33648), .DIN2(n33649), .Q(n33647) );
  and2s1 U25983 ( .DIN1(n33639), .DIN2(n32207), .Q(n33649) );
  and2s1 U25984 ( .DIN1(n33640), .DIN2(n32410), .Q(n33648) );
  and2s1 U25985 ( .DIN1(u0_csc[7]), .DIN2(n33641), .Q(n33646) );
  or2s1 U25986 ( .DIN1(n33650), .DIN2(n33651), .Q(n9489) );
  or2s1 U25987 ( .DIN1(n33652), .DIN2(n33653), .Q(n33651) );
  and2s1 U25988 ( .DIN1(n33639), .DIN2(n32210), .Q(n33653) );
  and2s1 U25989 ( .DIN1(n33640), .DIN2(n32413), .Q(n33652) );
  and2s1 U25990 ( .DIN1(u0_csc[6]), .DIN2(n33641), .Q(n33650) );
  or2s1 U25991 ( .DIN1(n33654), .DIN2(n33655), .Q(n9488) );
  or2s1 U25992 ( .DIN1(n33656), .DIN2(n33657), .Q(n33655) );
  and2s1 U25993 ( .DIN1(n33639), .DIN2(n32834), .Q(n33657) );
  and2s1 U25994 ( .DIN1(n33640), .DIN2(n32416), .Q(n33656) );
  and2s1 U25995 ( .DIN1(u0_csc[5]), .DIN2(n33641), .Q(n33654) );
  or2s1 U25996 ( .DIN1(n33658), .DIN2(n33659), .Q(n9487) );
  or2s1 U25997 ( .DIN1(n33660), .DIN2(n33661), .Q(n33659) );
  and2s1 U25998 ( .DIN1(n33639), .DIN2(n32842), .Q(n33661) );
  and2s1 U25999 ( .DIN1(n33640), .DIN2(n32419), .Q(n33660) );
  and2s1 U26000 ( .DIN1(u0_csc[4]), .DIN2(n33641), .Q(n33658) );
  or2s1 U26001 ( .DIN1(n33662), .DIN2(n33663), .Q(n9486) );
  or2s1 U26002 ( .DIN1(n33664), .DIN2(n33665), .Q(n33663) );
  and2s1 U26003 ( .DIN1(n33639), .DIN2(u0_csc0[3]), .Q(n33665) );
  and2s1 U26004 ( .DIN1(n33640), .DIN2(u0_csc1[3]), .Q(n33664) );
  and2s1 U26005 ( .DIN1(u0_csc[3]), .DIN2(n33641), .Q(n33662) );
  or2s1 U26006 ( .DIN1(n33666), .DIN2(n33667), .Q(n9485) );
  or2s1 U26007 ( .DIN1(n33668), .DIN2(n33669), .Q(n33667) );
  and2s1 U26008 ( .DIN1(n33639), .DIN2(u0_csc0[2]), .Q(n33669) );
  and2s1 U26009 ( .DIN1(n33640), .DIN2(u0_csc1[2]), .Q(n33668) );
  and2s1 U26010 ( .DIN1(u0_csc[2]), .DIN2(n33641), .Q(n33666) );
  or2s1 U26011 ( .DIN1(n33670), .DIN2(n33671), .Q(n9484) );
  or2s1 U26012 ( .DIN1(n33672), .DIN2(n33673), .Q(n33671) );
  and2s1 U26013 ( .DIN1(n33674), .DIN2(n9091), .Q(n33673) );
  and2s1 U26014 ( .DIN1(n33675), .DIN2(n9028), .Q(n33672) );
  or2s1 U26015 ( .DIN1(n33676), .DIN2(n33677), .Q(n33670) );
  or2s1 U26016 ( .DIN1(n33678), .DIN2(n33679), .Q(n33677) );
  and2s1 U26017 ( .DIN1(n33680), .DIN2(n32721), .Q(n33679) );
  and2s1 U26018 ( .DIN1(n33681), .DIN2(n32697), .Q(n33678) );
  and2s1 U26019 ( .DIN1(n33682), .DIN2(n32649), .Q(n33676) );
  hi1s1 U26020 ( .DIN1(n36598), .Q(n32649) );
  or2s1 U26021 ( .DIN1(n33683), .DIN2(n33684), .Q(n9483) );
  or2s1 U26022 ( .DIN1(n33685), .DIN2(n33686), .Q(n33684) );
  and2s1 U26023 ( .DIN1(n33674), .DIN2(n9090), .Q(n33686) );
  and2s1 U26024 ( .DIN1(n33675), .DIN2(n9029), .Q(n33685) );
  or2s1 U26025 ( .DIN1(n33687), .DIN2(n33688), .Q(n33683) );
  or2s1 U26026 ( .DIN1(n33689), .DIN2(n33690), .Q(n33688) );
  and2s1 U26027 ( .DIN1(n33680), .DIN2(n32724), .Q(n33690) );
  and2s1 U26028 ( .DIN1(n33681), .DIN2(n32700), .Q(n33689) );
  and2s1 U26029 ( .DIN1(n33682), .DIN2(n32652), .Q(n33687) );
  hi1s1 U26030 ( .DIN1(n36599), .Q(n32652) );
  or2s1 U26031 ( .DIN1(n33691), .DIN2(n33692), .Q(n9482) );
  or2s1 U26032 ( .DIN1(n33693), .DIN2(n33694), .Q(n33692) );
  and2s1 U26033 ( .DIN1(n33674), .DIN2(n9089), .Q(n33694) );
  and2s1 U26034 ( .DIN1(n33675), .DIN2(n9030), .Q(n33693) );
  or2s1 U26035 ( .DIN1(n33695), .DIN2(n33696), .Q(n33691) );
  or2s1 U26036 ( .DIN1(n33697), .DIN2(n33698), .Q(n33696) );
  and2s1 U26037 ( .DIN1(n33680), .DIN2(n32727), .Q(n33698) );
  and2s1 U26038 ( .DIN1(n33681), .DIN2(n32703), .Q(n33697) );
  and2s1 U26039 ( .DIN1(n33682), .DIN2(n32655), .Q(n33695) );
  hi1s1 U26040 ( .DIN1(n36600), .Q(n32655) );
  or2s1 U26041 ( .DIN1(n33699), .DIN2(n33700), .Q(n9481) );
  or2s1 U26042 ( .DIN1(n33701), .DIN2(n33702), .Q(n33700) );
  and2s1 U26043 ( .DIN1(n33674), .DIN2(n9088), .Q(n33702) );
  and2s1 U26044 ( .DIN1(n33675), .DIN2(n9031), .Q(n33701) );
  or2s1 U26045 ( .DIN1(n33703), .DIN2(n33704), .Q(n33699) );
  or2s1 U26046 ( .DIN1(n33705), .DIN2(n33706), .Q(n33704) );
  and2s1 U26047 ( .DIN1(n33680), .DIN2(n32730), .Q(n33706) );
  and2s1 U26048 ( .DIN1(n33681), .DIN2(n32706), .Q(n33705) );
  and2s1 U26049 ( .DIN1(n33682), .DIN2(n32658), .Q(n33703) );
  hi1s1 U26050 ( .DIN1(n36601), .Q(n32658) );
  or2s1 U26051 ( .DIN1(n33707), .DIN2(n33708), .Q(n9480) );
  or2s1 U26052 ( .DIN1(n33709), .DIN2(n33710), .Q(n33708) );
  and2s1 U26053 ( .DIN1(n33674), .DIN2(n9087), .Q(n33710) );
  and2s1 U26054 ( .DIN1(n33675), .DIN2(n9032), .Q(n33709) );
  or2s1 U26055 ( .DIN1(n33711), .DIN2(n33712), .Q(n33707) );
  or2s1 U26056 ( .DIN1(n33713), .DIN2(n33714), .Q(n33712) );
  and2s1 U26057 ( .DIN1(n33680), .DIN2(n32733), .Q(n33714) );
  and2s1 U26058 ( .DIN1(n33681), .DIN2(n32709), .Q(n33713) );
  and2s1 U26059 ( .DIN1(n33682), .DIN2(n32661), .Q(n33711) );
  hi1s1 U26060 ( .DIN1(n36602), .Q(n32661) );
  or2s1 U26061 ( .DIN1(n33715), .DIN2(n33716), .Q(n9479) );
  or2s1 U26062 ( .DIN1(n33717), .DIN2(n33718), .Q(n33716) );
  and2s1 U26063 ( .DIN1(n33674), .DIN2(n9086), .Q(n33718) );
  and2s1 U26064 ( .DIN1(n33675), .DIN2(n9033), .Q(n33717) );
  or2s1 U26065 ( .DIN1(n33719), .DIN2(n33720), .Q(n33715) );
  or2s1 U26066 ( .DIN1(n33721), .DIN2(n33722), .Q(n33720) );
  and2s1 U26067 ( .DIN1(n33680), .DIN2(n32740), .Q(n33722) );
  and2s1 U26068 ( .DIN1(n33681), .DIN2(n32712), .Q(n33721) );
  and2s1 U26069 ( .DIN1(n33682), .DIN2(n32664), .Q(n33719) );
  hi1s1 U26070 ( .DIN1(n36603), .Q(n32664) );
  or2s1 U26071 ( .DIN1(n33723), .DIN2(n33724), .Q(n9478) );
  or2s1 U26072 ( .DIN1(n33725), .DIN2(n33726), .Q(n33724) );
  and2s1 U26073 ( .DIN1(n33674), .DIN2(n9085), .Q(n33726) );
  and2s1 U26074 ( .DIN1(n33675), .DIN2(n9034), .Q(n33725) );
  or2s1 U26075 ( .DIN1(n33727), .DIN2(n33728), .Q(n33723) );
  or2s1 U26076 ( .DIN1(n33729), .DIN2(n33730), .Q(n33728) );
  and2s1 U26077 ( .DIN1(n33680), .DIN2(n32829), .Q(n33730) );
  and2s1 U26078 ( .DIN1(n33681), .DIN2(n32715), .Q(n33729) );
  and2s1 U26079 ( .DIN1(n33682), .DIN2(n32667), .Q(n33727) );
  hi1s1 U26080 ( .DIN1(n36604), .Q(n32667) );
  or2s1 U26081 ( .DIN1(n33731), .DIN2(n33732), .Q(n9477) );
  or2s1 U26082 ( .DIN1(n33733), .DIN2(n33734), .Q(n33732) );
  and2s1 U26083 ( .DIN1(n33674), .DIN2(n9084), .Q(n33734) );
  and2s1 U26084 ( .DIN1(n33675), .DIN2(n9035), .Q(n33733) );
  or2s1 U26085 ( .DIN1(n33735), .DIN2(n33736), .Q(n33731) );
  or2s1 U26086 ( .DIN1(n33737), .DIN2(n33738), .Q(n33736) );
  and2s1 U26087 ( .DIN1(n33680), .DIN2(n32837), .Q(n33738) );
  and2s1 U26088 ( .DIN1(n33681), .DIN2(n32718), .Q(n33737) );
  and2s1 U26089 ( .DIN1(n33682), .DIN2(n32670), .Q(n33735) );
  hi1s1 U26090 ( .DIN1(n36605), .Q(n32670) );
  or2s1 U26091 ( .DIN1(n33739), .DIN2(n33740), .Q(n9476) );
  or2s1 U26092 ( .DIN1(n33741), .DIN2(n33742), .Q(n33740) );
  and2s1 U26093 ( .DIN1(n33639), .DIN2(n32750), .Q(n33742) );
  and2s1 U26094 ( .DIN1(n33496), .DIN2(n33743), .Q(n33639) );
  and2s1 U26095 ( .DIN1(n33640), .DIN2(n32426), .Q(n33741) );
  and2s1 U26096 ( .DIN1(n33634), .DIN2(n33743), .Q(n33640) );
  and2s1 U26097 ( .DIN1(n33500), .DIN2(n33744), .Q(n33634) );
  and2s1 U26098 ( .DIN1(n33745), .DIN2(n33501), .Q(n33744) );
  hi1s1 U26099 ( .DIN1(n33746), .Q(n33501) );
  and2s1 U26100 ( .DIN1(wb_we_i), .DIN2(u0_csc1[8]), .Q(n33746) );
  hi1s1 U26101 ( .DIN1(n33496), .Q(n33745) );
  and2s1 U26102 ( .DIN1(n33747), .DIN2(n33517), .Q(n33496) );
  hi1s1 U26103 ( .DIN1(n33748), .Q(n33517) );
  or2s1 U26104 ( .DIN1(n33749), .DIN2(n33750), .Q(n33748) );
  or2s1 U26105 ( .DIN1(n33751), .DIN2(n33752), .Q(n33750) );
  or2s1 U26106 ( .DIN1(n33753), .DIN2(n33754), .Q(n33752) );
  hi1s1 U26107 ( .DIN1(n33755), .Q(n33753) );
  or2s1 U26108 ( .DIN1(n33756), .DIN2(u0_csc0[17]), .Q(n33755) );
  or2s1 U26109 ( .DIN1(n33757), .DIN2(n33758), .Q(n33751) );
  or2s1 U26110 ( .DIN1(n33759), .DIN2(n33760), .Q(n33758) );
  and2s1 U26111 ( .DIN1(u0_csc_mask_r[7]), .DIN2(n33761), .Q(n33760) );
  or2s1 U26112 ( .DIN1(n33762), .DIN2(n33763), .Q(n33761) );
  and2s1 U26113 ( .DIN1(u0_csc0[23]), .DIN2(n33764), .Q(n33763) );
  hi1s1 U26114 ( .DIN1(n33765), .Q(n33762) );
  or2s1 U26115 ( .DIN1(n33764), .DIN2(u0_csc0[23]), .Q(n33765) );
  and2s1 U26116 ( .DIN1(u0_csc_mask_r[6]), .DIN2(n33766), .Q(n33759) );
  or2s1 U26117 ( .DIN1(n33767), .DIN2(n33768), .Q(n33766) );
  and2s1 U26118 ( .DIN1(u0_csc0[22]), .DIN2(n33769), .Q(n33768) );
  hi1s1 U26119 ( .DIN1(n33770), .Q(n33767) );
  or2s1 U26120 ( .DIN1(n33769), .DIN2(u0_csc0[22]), .Q(n33770) );
  hi1s1 U26121 ( .DIN1(n33771), .Q(n33757) );
  or2s1 U26122 ( .DIN1(n33772), .DIN2(u0_csc0[16]), .Q(n33771) );
  or2s1 U26123 ( .DIN1(n33773), .DIN2(n33774), .Q(n33749) );
  or2s1 U26124 ( .DIN1(n33775), .DIN2(n33776), .Q(n33774) );
  or2s1 U26125 ( .DIN1(n33777), .DIN2(n33778), .Q(n33776) );
  and2s1 U26126 ( .DIN1(u0_csc_mask_r[4]), .DIN2(n33779), .Q(n33778) );
  or2s1 U26127 ( .DIN1(n33780), .DIN2(n33781), .Q(n33779) );
  and2s1 U26128 ( .DIN1(u0_csc0[20]), .DIN2(n33782), .Q(n33781) );
  hi1s1 U26129 ( .DIN1(n33783), .Q(n33780) );
  or2s1 U26130 ( .DIN1(n33782), .DIN2(u0_csc0[20]), .Q(n33783) );
  and2s1 U26131 ( .DIN1(u0_csc_mask_r[3]), .DIN2(n33784), .Q(n33777) );
  or2s1 U26132 ( .DIN1(n33785), .DIN2(n33786), .Q(n33784) );
  and2s1 U26133 ( .DIN1(u0_csc0[19]), .DIN2(n33787), .Q(n33786) );
  hi1s1 U26134 ( .DIN1(n33788), .Q(n33785) );
  or2s1 U26135 ( .DIN1(n33787), .DIN2(u0_csc0[19]), .Q(n33788) );
  and2s1 U26136 ( .DIN1(u0_csc_mask_r[5]), .DIN2(n33789), .Q(n33775) );
  or2s1 U26137 ( .DIN1(n33790), .DIN2(n33791), .Q(n33789) );
  and2s1 U26138 ( .DIN1(u0_csc0[21]), .DIN2(n33792), .Q(n33791) );
  hi1s1 U26139 ( .DIN1(n33793), .Q(n33790) );
  or2s1 U26140 ( .DIN1(n33792), .DIN2(u0_csc0[21]), .Q(n33793) );
  or2s1 U26141 ( .DIN1(n33794), .DIN2(n33795), .Q(n33773) );
  or2s1 U26142 ( .DIN1(n33796), .DIN2(n33797), .Q(n33795) );
  and2s1 U26143 ( .DIN1(n33798), .DIN2(u0_csc0[17]), .Q(n33797) );
  and2s1 U26144 ( .DIN1(n33799), .DIN2(u0_csc0[16]), .Q(n33796) );
  and2s1 U26145 ( .DIN1(u0_csc_mask_r[2]), .DIN2(n33800), .Q(n33794) );
  or2s1 U26146 ( .DIN1(n33801), .DIN2(n33802), .Q(n33800) );
  and2s1 U26147 ( .DIN1(u0_csc0[18]), .DIN2(n33803), .Q(n33802) );
  hi1s1 U26148 ( .DIN1(n33804), .Q(n33801) );
  or2s1 U26149 ( .DIN1(n33803), .DIN2(u0_csc0[18]), .Q(n33804) );
  hi1s1 U26150 ( .DIN1(n33805), .Q(n33747) );
  and2s1 U26151 ( .DIN1(u0_csc0[8]), .DIN2(wb_we_i), .Q(n33805) );
  hi1s1 U26152 ( .DIN1(n33806), .Q(n33500) );
  or2s1 U26153 ( .DIN1(n33807), .DIN2(n33808), .Q(n33806) );
  or2s1 U26154 ( .DIN1(n33809), .DIN2(n33810), .Q(n33808) );
  or2s1 U26155 ( .DIN1(n33811), .DIN2(n33812), .Q(n33810) );
  hi1s1 U26156 ( .DIN1(n33813), .Q(n33811) );
  or2s1 U26157 ( .DIN1(n33756), .DIN2(u0_csc1[17]), .Q(n33813) );
  or2s1 U26158 ( .DIN1(n33814), .DIN2(n33815), .Q(n33809) );
  or2s1 U26159 ( .DIN1(n33816), .DIN2(n33817), .Q(n33815) );
  and2s1 U26160 ( .DIN1(u0_csc_mask_r[7]), .DIN2(n33818), .Q(n33817) );
  or2s1 U26161 ( .DIN1(n33819), .DIN2(n33820), .Q(n33818) );
  and2s1 U26162 ( .DIN1(u0_csc1[23]), .DIN2(n33764), .Q(n33820) );
  hi1s1 U26163 ( .DIN1(n33821), .Q(n33819) );
  or2s1 U26164 ( .DIN1(n33764), .DIN2(u0_csc1[23]), .Q(n33821) );
  hi1s1 U26165 ( .DIN1(wb_addr_i[28]), .Q(n33764) );
  and2s1 U26166 ( .DIN1(u0_csc_mask_r[6]), .DIN2(n33822), .Q(n33816) );
  or2s1 U26167 ( .DIN1(n33823), .DIN2(n33824), .Q(n33822) );
  and2s1 U26168 ( .DIN1(u0_csc1[22]), .DIN2(n33769), .Q(n33824) );
  hi1s1 U26169 ( .DIN1(n33825), .Q(n33823) );
  or2s1 U26170 ( .DIN1(n33769), .DIN2(u0_csc1[22]), .Q(n33825) );
  hi1s1 U26171 ( .DIN1(wb_addr_i[27]), .Q(n33769) );
  hi1s1 U26172 ( .DIN1(n33826), .Q(n33814) );
  or2s1 U26173 ( .DIN1(n33772), .DIN2(u0_csc1[16]), .Q(n33826) );
  or2s1 U26174 ( .DIN1(n33827), .DIN2(n33828), .Q(n33807) );
  or2s1 U26175 ( .DIN1(n33829), .DIN2(n33830), .Q(n33828) );
  or2s1 U26176 ( .DIN1(n33831), .DIN2(n33832), .Q(n33830) );
  and2s1 U26177 ( .DIN1(u0_csc_mask_r[4]), .DIN2(n33833), .Q(n33832) );
  or2s1 U26178 ( .DIN1(n33834), .DIN2(n33835), .Q(n33833) );
  and2s1 U26179 ( .DIN1(u0_csc1[20]), .DIN2(n33782), .Q(n33835) );
  hi1s1 U26180 ( .DIN1(n33836), .Q(n33834) );
  or2s1 U26181 ( .DIN1(n33782), .DIN2(u0_csc1[20]), .Q(n33836) );
  hi1s1 U26182 ( .DIN1(wb_addr_i[25]), .Q(n33782) );
  and2s1 U26183 ( .DIN1(u0_csc_mask_r[3]), .DIN2(n33837), .Q(n33831) );
  or2s1 U26184 ( .DIN1(n33838), .DIN2(n33839), .Q(n33837) );
  and2s1 U26185 ( .DIN1(u0_csc1[19]), .DIN2(n33787), .Q(n33839) );
  hi1s1 U26186 ( .DIN1(n33840), .Q(n33838) );
  or2s1 U26187 ( .DIN1(n33787), .DIN2(u0_csc1[19]), .Q(n33840) );
  hi1s1 U26188 ( .DIN1(wb_addr_i[24]), .Q(n33787) );
  and2s1 U26189 ( .DIN1(u0_csc_mask_r[5]), .DIN2(n33841), .Q(n33829) );
  or2s1 U26190 ( .DIN1(n33842), .DIN2(n33843), .Q(n33841) );
  and2s1 U26191 ( .DIN1(u0_csc1[21]), .DIN2(n33792), .Q(n33843) );
  hi1s1 U26192 ( .DIN1(n33844), .Q(n33842) );
  or2s1 U26193 ( .DIN1(n33792), .DIN2(u0_csc1[21]), .Q(n33844) );
  hi1s1 U26194 ( .DIN1(wb_addr_i[26]), .Q(n33792) );
  or2s1 U26195 ( .DIN1(n33845), .DIN2(n33846), .Q(n33827) );
  or2s1 U26196 ( .DIN1(n33847), .DIN2(n33848), .Q(n33846) );
  and2s1 U26197 ( .DIN1(n33798), .DIN2(u0_csc1[17]), .Q(n33848) );
  and2s1 U26198 ( .DIN1(u0_csc_mask_r[1]), .DIN2(n33756), .Q(n33798) );
  hi1s1 U26199 ( .DIN1(n33849), .Q(n33756) );
  and2s1 U26200 ( .DIN1(u0_csc_mask_r[1]), .DIN2(wb_addr_i[22]), .Q(n33849) );
  and2s1 U26201 ( .DIN1(n33799), .DIN2(u0_csc1[16]), .Q(n33847) );
  and2s1 U26202 ( .DIN1(u0_csc_mask_r[0]), .DIN2(n33772), .Q(n33799) );
  hi1s1 U26203 ( .DIN1(n33850), .Q(n33772) );
  and2s1 U26204 ( .DIN1(u0_csc_mask_r[0]), .DIN2(wb_addr_i[21]), .Q(n33850) );
  and2s1 U26205 ( .DIN1(u0_csc_mask_r[2]), .DIN2(n33851), .Q(n33845) );
  or2s1 U26206 ( .DIN1(n33852), .DIN2(n33853), .Q(n33851) );
  and2s1 U26207 ( .DIN1(u0_csc1[18]), .DIN2(n33803), .Q(n33853) );
  hi1s1 U26208 ( .DIN1(n33854), .Q(n33852) );
  or2s1 U26209 ( .DIN1(n33803), .DIN2(u0_csc1[18]), .Q(n33854) );
  hi1s1 U26210 ( .DIN1(wb_addr_i[23]), .Q(n33803) );
  and2s1 U26211 ( .DIN1(u0_csc[1]), .DIN2(n33641), .Q(n33739) );
  or2s1 U26212 ( .DIN1(n33855), .DIN2(n33856), .Q(n9475) );
  or2s1 U26213 ( .DIN1(n33857), .DIN2(n33858), .Q(n33856) );
  and2s1 U26214 ( .DIN1(n33859), .DIN2(n33860), .Q(n33858) );
  and2s1 U26215 ( .DIN1(n33861), .DIN2(n33862), .Q(n33857) );
  and2s1 U26216 ( .DIN1(u5_timer2[8]), .DIN2(n33863), .Q(n33861) );
  and2s1 U26217 ( .DIN1(n33864), .DIN2(n33865), .Q(n33855) );
  and2s1 U26218 ( .DIN1(n33866), .DIN2(n33867), .Q(n9474) );
  hi1s1 U26219 ( .DIN1(n33868), .Q(n33867) );
  or2s1 U26220 ( .DIN1(n33869), .DIN2(n33870), .Q(n9473) );
  and2s1 U26221 ( .DIN1(u5_state[51]), .DIN2(n32855), .Q(n33870) );
  and2s1 U26222 ( .DIN1(n33871), .DIN2(u5_tmr2_done), .Q(n33869) );
  or2s1 U26223 ( .DIN1(n33872), .DIN2(n33873), .Q(n9472) );
  and2s1 U26224 ( .DIN1(u5_state[65]), .DIN2(n32844), .Q(n33873) );
  and2s1 U26225 ( .DIN1(n33874), .DIN2(n15513), .Q(n33872) );
  and2s1 U26226 ( .DIN1(u5_tmr2_done), .DIN2(n33875), .Q(n33874) );
  and2s1 U26227 ( .DIN1(n33876), .DIN2(n32638), .Q(n9471) );
  and2s1 U26228 ( .DIN1(n33877), .DIN2(n33878), .Q(n33876) );
  or2s1 U26229 ( .DIN1(n33879), .DIN2(n33512), .Q(n33877) );
  hi1s1 U26230 ( .DIN1(n36606), .Q(n33512) );
  or2s1 U26231 ( .DIN1(n33880), .DIN2(n33881), .Q(n9470) );
  and2s1 U26232 ( .DIN1(n33882), .DIN2(n33883), .Q(n33880) );
  or2s1 U26233 ( .DIN1(n33884), .DIN2(n33885), .Q(n9469) );
  or2s1 U26234 ( .DIN1(u5_wb_stb_first), .DIN2(n33881), .Q(n33885) );
  and2s1 U26235 ( .DIN1(n15473), .DIN2(n33886), .Q(n33881) );
  and2s1 U26236 ( .DIN1(n32638), .DIN2(n15472), .Q(n33886) );
  and2s1 U26237 ( .DIN1(n32625), .DIN2(n32614), .Q(n32638) );
  and2s1 U26238 ( .DIN1(n33887), .DIN2(n33882), .Q(n33884) );
  and2s1 U26239 ( .DIN1(n32626), .DIN2(n33878), .Q(n33882) );
  hi1s1 U26240 ( .DIN1(wb_err_o), .Q(n33878) );
  hi1s1 U26241 ( .DIN1(wb_ack_o), .Q(n32626) );
  and2s1 U26242 ( .DIN1(wb_stb_i), .DIN2(n33883), .Q(n33887) );
  hi1s1 U26243 ( .DIN1(n36607), .Q(n33883) );
  or2s1 U26244 ( .DIN1(n33888), .DIN2(n33889), .Q(n9468) );
  and2s1 U26245 ( .DIN1(u5_state[3]), .DIN2(n32844), .Q(n33888) );
  or2s1 U26246 ( .DIN1(n33890), .DIN2(n33891), .Q(n9467) );
  or2s1 U26247 ( .DIN1(n33892), .DIN2(n33893), .Q(n33891) );
  and2s1 U26248 ( .DIN1(u5_state[1]), .DIN2(n32965), .Q(n33893) );
  and2s1 U26249 ( .DIN1(n33894), .DIN2(n33895), .Q(n33892) );
  or2s1 U26250 ( .DIN1(n33896), .DIN2(n33897), .Q(n33890) );
  and2s1 U26251 ( .DIN1(u5_tmr_done), .DIN2(n33898), .Q(n33897) );
  or2s1 U26252 ( .DIN1(n33899), .DIN2(n33900), .Q(n33898) );
  and2s1 U26253 ( .DIN1(n33901), .DIN2(n33902), .Q(n33899) );
  or2s1 U26254 ( .DIN1(n33903), .DIN2(n33904), .Q(n9466) );
  or2s1 U26255 ( .DIN1(n33905), .DIN2(n33906), .Q(n33904) );
  and2s1 U26256 ( .DIN1(u5_state[9]), .DIN2(n32965), .Q(n33906) );
  and2s1 U26257 ( .DIN1(n33907), .DIN2(n33908), .Q(n33905) );
  or2s1 U26258 ( .DIN1(n33909), .DIN2(n33910), .Q(n33907) );
  and2s1 U26259 ( .DIN1(n33911), .DIN2(u5_tmr_done), .Q(n33909) );
  and2s1 U26260 ( .DIN1(n32962), .DIN2(n33910), .Q(n33903) );
  or2s1 U26261 ( .DIN1(n33912), .DIN2(n33913), .Q(n9465) );
  and2s1 U26262 ( .DIN1(u5_state[25]), .DIN2(n32965), .Q(n33912) );
  or2s1 U26263 ( .DIN1(n33914), .DIN2(n33915), .Q(n9464) );
  hi1s1 U26264 ( .DIN1(n33916), .Q(n33915) );
  and2s1 U26265 ( .DIN1(n33917), .DIN2(n33918), .Q(n33916) );
  and2s1 U26266 ( .DIN1(n33919), .DIN2(n33920), .Q(n33914) );
  or2s1 U26267 ( .DIN1(n33921), .DIN2(n33922), .Q(n9463) );
  and2s1 U26268 ( .DIN1(u0_spec_req_cs[1]), .DIN2(n15511), .Q(n33922) );
  and2s1 U26269 ( .DIN1(n33923), .DIN2(n33924), .Q(n33921) );
  or2s1 U26270 ( .DIN1(n33925), .DIN2(n33926), .Q(n33923) );
  and2s1 U26271 ( .DIN1(n33927), .DIN2(n15509), .Q(n33926) );
  and2s1 U26272 ( .DIN1(u0_init_req), .DIN2(n33928), .Q(n33927) );
  and2s1 U26273 ( .DIN1(n33929), .DIN2(n15506), .Q(n33925) );
  and2s1 U26274 ( .DIN1(n33930), .DIN2(n33920), .Q(n33929) );
  or2s1 U26275 ( .DIN1(n33931), .DIN2(n33932), .Q(n9462) );
  hi1s1 U26276 ( .DIN1(n15483), .Q(n33932) );
  and2s1 U26277 ( .DIN1(n33933), .DIN2(u0_spec_req_cs[1]), .Q(n33931) );
  or2s1 U26278 ( .DIN1(n33934), .DIN2(n33935), .Q(n9461) );
  and2s1 U26279 ( .DIN1(n33936), .DIN2(n33928), .Q(n33935) );
  or2s1 U26280 ( .DIN1(n33937), .DIN2(n33917), .Q(n33936) );
  and2s1 U26281 ( .DIN1(n33938), .DIN2(n32752), .Q(n33934) );
  hi1s1 U26282 ( .DIN1(n33939), .Q(n32752) );
  and2s1 U26283 ( .DIN1(n15483), .DIN2(n4618), .Q(n33938) );
  or2s1 U26284 ( .DIN1(n33940), .DIN2(n33928), .Q(n9460) );
  hi1s1 U26285 ( .DIN1(n36608), .Q(n33928) );
  or2s1 U26286 ( .DIN1(n33941), .DIN2(n33942), .Q(n9459) );
  and2s1 U26287 ( .DIN1(u0_spec_req_cs[0]), .DIN2(n15511), .Q(n33942) );
  and2s1 U26288 ( .DIN1(n33943), .DIN2(n33924), .Q(n33941) );
  or2s1 U26289 ( .DIN1(n33944), .DIN2(n33945), .Q(n33943) );
  and2s1 U26290 ( .DIN1(u0_init_req), .DIN2(n33940), .Q(n33945) );
  and2s1 U26291 ( .DIN1(n33946), .DIN2(n33920), .Q(n33944) );
  hi1s1 U26292 ( .DIN1(u0_init_req), .Q(n33920) );
  or2s1 U26293 ( .DIN1(n33947), .DIN2(n33948), .Q(n9458) );
  hi1s1 U26294 ( .DIN1(n15510), .Q(n33948) );
  and2s1 U26295 ( .DIN1(u0_spec_req_cs[0]), .DIN2(n33933), .Q(n33947) );
  hi1s1 U26296 ( .DIN1(n33917), .Q(n33933) );
  or2s1 U26297 ( .DIN1(n33949), .DIN2(n33950), .Q(n9457) );
  and2s1 U26298 ( .DIN1(n33951), .DIN2(n33940), .Q(n33950) );
  hi1s1 U26299 ( .DIN1(n15509), .Q(n33940) );
  or2s1 U26300 ( .DIN1(n33917), .DIN2(n33952), .Q(n33951) );
  or2s1 U26301 ( .DIN1(u5_init_ack), .DIN2(n4989), .Q(n33917) );
  and2s1 U26302 ( .DIN1(n33953), .DIN2(n32751), .Q(n33949) );
  hi1s1 U26303 ( .DIN1(n33954), .Q(n32751) );
  and2s1 U26304 ( .DIN1(n15510), .DIN2(n4616), .Q(n33953) );
  or2s1 U26305 ( .DIN1(n33955), .DIN2(n33956), .Q(n9456) );
  or2s1 U26306 ( .DIN1(n33957), .DIN2(n33958), .Q(n33956) );
  and2s1 U26307 ( .DIN1(n33959), .DIN2(n32447), .Q(n33958) );
  and2s1 U26308 ( .DIN1(n33960), .DIN2(n32234), .Q(n33957) );
  and2s1 U26309 ( .DIN1(u0_sp_tms[27]), .DIN2(n33524), .Q(n33955) );
  or2s1 U26310 ( .DIN1(n33961), .DIN2(n33962), .Q(n9455) );
  or2s1 U26311 ( .DIN1(n33963), .DIN2(n33964), .Q(n33962) );
  and2s1 U26312 ( .DIN1(n33959), .DIN2(n32450), .Q(n33964) );
  and2s1 U26313 ( .DIN1(n33960), .DIN2(n32238), .Q(n33963) );
  and2s1 U26314 ( .DIN1(u0_sp_tms[26]), .DIN2(n33524), .Q(n33961) );
  or2s1 U26315 ( .DIN1(n33965), .DIN2(n33966), .Q(n9454) );
  or2s1 U26316 ( .DIN1(n33967), .DIN2(n33968), .Q(n33966) );
  and2s1 U26317 ( .DIN1(n33959), .DIN2(n32453), .Q(n33968) );
  and2s1 U26318 ( .DIN1(n33960), .DIN2(n32242), .Q(n33967) );
  and2s1 U26319 ( .DIN1(n33524), .DIN2(u0_sp_tms[25]), .Q(n33965) );
  or2s1 U26320 ( .DIN1(n33969), .DIN2(n33970), .Q(n9453) );
  or2s1 U26321 ( .DIN1(n33971), .DIN2(n33972), .Q(n33970) );
  and2s1 U26322 ( .DIN1(n33959), .DIN2(n32456), .Q(n33972) );
  and2s1 U26323 ( .DIN1(n33960), .DIN2(n32246), .Q(n33971) );
  and2s1 U26324 ( .DIN1(u0_sp_tms[24]), .DIN2(n33524), .Q(n33969) );
  or2s1 U26325 ( .DIN1(n33973), .DIN2(n33974), .Q(n9452) );
  or2s1 U26326 ( .DIN1(n33975), .DIN2(n33976), .Q(n33974) );
  and2s1 U26327 ( .DIN1(n33959), .DIN2(n32459), .Q(n33976) );
  and2s1 U26328 ( .DIN1(n33960), .DIN2(n32250), .Q(n33975) );
  and2s1 U26329 ( .DIN1(u0_sp_tms[23]), .DIN2(n33524), .Q(n33973) );
  or2s1 U26330 ( .DIN1(n33977), .DIN2(n33978), .Q(n9451) );
  or2s1 U26331 ( .DIN1(n33979), .DIN2(n33980), .Q(n33978) );
  and2s1 U26332 ( .DIN1(n33959), .DIN2(n32462), .Q(n33980) );
  and2s1 U26333 ( .DIN1(n33960), .DIN2(n32254), .Q(n33979) );
  and2s1 U26334 ( .DIN1(u0_sp_tms[22]), .DIN2(n33524), .Q(n33977) );
  or2s1 U26335 ( .DIN1(n33981), .DIN2(n33982), .Q(n9450) );
  or2s1 U26336 ( .DIN1(n33983), .DIN2(n33984), .Q(n33982) );
  and2s1 U26337 ( .DIN1(n33959), .DIN2(n32465), .Q(n33984) );
  and2s1 U26338 ( .DIN1(n33960), .DIN2(n32258), .Q(n33983) );
  and2s1 U26339 ( .DIN1(n33524), .DIN2(u0_sp_tms[21]), .Q(n33981) );
  or2s1 U26340 ( .DIN1(n33985), .DIN2(n33986), .Q(n9449) );
  or2s1 U26341 ( .DIN1(n33987), .DIN2(n33988), .Q(n33986) );
  and2s1 U26342 ( .DIN1(n33959), .DIN2(n32468), .Q(n33988) );
  and2s1 U26343 ( .DIN1(n33960), .DIN2(n32262), .Q(n33987) );
  and2s1 U26344 ( .DIN1(n33524), .DIN2(u0_sp_tms[20]), .Q(n33985) );
  or2s1 U26345 ( .DIN1(n33989), .DIN2(n33990), .Q(n9448) );
  or2s1 U26346 ( .DIN1(n33991), .DIN2(n33992), .Q(n33990) );
  and2s1 U26347 ( .DIN1(n33959), .DIN2(n32471), .Q(n33992) );
  and2s1 U26348 ( .DIN1(n33960), .DIN2(n32266), .Q(n33991) );
  and2s1 U26349 ( .DIN1(n33524), .DIN2(u0_sp_tms[19]), .Q(n33989) );
  or2s1 U26350 ( .DIN1(n33993), .DIN2(n33994), .Q(n9447) );
  or2s1 U26351 ( .DIN1(n33995), .DIN2(n33996), .Q(n33994) );
  and2s1 U26352 ( .DIN1(n33959), .DIN2(n32474), .Q(n33996) );
  and2s1 U26353 ( .DIN1(n33960), .DIN2(n32270), .Q(n33995) );
  and2s1 U26354 ( .DIN1(n33524), .DIN2(u0_sp_tms[18]), .Q(n33993) );
  or2s1 U26355 ( .DIN1(n33997), .DIN2(n33998), .Q(n9446) );
  or2s1 U26356 ( .DIN1(n33999), .DIN2(n34000), .Q(n33998) );
  and2s1 U26357 ( .DIN1(n33959), .DIN2(n32477), .Q(n34000) );
  and2s1 U26358 ( .DIN1(n33960), .DIN2(n32274), .Q(n33999) );
  and2s1 U26359 ( .DIN1(n33524), .DIN2(u0_sp_tms[17]), .Q(n33997) );
  or2s1 U26360 ( .DIN1(n34001), .DIN2(n34002), .Q(n9445) );
  or2s1 U26361 ( .DIN1(n34003), .DIN2(n34004), .Q(n34002) );
  and2s1 U26362 ( .DIN1(n33959), .DIN2(n32480), .Q(n34004) );
  and2s1 U26363 ( .DIN1(n33960), .DIN2(n32278), .Q(n34003) );
  and2s1 U26364 ( .DIN1(n33524), .DIN2(u0_sp_tms[16]), .Q(n34001) );
  or2s1 U26365 ( .DIN1(n34005), .DIN2(n34006), .Q(n9444) );
  or2s1 U26366 ( .DIN1(n34007), .DIN2(n34008), .Q(n34006) );
  and2s1 U26367 ( .DIN1(n33959), .DIN2(n32483), .Q(n34008) );
  and2s1 U26368 ( .DIN1(n33960), .DIN2(n32282), .Q(n34007) );
  and2s1 U26369 ( .DIN1(n33524), .DIN2(u0_sp_tms[15]), .Q(n34005) );
  or2s1 U26370 ( .DIN1(n34009), .DIN2(n34010), .Q(n9443) );
  or2s1 U26371 ( .DIN1(n34011), .DIN2(n34012), .Q(n34010) );
  and2s1 U26372 ( .DIN1(n33959), .DIN2(n32486), .Q(n34012) );
  and2s1 U26373 ( .DIN1(n33960), .DIN2(n32286), .Q(n34011) );
  and2s1 U26374 ( .DIN1(u0_sp_tms[14]), .DIN2(n33524), .Q(n34009) );
  or2s1 U26375 ( .DIN1(n34013), .DIN2(n34014), .Q(n9442) );
  or2s1 U26376 ( .DIN1(n34015), .DIN2(n34016), .Q(n34014) );
  and2s1 U26377 ( .DIN1(n33959), .DIN2(n32489), .Q(n34016) );
  and2s1 U26378 ( .DIN1(n33960), .DIN2(n32290), .Q(n34015) );
  and2s1 U26379 ( .DIN1(n33524), .DIN2(u0_sp_tms[13]), .Q(n34013) );
  or2s1 U26380 ( .DIN1(n34017), .DIN2(n34018), .Q(n9441) );
  or2s1 U26381 ( .DIN1(n34019), .DIN2(n34020), .Q(n34018) );
  and2s1 U26382 ( .DIN1(n33959), .DIN2(n32492), .Q(n34020) );
  and2s1 U26383 ( .DIN1(n33960), .DIN2(n32294), .Q(n34019) );
  and2s1 U26384 ( .DIN1(u0_sp_tms[12]), .DIN2(n33524), .Q(n34017) );
  or2s1 U26385 ( .DIN1(n34021), .DIN2(n34022), .Q(n9440) );
  or2s1 U26386 ( .DIN1(n34023), .DIN2(n34024), .Q(n34022) );
  and2s1 U26387 ( .DIN1(n33959), .DIN2(n32495), .Q(n34024) );
  and2s1 U26388 ( .DIN1(n33960), .DIN2(n32298), .Q(n34023) );
  and2s1 U26389 ( .DIN1(u0_sp_tms[11]), .DIN2(n33524), .Q(n34021) );
  or2s1 U26390 ( .DIN1(n34025), .DIN2(n34026), .Q(n9439) );
  or2s1 U26391 ( .DIN1(n34027), .DIN2(n34028), .Q(n34026) );
  and2s1 U26392 ( .DIN1(n33959), .DIN2(n32498), .Q(n34028) );
  and2s1 U26393 ( .DIN1(n33960), .DIN2(n32302), .Q(n34027) );
  and2s1 U26394 ( .DIN1(u0_sp_tms[10]), .DIN2(n33524), .Q(n34025) );
  or2s1 U26395 ( .DIN1(n34029), .DIN2(n34030), .Q(n9438) );
  or2s1 U26396 ( .DIN1(n34031), .DIN2(n34032), .Q(n34030) );
  and2s1 U26397 ( .DIN1(n33959), .DIN2(n32501), .Q(n34032) );
  and2s1 U26398 ( .DIN1(n33960), .DIN2(n32306), .Q(n34031) );
  and2s1 U26399 ( .DIN1(n33524), .DIN2(u0_sp_tms[9]), .Q(n34029) );
  or2s1 U26400 ( .DIN1(n34033), .DIN2(n34034), .Q(n9437) );
  or2s1 U26401 ( .DIN1(n34035), .DIN2(n34036), .Q(n34034) );
  and2s1 U26402 ( .DIN1(n33959), .DIN2(n32504), .Q(n34036) );
  and2s1 U26403 ( .DIN1(n33960), .DIN2(n32310), .Q(n34035) );
  and2s1 U26404 ( .DIN1(u0_sp_tms[8]), .DIN2(n33524), .Q(n34033) );
  or2s1 U26405 ( .DIN1(n34037), .DIN2(n34038), .Q(n9436) );
  or2s1 U26406 ( .DIN1(n34039), .DIN2(n34040), .Q(n34038) );
  and2s1 U26407 ( .DIN1(n33959), .DIN2(n32507), .Q(n34040) );
  and2s1 U26408 ( .DIN1(n33960), .DIN2(n32314), .Q(n34039) );
  and2s1 U26409 ( .DIN1(u0_sp_tms[7]), .DIN2(n33524), .Q(n34037) );
  or2s1 U26410 ( .DIN1(n34041), .DIN2(n34042), .Q(n9435) );
  or2s1 U26411 ( .DIN1(n34043), .DIN2(n34044), .Q(n34042) );
  and2s1 U26412 ( .DIN1(n33959), .DIN2(n32510), .Q(n34044) );
  and2s1 U26413 ( .DIN1(n33960), .DIN2(n32318), .Q(n34043) );
  and2s1 U26414 ( .DIN1(u0_sp_tms[6]), .DIN2(n33524), .Q(n34041) );
  or2s1 U26415 ( .DIN1(n34045), .DIN2(n34046), .Q(n9434) );
  or2s1 U26416 ( .DIN1(n34047), .DIN2(n34048), .Q(n34046) );
  and2s1 U26417 ( .DIN1(n33959), .DIN2(n32513), .Q(n34048) );
  and2s1 U26418 ( .DIN1(n33960), .DIN2(n32322), .Q(n34047) );
  and2s1 U26419 ( .DIN1(n33524), .DIN2(u0_sp_tms[5]), .Q(n34045) );
  or2s1 U26420 ( .DIN1(n34049), .DIN2(n34050), .Q(n9433) );
  or2s1 U26421 ( .DIN1(n34051), .DIN2(n34052), .Q(n34050) );
  and2s1 U26422 ( .DIN1(n33959), .DIN2(n32516), .Q(n34052) );
  and2s1 U26423 ( .DIN1(n33960), .DIN2(n32326), .Q(n34051) );
  and2s1 U26424 ( .DIN1(u0_sp_tms[4]), .DIN2(n33524), .Q(n34049) );
  or2s1 U26425 ( .DIN1(n34053), .DIN2(n34054), .Q(n9432) );
  or2s1 U26426 ( .DIN1(n34055), .DIN2(n34056), .Q(n34054) );
  and2s1 U26427 ( .DIN1(n33959), .DIN2(n32519), .Q(n34056) );
  and2s1 U26428 ( .DIN1(n33960), .DIN2(n32330), .Q(n34055) );
  and2s1 U26429 ( .DIN1(u0_sp_tms[3]), .DIN2(n33524), .Q(n34053) );
  or2s1 U26430 ( .DIN1(n34057), .DIN2(n34058), .Q(n9431) );
  or2s1 U26431 ( .DIN1(n34059), .DIN2(n34060), .Q(n34058) );
  and2s1 U26432 ( .DIN1(n33959), .DIN2(n32522), .Q(n34060) );
  and2s1 U26433 ( .DIN1(n33960), .DIN2(n32334), .Q(n34059) );
  and2s1 U26434 ( .DIN1(n33524), .DIN2(u0_sp_tms[2]), .Q(n34057) );
  or2s1 U26435 ( .DIN1(n34061), .DIN2(n34062), .Q(n9430) );
  or2s1 U26436 ( .DIN1(n34063), .DIN2(n34064), .Q(n34062) );
  and2s1 U26437 ( .DIN1(n33959), .DIN2(n32525), .Q(n34064) );
  and2s1 U26438 ( .DIN1(n33960), .DIN2(n32338), .Q(n34063) );
  and2s1 U26439 ( .DIN1(n33524), .DIN2(u0_sp_tms[1]), .Q(n34061) );
  or2s1 U26440 ( .DIN1(n34065), .DIN2(n34066), .Q(n9429) );
  or2s1 U26441 ( .DIN1(n34067), .DIN2(n34068), .Q(n34066) );
  and2s1 U26442 ( .DIN1(n33959), .DIN2(n32528), .Q(n34068) );
  and2s1 U26443 ( .DIN1(u0_spec_req_cs[1]), .DIN2(n34069), .Q(n33959) );
  and2s1 U26444 ( .DIN1(n33952), .DIN2(n33633), .Q(n34069) );
  and2s1 U26445 ( .DIN1(n33960), .DIN2(n32342), .Q(n34067) );
  and2s1 U26446 ( .DIN1(n33633), .DIN2(u0_spec_req_cs[0]), .Q(n33960) );
  hi1s1 U26447 ( .DIN1(n33524), .Q(n33633) );
  and2s1 U26448 ( .DIN1(n33524), .DIN2(u0_sp_tms[0]), .Q(n34065) );
  and2s1 U26449 ( .DIN1(n33641), .DIN2(n34070), .Q(n33524) );
  or2s1 U26450 ( .DIN1(n32033), .DIN2(n32621), .Q(n34070) );
  or2s1 U26451 ( .DIN1(n34071), .DIN2(n34072), .Q(n9428) );
  or2s1 U26452 ( .DIN1(n34073), .DIN2(n34074), .Q(n34072) );
  and2s1 U26453 ( .DIN1(n34075), .DIN2(n32402), .Q(n34074) );
  and2s1 U26454 ( .DIN1(n34076), .DIN2(n32199), .Q(n34073) );
  and2s1 U26455 ( .DIN1(u0_sp_csc_10), .DIN2(n33641), .Q(n34071) );
  or2s1 U26456 ( .DIN1(n34077), .DIN2(n34078), .Q(n9427) );
  or2s1 U26457 ( .DIN1(n34079), .DIN2(n34080), .Q(n34078) );
  and2s1 U26458 ( .DIN1(n34075), .DIN2(n32405), .Q(n34080) );
  and2s1 U26459 ( .DIN1(n34076), .DIN2(n32202), .Q(n34079) );
  and2s1 U26460 ( .DIN1(u0_sp_csc_9), .DIN2(n33641), .Q(n34077) );
  or2s1 U26461 ( .DIN1(n34081), .DIN2(n34082), .Q(n9426) );
  or2s1 U26462 ( .DIN1(n34083), .DIN2(n34084), .Q(n34082) );
  and2s1 U26463 ( .DIN1(n34075), .DIN2(n32410), .Q(n34084) );
  and2s1 U26464 ( .DIN1(n34076), .DIN2(n32207), .Q(n34083) );
  and2s1 U26465 ( .DIN1(u0_sp_csc[7]), .DIN2(n33641), .Q(n34081) );
  or2s1 U26466 ( .DIN1(n34085), .DIN2(n34086), .Q(n9425) );
  or2s1 U26467 ( .DIN1(n34087), .DIN2(n34088), .Q(n34086) );
  and2s1 U26468 ( .DIN1(n34075), .DIN2(n32413), .Q(n34088) );
  and2s1 U26469 ( .DIN1(n34076), .DIN2(n32210), .Q(n34087) );
  and2s1 U26470 ( .DIN1(u0_sp_csc[6]), .DIN2(n33641), .Q(n34085) );
  or2s1 U26471 ( .DIN1(n34089), .DIN2(n34090), .Q(n9424) );
  or2s1 U26472 ( .DIN1(n34091), .DIN2(n34092), .Q(n34090) );
  and2s1 U26473 ( .DIN1(n34075), .DIN2(n32416), .Q(n34092) );
  and2s1 U26474 ( .DIN1(n34076), .DIN2(n32834), .Q(n34091) );
  and2s1 U26475 ( .DIN1(n33641), .DIN2(n34093), .Q(n34089) );
  or2s1 U26476 ( .DIN1(n34094), .DIN2(n34095), .Q(n9423) );
  or2s1 U26477 ( .DIN1(n34096), .DIN2(n34097), .Q(n34095) );
  and2s1 U26478 ( .DIN1(n34075), .DIN2(n32419), .Q(n34097) );
  and2s1 U26479 ( .DIN1(n34076), .DIN2(n32842), .Q(n34096) );
  and2s1 U26480 ( .DIN1(u0_sp_csc[4]), .DIN2(n33641), .Q(n34094) );
  or2s1 U26481 ( .DIN1(n34098), .DIN2(n34099), .Q(n9422) );
  and2s1 U26482 ( .DIN1(u5_state[41]), .DIN2(n32844), .Q(n34099) );
  and2s1 U26483 ( .DIN1(n34100), .DIN2(n32849), .Q(n34098) );
  or2s1 U26484 ( .DIN1(n34101), .DIN2(n34102), .Q(n9421) );
  and2s1 U26485 ( .DIN1(u5_state[42]), .DIN2(n32844), .Q(n34101) );
  or2s1 U26486 ( .DIN1(n34103), .DIN2(n34104), .Q(n9420) );
  and2s1 U26487 ( .DIN1(u5_state[43]), .DIN2(n32925), .Q(n34104) );
  and2s1 U26488 ( .DIN1(n34105), .DIN2(n34106), .Q(n34103) );
  and2s1 U26489 ( .DIN1(n34107), .DIN2(u5_tmr2_done), .Q(n34105) );
  or2s1 U26490 ( .DIN1(n34108), .DIN2(n19411), .Q(n9419) );
  and2s1 U26491 ( .DIN1(u5_state[44]), .DIN2(n32844), .Q(n34108) );
  or2s1 U26492 ( .DIN1(n34109), .DIN2(n34110), .Q(n9418) );
  and2s1 U26493 ( .DIN1(n34111), .DIN2(n32921), .Q(n34110) );
  and2s1 U26494 ( .DIN1(u5_state[53]), .DIN2(n32855), .Q(n34109) );
  or2s1 U26495 ( .DIN1(n34112), .DIN2(n34113), .Q(n9417) );
  and2s1 U26496 ( .DIN1(u5_state[54]), .DIN2(n32925), .Q(n34113) );
  and2s1 U26497 ( .DIN1(n34114), .DIN2(u5_tmr2_done), .Q(n34112) );
  or2s1 U26498 ( .DIN1(n34115), .DIN2(n34116), .Q(n9416) );
  and2s1 U26499 ( .DIN1(u5_state[55]), .DIN2(n32844), .Q(n34115) );
  or2s1 U26500 ( .DIN1(n34117), .DIN2(n34118), .Q(n9415) );
  or2s1 U26501 ( .DIN1(n34119), .DIN2(n34120), .Q(n34118) );
  and2s1 U26502 ( .DIN1(n34121), .DIN2(n32921), .Q(n34120) );
  and2s1 U26503 ( .DIN1(u5_state[57]), .DIN2(n32922), .Q(n34119) );
  or2s1 U26504 ( .DIN1(n34122), .DIN2(n34123), .Q(n9414) );
  and2s1 U26505 ( .DIN1(u5_state[6]), .DIN2(n32844), .Q(n34123) );
  and2s1 U26506 ( .DIN1(n34124), .DIN2(u5_tmr_done), .Q(n34122) );
  and2s1 U26507 ( .DIN1(n34125), .DIN2(n34126), .Q(n34124) );
  or2s1 U26508 ( .DIN1(n34127), .DIN2(n34128), .Q(n9413) );
  and2s1 U26509 ( .DIN1(n32896), .DIN2(n34129), .Q(n34128) );
  and2s1 U26510 ( .DIN1(u5_state[64]), .DIN2(n32844), .Q(n34127) );
  or2s1 U26511 ( .DIN1(n34130), .DIN2(n34131), .Q(n9412) );
  hi1s1 U26512 ( .DIN1(n34132), .Q(n34131) );
  and2s1 U26513 ( .DIN1(n34133), .DIN2(u5_ir_cnt[0]), .Q(n34130) );
  or2s1 U26514 ( .DIN1(n34134), .DIN2(n34135), .Q(n9411) );
  or2s1 U26515 ( .DIN1(n34136), .DIN2(n34137), .Q(n34135) );
  and2s1 U26516 ( .DIN1(u5_ir_cnt[1]), .DIN2(n34132), .Q(n34137) );
  or2s1 U26517 ( .DIN1(u5_ir_cnt[0]), .DIN2(n34138), .Q(n34132) );
  or2s1 U26518 ( .DIN1(n34139), .DIN2(n34140), .Q(n9410) );
  and2s1 U26519 ( .DIN1(n34141), .DIN2(n34142), .Q(n34140) );
  and2s1 U26520 ( .DIN1(n34134), .DIN2(n15508), .Q(n34139) );
  and2s1 U26521 ( .DIN1(n34143), .DIN2(n33913), .Q(n34134) );
  or2s1 U26522 ( .DIN1(n34144), .DIN2(n34145), .Q(n9408) );
  and2s1 U26523 ( .DIN1(n19413), .DIN2(n33913), .Q(n34145) );
  and2s1 U26524 ( .DIN1(n34146), .DIN2(n34147), .Q(n34144) );
  hi1s1 U26525 ( .DIN1(n15474), .Q(n34147) );
  or2s1 U26526 ( .DIN1(n34148), .DIN2(n34141), .Q(n34146) );
  or2s1 U26527 ( .DIN1(n34149), .DIN2(n34133), .Q(n34141) );
  and2s1 U26528 ( .DIN1(n34138), .DIN2(n34150), .Q(n34133) );
  hi1s1 U26529 ( .DIN1(n33913), .Q(n34138) );
  and2s1 U26530 ( .DIN1(n33913), .DIN2(n34151), .Q(n34149) );
  and2s1 U26531 ( .DIN1(n33913), .DIN2(n34142), .Q(n34148) );
  hi1s1 U26532 ( .DIN1(n15508), .Q(n34142) );
  and2s1 U26533 ( .DIN1(n32921), .DIN2(n34152), .Q(n33913) );
  or2s1 U26534 ( .DIN1(n34153), .DIN2(n34154), .Q(n9407) );
  and2s1 U26535 ( .DIN1(n34136), .DIN2(n32921), .Q(n34154) );
  and2s1 U26536 ( .DIN1(u5_state[23]), .DIN2(n32965), .Q(n34153) );
  or2s1 U26537 ( .DIN1(n34155), .DIN2(n34156), .Q(n9406) );
  and2s1 U26538 ( .DIN1(u5_state[29]), .DIN2(n32925), .Q(n34156) );
  and2s1 U26539 ( .DIN1(n34157), .DIN2(n34158), .Q(n34155) );
  and2s1 U26540 ( .DIN1(u5_state[28]), .DIN2(u5_tmr_done), .Q(n34157) );
  or2s1 U26541 ( .DIN1(n34159), .DIN2(n34160), .Q(n9405) );
  and2s1 U26542 ( .DIN1(n34161), .DIN2(n32921), .Q(n34160) );
  and2s1 U26543 ( .DIN1(u5_state[30]), .DIN2(n32922), .Q(n34159) );
  or2s1 U26544 ( .DIN1(n34162), .DIN2(n32855), .Q(n32922) );
  or2s1 U26545 ( .DIN1(n34163), .DIN2(n34164), .Q(n9404) );
  and2s1 U26546 ( .DIN1(u4_rfr_cnt[7]), .DIN2(n34165), .Q(n34164) );
  or2s1 U26547 ( .DIN1(n34166), .DIN2(n34167), .Q(n34165) );
  and2s1 U26548 ( .DIN1(n34168), .DIN2(n34169), .Q(n34166) );
  and2s1 U26549 ( .DIN1(n34170), .DIN2(u4_rfr_cnt[6]), .Q(n34163) );
  and2s1 U26550 ( .DIN1(n34171), .DIN2(n34172), .Q(n34170) );
  hi1s1 U26551 ( .DIN1(u4_rfr_cnt[7]), .Q(n34172) );
  or2s1 U26552 ( .DIN1(n34173), .DIN2(n34174), .Q(n9403) );
  and2s1 U26553 ( .DIN1(n34175), .DIN2(u4_rfr_cnt[0]), .Q(n34173) );
  or2s1 U26554 ( .DIN1(n34176), .DIN2(n34177), .Q(n9402) );
  and2s1 U26555 ( .DIN1(u4_rfr_cnt[1]), .DIN2(n34178), .Q(n34177) );
  and2s1 U26556 ( .DIN1(n34179), .DIN2(n34168), .Q(n34176) );
  and2s1 U26557 ( .DIN1(u4_rfr_cnt[0]), .DIN2(n34180), .Q(n34179) );
  or2s1 U26558 ( .DIN1(n34181), .DIN2(n34182), .Q(n9401) );
  and2s1 U26559 ( .DIN1(u4_rfr_cnt[2]), .DIN2(n34183), .Q(n34182) );
  or2s1 U26560 ( .DIN1(n34184), .DIN2(n34178), .Q(n34183) );
  or2s1 U26561 ( .DIN1(n34174), .DIN2(n34175), .Q(n34178) );
  and2s1 U26562 ( .DIN1(n34168), .DIN2(n34185), .Q(n34174) );
  and2s1 U26563 ( .DIN1(n34168), .DIN2(n34180), .Q(n34184) );
  and2s1 U26564 ( .DIN1(n34186), .DIN2(n34187), .Q(n34181) );
  and2s1 U26565 ( .DIN1(u4_rfr_cnt[0]), .DIN2(n34188), .Q(n34187) );
  and2s1 U26566 ( .DIN1(n34168), .DIN2(u4_rfr_cnt[1]), .Q(n34186) );
  or2s1 U26567 ( .DIN1(n34189), .DIN2(n34190), .Q(n9400) );
  and2s1 U26568 ( .DIN1(u4_rfr_cnt[3]), .DIN2(n34191), .Q(n34190) );
  and2s1 U26569 ( .DIN1(n34192), .DIN2(n34168), .Q(n34189) );
  and2s1 U26570 ( .DIN1(n34193), .DIN2(n34194), .Q(n34192) );
  or2s1 U26571 ( .DIN1(n34195), .DIN2(n34196), .Q(n9399) );
  and2s1 U26572 ( .DIN1(u4_rfr_cnt[4]), .DIN2(n34197), .Q(n34196) );
  or2s1 U26573 ( .DIN1(n34198), .DIN2(n34191), .Q(n34197) );
  or2s1 U26574 ( .DIN1(n34199), .DIN2(n34175), .Q(n34191) );
  and2s1 U26575 ( .DIN1(n34168), .DIN2(n34200), .Q(n34199) );
  and2s1 U26576 ( .DIN1(n34168), .DIN2(n34194), .Q(n34198) );
  and2s1 U26577 ( .DIN1(n34201), .DIN2(n34202), .Q(n34195) );
  and2s1 U26578 ( .DIN1(n34193), .DIN2(n34203), .Q(n34202) );
  hi1s1 U26579 ( .DIN1(n34200), .Q(n34193) );
  and2s1 U26580 ( .DIN1(n34168), .DIN2(u4_rfr_cnt[3]), .Q(n34201) );
  or2s1 U26581 ( .DIN1(n34204), .DIN2(n34205), .Q(n9398) );
  and2s1 U26582 ( .DIN1(u4_rfr_cnt[5]), .DIN2(n34206), .Q(n34205) );
  and2s1 U26583 ( .DIN1(n34207), .DIN2(n34208), .Q(n34204) );
  or2s1 U26584 ( .DIN1(n34209), .DIN2(n34210), .Q(n9397) );
  and2s1 U26585 ( .DIN1(u4_rfr_cnt[6]), .DIN2(n34167), .Q(n34210) );
  or2s1 U26586 ( .DIN1(n34207), .DIN2(n34206), .Q(n34167) );
  or2s1 U26587 ( .DIN1(n34211), .DIN2(n34175), .Q(n34206) );
  and2s1 U26588 ( .DIN1(n34126), .DIN2(n34212), .Q(n34175) );
  hi1s1 U26589 ( .DIN1(n36610), .Q(n34212) );
  and2s1 U26590 ( .DIN1(n34168), .DIN2(n34213), .Q(n34211) );
  and2s1 U26591 ( .DIN1(n34168), .DIN2(n34214), .Q(n34207) );
  hi1s1 U26592 ( .DIN1(u4_rfr_cnt[5]), .Q(n34214) );
  and2s1 U26593 ( .DIN1(n34171), .DIN2(n34169), .Q(n34209) );
  hi1s1 U26594 ( .DIN1(u4_rfr_cnt[6]), .Q(n34169) );
  and2s1 U26595 ( .DIN1(u4_rfr_cnt[5]), .DIN2(n34215), .Q(n34171) );
  and2s1 U26596 ( .DIN1(n34168), .DIN2(n34208), .Q(n34215) );
  hi1s1 U26597 ( .DIN1(n34213), .Q(n34208) );
  or2s1 U26598 ( .DIN1(n34203), .DIN2(n34216), .Q(n34213) );
  or2s1 U26599 ( .DIN1(n34200), .DIN2(n34194), .Q(n34216) );
  hi1s1 U26600 ( .DIN1(u4_rfr_cnt[3]), .Q(n34194) );
  or2s1 U26601 ( .DIN1(n34188), .DIN2(n34217), .Q(n34200) );
  or2s1 U26602 ( .DIN1(n34185), .DIN2(n34180), .Q(n34217) );
  hi1s1 U26603 ( .DIN1(u4_rfr_cnt[1]), .Q(n34180) );
  hi1s1 U26604 ( .DIN1(u4_rfr_cnt[0]), .Q(n34185) );
  hi1s1 U26605 ( .DIN1(u4_rfr_cnt[2]), .Q(n34188) );
  hi1s1 U26606 ( .DIN1(u4_rfr_cnt[4]), .Q(n34203) );
  and2s1 U26607 ( .DIN1(n34126), .DIN2(n36610), .Q(n34168) );
  and2s1 U26608 ( .DIN1(n34218), .DIN2(u4_rfr_cnt[0]), .Q(n9396) );
  and2s1 U26609 ( .DIN1(n34219), .DIN2(n4612), .Q(n34218) );
  or2s1 U26610 ( .DIN1(n34220), .DIN2(n34221), .Q(n34219) );
  and2s1 U26611 ( .DIN1(n34222), .DIN2(u4_rfr_cnt[2]), .Q(n34221) );
  and2s1 U26612 ( .DIN1(u4_rfr_cnt[1]), .DIN2(n34223), .Q(n34222) );
  or2s1 U26613 ( .DIN1(n34224), .DIN2(n34225), .Q(n34223) );
  and2s1 U26614 ( .DIN1(n34226), .DIN2(n34227), .Q(n34225) );
  and2s1 U26615 ( .DIN1(u4_rfr_cnt[3]), .DIN2(n34228), .Q(n34224) );
  or2s1 U26616 ( .DIN1(n34229), .DIN2(n34226), .Q(n34228) );
  and2s1 U26617 ( .DIN1(u4_rfr_cnt[4]), .DIN2(n34230), .Q(n34229) );
  or2s1 U26618 ( .DIN1(n34231), .DIN2(n34232), .Q(n34230) );
  and2s1 U26619 ( .DIN1(n34227), .DIN2(n34233), .Q(n34232) );
  and2s1 U26620 ( .DIN1(u4_rfr_cnt[5]), .DIN2(n34234), .Q(n34231) );
  or2s1 U26621 ( .DIN1(n34235), .DIN2(n34233), .Q(n34234) );
  and2s1 U26622 ( .DIN1(u4_rfr_cnt[6]), .DIN2(n34236), .Q(n34235) );
  or2s1 U26623 ( .DIN1(u4_rfr_cnt[7]), .DIN2(n34227), .Q(n34236) );
  and2s1 U26624 ( .DIN1(n34237), .DIN2(n34238), .Q(n34220) );
  or2s1 U26625 ( .DIN1(u4_rfr_cnt[1]), .DIN2(n34227), .Q(n34238) );
  hi1s1 U26626 ( .DIN1(u0_csr_r[8]), .Q(n34227) );
  and2s1 U26627 ( .DIN1(n34226), .DIN2(n34233), .Q(n34237) );
  hi1s1 U26628 ( .DIN1(u0_csr_r[9]), .Q(n34233) );
  hi1s1 U26629 ( .DIN1(u0_csr_r[10]), .Q(n34226) );
  and2s1 U26630 ( .DIN1(n34239), .DIN2(n34126), .Q(n9395) );
  or2s1 U26631 ( .DIN1(u4_rfr_req), .DIN2(n4611), .Q(n34239) );
  or2s1 U26632 ( .DIN1(n34240), .DIN2(n34241), .Q(n9394) );
  and2s1 U26633 ( .DIN1(u5_state[21]), .DIN2(n32844), .Q(n34240) );
  or2s1 U26634 ( .DIN1(n34242), .DIN2(n34243), .Q(n9393) );
  and2s1 U26635 ( .DIN1(u5_state[22]), .DIN2(n32844), .Q(n34242) );
  or2s1 U26636 ( .DIN1(n34244), .DIN2(n34245), .Q(n9392) );
  and2s1 U26637 ( .DIN1(n32878), .DIN2(n34129), .Q(n34245) );
  hi1s1 U26638 ( .DIN1(n15513), .Q(n34129) );
  and2s1 U26639 ( .DIN1(u5_state[61]), .DIN2(n32844), .Q(n34244) );
  or2s1 U26640 ( .DIN1(n34246), .DIN2(n34247), .Q(n9391) );
  and2s1 U26641 ( .DIN1(u5_state[46]), .DIN2(n32844), .Q(n34246) );
  or2s1 U26642 ( .DIN1(n34248), .DIN2(n34249), .Q(n9390) );
  and2s1 U26643 ( .DIN1(u5_state[48]), .DIN2(n32844), .Q(n34248) );
  or2s1 U26644 ( .DIN1(n34250), .DIN2(n34251), .Q(n9389) );
  and2s1 U26645 ( .DIN1(u5_state[49]), .DIN2(n32855), .Q(n34250) );
  or2s1 U26646 ( .DIN1(n34252), .DIN2(n34253), .Q(n9388) );
  and2s1 U26647 ( .DIN1(u5_state[5]), .DIN2(n32965), .Q(n34253) );
  and2s1 U26648 ( .DIN1(n34254), .DIN2(n32921), .Q(n34252) );
  or2s1 U26649 ( .DIN1(n34255), .DIN2(n34256), .Q(n9387) );
  and2s1 U26650 ( .DIN1(u5_resume_req_r), .DIN2(n34257), .Q(n34256) );
  and2s1 U26651 ( .DIN1(u5_state[31]), .DIN2(n32855), .Q(n34255) );
  or2s1 U26652 ( .DIN1(n34258), .DIN2(n34259), .Q(n32855) );
  or2s1 U26653 ( .DIN1(n34260), .DIN2(n34261), .Q(n9386) );
  and2s1 U26654 ( .DIN1(u5_state[34]), .DIN2(n32844), .Q(n34260) );
  or2s1 U26655 ( .DIN1(n34262), .DIN2(n34263), .Q(n9385) );
  and2s1 U26656 ( .DIN1(u5_state[35]), .DIN2(n32844), .Q(n34262) );
  or2s1 U26657 ( .DIN1(n34264), .DIN2(n34265), .Q(n9384) );
  and2s1 U26658 ( .DIN1(u5_state[28]), .DIN2(n32965), .Q(n34265) );
  and2s1 U26659 ( .DIN1(n34266), .DIN2(n34267), .Q(n34264) );
  and2s1 U26660 ( .DIN1(n34268), .DIN2(n32921), .Q(n34267) );
  or2s1 U26661 ( .DIN1(n34269), .DIN2(n34270), .Q(n9383) );
  and2s1 U26662 ( .DIN1(u5_state[24]), .DIN2(n32925), .Q(n34270) );
  and2s1 U26663 ( .DIN1(u5_tmr_done), .DIN2(n34271), .Q(n34269) );
  or2s1 U26664 ( .DIN1(n34272), .DIN2(n34273), .Q(n34271) );
  and2s1 U26665 ( .DIN1(n15507), .DIN2(n34274), .Q(n34272) );
  or2s1 U26666 ( .DIN1(n34275), .DIN2(n34276), .Q(n9382) );
  and2s1 U26667 ( .DIN1(u5_state[26]), .DIN2(n32844), .Q(n34276) );
  and2s1 U26668 ( .DIN1(n34277), .DIN2(n34274), .Q(n34275) );
  and2s1 U26669 ( .DIN1(u5_tmr_done), .DIN2(n34278), .Q(n34277) );
  hi1s1 U26670 ( .DIN1(n15507), .Q(n34278) );
  or2s1 U26671 ( .DIN1(n34279), .DIN2(n34280), .Q(n9381) );
  and2s1 U26672 ( .DIN1(u5_state[18]), .DIN2(n32844), .Q(n34279) );
  or2s1 U26673 ( .DIN1(n34281), .DIN2(n34282), .Q(n9380) );
  and2s1 U26674 ( .DIN1(n34283), .DIN2(n32921), .Q(n34282) );
  and2s1 U26675 ( .DIN1(u5_state[19]), .DIN2(n32965), .Q(n34281) );
  or2s1 U26676 ( .DIN1(n34284), .DIN2(n34285), .Q(n32965) );
  or2s1 U26677 ( .DIN1(n34286), .DIN2(n34287), .Q(n9379) );
  and2s1 U26678 ( .DIN1(n32868), .DIN2(u5_tmr_done), .Q(n34287) );
  and2s1 U26679 ( .DIN1(u5_state[20]), .DIN2(n32925), .Q(n34286) );
  or2s1 U26680 ( .DIN1(n34288), .DIN2(n34289), .Q(n9378) );
  or2s1 U26681 ( .DIN1(n32868), .DIN2(n34290), .Q(n34289) );
  or2s1 U26682 ( .DIN1(n34283), .DIN2(n34280), .Q(n34288) );
  or2s1 U26683 ( .DIN1(n34291), .DIN2(n34292), .Q(n9377) );
  or2s1 U26684 ( .DIN1(n34293), .DIN2(n34294), .Q(n34292) );
  and2s1 U26685 ( .DIN1(n34295), .DIN2(u5_tmr2_done), .Q(n34294) );
  and2s1 U26686 ( .DIN1(n34296), .DIN2(n32849), .Q(n34293) );
  and2s1 U26687 ( .DIN1(u5_tmr2_done), .DIN2(n34297), .Q(n32849) );
  and2s1 U26688 ( .DIN1(u5_state[45]), .DIN2(n32925), .Q(n34291) );
  or2s1 U26689 ( .DIN1(n34298), .DIN2(n34299), .Q(n9376) );
  hi1s1 U26690 ( .DIN1(n34300), .Q(n34299) );
  or2s1 U26691 ( .DIN1(n34301), .DIN2(n15483), .Q(n34300) );
  and2s1 U26692 ( .DIN1(n34302), .DIN2(n34301), .Q(n34298) );
  or2s1 U26693 ( .DIN1(n34303), .DIN2(n4991), .Q(n34301) );
  and2s1 U26694 ( .DIN1(n34304), .DIN2(n33930), .Q(n34302) );
  or2s1 U26695 ( .DIN1(n33937), .DIN2(n33918), .Q(n34304) );
  or2s1 U26696 ( .DIN1(n34305), .DIN2(n34306), .Q(n9375) );
  hi1s1 U26697 ( .DIN1(n34307), .Q(n34306) );
  or2s1 U26698 ( .DIN1(n34308), .DIN2(n15510), .Q(n34307) );
  and2s1 U26699 ( .DIN1(n34309), .DIN2(n34308), .Q(n34305) );
  or2s1 U26700 ( .DIN1(n34310), .DIN2(n4992), .Q(n34308) );
  and2s1 U26701 ( .DIN1(n34311), .DIN2(n33946), .Q(n34309) );
  or2s1 U26702 ( .DIN1(n33952), .DIN2(n33918), .Q(n34311) );
  or2s1 U26703 ( .DIN1(u5_lmr_ack), .DIN2(n4988), .Q(n33918) );
  or2s1 U26704 ( .DIN1(n33946), .DIN2(n33930), .Q(n9374) );
  hi1s1 U26705 ( .DIN1(n36611), .Q(n33930) );
  hi1s1 U26706 ( .DIN1(n15506), .Q(n33946) );
  or2s1 U26707 ( .DIN1(n34312), .DIN2(n34313), .Q(n9373) );
  and2s1 U26708 ( .DIN1(u5_state[33]), .DIN2(n32988), .Q(n34313) );
  hi1s1 U26709 ( .DIN1(n34314), .Q(n34312) );
  or2s1 U26710 ( .DIN1(n32871), .DIN2(n34315), .Q(n34314) );
  or2s1 U26711 ( .DIN1(n32979), .DIN2(n34316), .Q(n32871) );
  or2s1 U26712 ( .DIN1(u5_cmd_asserted2), .DIN2(n34317), .Q(n34316) );
  hi1s1 U26713 ( .DIN1(n34318), .Q(n34317) );
  or2s1 U26714 ( .DIN1(n34319), .DIN2(n34320), .Q(n9372) );
  hi1s1 U26715 ( .DIN1(n34321), .Q(n34319) );
  or2s1 U26716 ( .DIN1(n34322), .DIN2(n34323), .Q(n34321) );
  and2s1 U26717 ( .DIN1(n32921), .DIN2(n34324), .Q(n34323) );
  or2s1 U26718 ( .DIN1(n34325), .DIN2(n34320), .Q(n9371) );
  and2s1 U26719 ( .DIN1(u5_state[27]), .DIN2(n32844), .Q(n34325) );
  or2s1 U26720 ( .DIN1(n34326), .DIN2(n34327), .Q(n9370) );
  and2s1 U26721 ( .DIN1(u5_state[4]), .DIN2(n32844), .Q(n34326) );
  or2s1 U26722 ( .DIN1(n34328), .DIN2(n34329), .Q(n9369) );
  and2s1 U26723 ( .DIN1(u5_ap_en), .DIN2(n34315), .Q(n34329) );
  and2s1 U26724 ( .DIN1(n34330), .DIN2(n34331), .Q(n34328) );
  and2s1 U26725 ( .DIN1(n32962), .DIN2(n32870), .Q(n34330) );
  or2s1 U26726 ( .DIN1(n34332), .DIN2(n34333), .Q(n9368) );
  and2s1 U26727 ( .DIN1(u5_state[62]), .DIN2(n32925), .Q(n34332) );
  or2s1 U26728 ( .DIN1(n34334), .DIN2(n33013), .Q(n9367) );
  and2s1 U26729 ( .DIN1(u5_state[32]), .DIN2(n32844), .Q(n34334) );
  or2s1 U26730 ( .DIN1(n34285), .DIN2(n32925), .Q(n32844) );
  or2s1 U26731 ( .DIN1(n34335), .DIN2(n32988), .Q(n32925) );
  or2s1 U26732 ( .DIN1(n34284), .DIN2(n34336), .Q(n32988) );
  or2s1 U26733 ( .DIN1(n34337), .DIN2(n34338), .Q(n34284) );
  or2s1 U26734 ( .DIN1(n34162), .DIN2(n34339), .Q(n34338) );
  or2s1 U26735 ( .DIN1(n34340), .DIN2(n34341), .Q(n34162) );
  hi1s1 U26736 ( .DIN1(n34342), .Q(n34340) );
  or2s1 U26737 ( .DIN1(n34343), .DIN2(u5_resume_req_r), .Q(n34342) );
  or2s1 U26738 ( .DIN1(n34344), .DIN2(n34345), .Q(n34337) );
  and2s1 U26739 ( .DIN1(n15512), .DIN2(n34346), .Q(n34345) );
  or2s1 U26740 ( .DIN1(n34347), .DIN2(n34348), .Q(n34346) );
  and2s1 U26741 ( .DIN1(n34349), .DIN2(n34350), .Q(n34344) );
  or2s1 U26742 ( .DIN1(n34351), .DIN2(n32856), .Q(n34349) );
  and2s1 U26743 ( .DIN1(n15512), .DIN2(n34352), .Q(n34335) );
  or2s1 U26744 ( .DIN1(n34258), .DIN2(n34353), .Q(n34285) );
  or2s1 U26745 ( .DIN1(n34354), .DIN2(n34355), .Q(n34353) );
  and2s1 U26746 ( .DIN1(u7_mc_br_r), .DIN2(n34356), .Q(n34354) );
  or2s1 U26747 ( .DIN1(n34357), .DIN2(n32865), .Q(n34356) );
  and2s1 U26748 ( .DIN1(n34358), .DIN2(u5_cmd_asserted2), .Q(n34357) );
  and2s1 U26749 ( .DIN1(n34318), .DIN2(n32870), .Q(n34358) );
  or2s1 U26750 ( .DIN1(n34359), .DIN2(n34360), .Q(n34258) );
  and2s1 U26751 ( .DIN1(n34361), .DIN2(n34350), .Q(n34360) );
  and2s1 U26752 ( .DIN1(n34362), .DIN2(n34363), .Q(n34359) );
  or2s1 U26753 ( .DIN1(n34364), .DIN2(n34365), .Q(n34362) );
  or2s1 U26754 ( .DIN1(n32868), .DIN2(n34366), .Q(n34365) );
  or2s1 U26755 ( .DIN1(n33492), .DIN2(n34367), .Q(n34364) );
  or2s1 U26756 ( .DIN1(n34273), .DIN2(n34368), .Q(n34367) );
  or2s1 U26757 ( .DIN1(n34369), .DIN2(n34102), .Q(n9365) );
  and2s1 U26758 ( .DIN1(n34247), .DIN2(n34296), .Q(n34369) );
  or2s1 U26759 ( .DIN1(n34370), .DIN2(n34371), .Q(n9364) );
  and2s1 U26760 ( .DIN1(n15504), .DIN2(n34372), .Q(n34371) );
  and2s1 U26761 ( .DIN1(n34373), .DIN2(n32837), .Q(n34370) );
  or2s1 U26762 ( .DIN1(n34374), .DIN2(n34375), .Q(n9363) );
  or2s1 U26763 ( .DIN1(n34376), .DIN2(n34377), .Q(n34375) );
  and2s1 U26764 ( .DIN1(n33674), .DIN2(n9061), .Q(n34377) );
  and2s1 U26765 ( .DIN1(n33675), .DIN2(n9059), .Q(n34376) );
  or2s1 U26766 ( .DIN1(n34378), .DIN2(n34379), .Q(n34374) );
  and2s1 U26767 ( .DIN1(n33682), .DIN2(n32837), .Q(n34379) );
  and2s1 U26768 ( .DIN1(n34380), .DIN2(n34372), .Q(n34378) );
  hi1s1 U26769 ( .DIN1(n36612), .Q(n34372) );
  or2s1 U26770 ( .DIN1(n34381), .DIN2(n34382), .Q(n9362) );
  and2s1 U26771 ( .DIN1(n15504), .DIN2(n34383), .Q(n34382) );
  and2s1 U26772 ( .DIN1(n34373), .DIN2(n32829), .Q(n34381) );
  or2s1 U26773 ( .DIN1(n34384), .DIN2(n34385), .Q(n9361) );
  or2s1 U26774 ( .DIN1(n34386), .DIN2(n34387), .Q(n34385) );
  and2s1 U26775 ( .DIN1(n33674), .DIN2(n9063), .Q(n34387) );
  and2s1 U26776 ( .DIN1(n33675), .DIN2(n9058), .Q(n34386) );
  or2s1 U26777 ( .DIN1(n34388), .DIN2(n34389), .Q(n34384) );
  and2s1 U26778 ( .DIN1(n33682), .DIN2(n32829), .Q(n34389) );
  and2s1 U26779 ( .DIN1(n34380), .DIN2(n34383), .Q(n34388) );
  hi1s1 U26780 ( .DIN1(n36613), .Q(n34383) );
  or2s1 U26781 ( .DIN1(n34390), .DIN2(n34391), .Q(n9360) );
  and2s1 U26782 ( .DIN1(n15504), .DIN2(n34392), .Q(n34391) );
  and2s1 U26783 ( .DIN1(n34373), .DIN2(n32740), .Q(n34390) );
  or2s1 U26784 ( .DIN1(n34393), .DIN2(n34394), .Q(n9359) );
  or2s1 U26785 ( .DIN1(n34395), .DIN2(n34396), .Q(n34394) );
  and2s1 U26786 ( .DIN1(n33674), .DIN2(n9064), .Q(n34396) );
  and2s1 U26787 ( .DIN1(n33675), .DIN2(n9057), .Q(n34395) );
  or2s1 U26788 ( .DIN1(n34397), .DIN2(n34398), .Q(n34393) );
  and2s1 U26789 ( .DIN1(n33682), .DIN2(n32740), .Q(n34398) );
  and2s1 U26790 ( .DIN1(n34380), .DIN2(n34392), .Q(n34397) );
  hi1s1 U26791 ( .DIN1(n36614), .Q(n34392) );
  or2s1 U26792 ( .DIN1(n34399), .DIN2(n34400), .Q(n9358) );
  and2s1 U26793 ( .DIN1(n15504), .DIN2(n34401), .Q(n34400) );
  and2s1 U26794 ( .DIN1(n34373), .DIN2(n32733), .Q(n34399) );
  or2s1 U26795 ( .DIN1(n34402), .DIN2(n34403), .Q(n9357) );
  or2s1 U26796 ( .DIN1(n34404), .DIN2(n34405), .Q(n34403) );
  and2s1 U26797 ( .DIN1(n33674), .DIN2(n9065), .Q(n34405) );
  and2s1 U26798 ( .DIN1(n33675), .DIN2(n9056), .Q(n34404) );
  or2s1 U26799 ( .DIN1(n34406), .DIN2(n34407), .Q(n34402) );
  and2s1 U26800 ( .DIN1(n33682), .DIN2(n32733), .Q(n34407) );
  and2s1 U26801 ( .DIN1(n34380), .DIN2(n34401), .Q(n34406) );
  hi1s1 U26802 ( .DIN1(n36615), .Q(n34401) );
  or2s1 U26803 ( .DIN1(n34408), .DIN2(n34409), .Q(n9356) );
  and2s1 U26804 ( .DIN1(n15504), .DIN2(n34410), .Q(n34409) );
  and2s1 U26805 ( .DIN1(n34373), .DIN2(n32730), .Q(n34408) );
  or2s1 U26806 ( .DIN1(n34411), .DIN2(n34412), .Q(n9355) );
  or2s1 U26807 ( .DIN1(n34413), .DIN2(n34414), .Q(n34412) );
  and2s1 U26808 ( .DIN1(n33674), .DIN2(n9060), .Q(n34414) );
  and2s1 U26809 ( .DIN1(n33675), .DIN2(n9055), .Q(n34413) );
  or2s1 U26810 ( .DIN1(n34415), .DIN2(n34416), .Q(n34411) );
  and2s1 U26811 ( .DIN1(n33682), .DIN2(n32730), .Q(n34416) );
  and2s1 U26812 ( .DIN1(n34380), .DIN2(n34410), .Q(n34415) );
  hi1s1 U26813 ( .DIN1(n36616), .Q(n34410) );
  or2s1 U26814 ( .DIN1(n34417), .DIN2(n34418), .Q(n9354) );
  and2s1 U26815 ( .DIN1(n15504), .DIN2(n34419), .Q(n34418) );
  and2s1 U26816 ( .DIN1(n34373), .DIN2(n32727), .Q(n34417) );
  or2s1 U26817 ( .DIN1(n34420), .DIN2(n34421), .Q(n9353) );
  or2s1 U26818 ( .DIN1(n34422), .DIN2(n34423), .Q(n34421) );
  and2s1 U26819 ( .DIN1(n33674), .DIN2(n9062), .Q(n34423) );
  and2s1 U26820 ( .DIN1(n33675), .DIN2(n9054), .Q(n34422) );
  or2s1 U26821 ( .DIN1(n34424), .DIN2(n34425), .Q(n34420) );
  and2s1 U26822 ( .DIN1(n33682), .DIN2(n32727), .Q(n34425) );
  and2s1 U26823 ( .DIN1(n34380), .DIN2(n34419), .Q(n34424) );
  hi1s1 U26824 ( .DIN1(n36617), .Q(n34419) );
  or2s1 U26825 ( .DIN1(n34426), .DIN2(n34427), .Q(n9352) );
  and2s1 U26826 ( .DIN1(n15504), .DIN2(n34428), .Q(n34427) );
  and2s1 U26827 ( .DIN1(n34373), .DIN2(n32724), .Q(n34426) );
  or2s1 U26828 ( .DIN1(n34429), .DIN2(n34430), .Q(n9351) );
  or2s1 U26829 ( .DIN1(n34431), .DIN2(n34432), .Q(n34430) );
  and2s1 U26830 ( .DIN1(n33674), .DIN2(n9066), .Q(n34432) );
  and2s1 U26831 ( .DIN1(n33675), .DIN2(n9053), .Q(n34431) );
  or2s1 U26832 ( .DIN1(n34433), .DIN2(n34434), .Q(n34429) );
  and2s1 U26833 ( .DIN1(n33682), .DIN2(n32724), .Q(n34434) );
  and2s1 U26834 ( .DIN1(n34380), .DIN2(n34428), .Q(n34433) );
  hi1s1 U26835 ( .DIN1(n36618), .Q(n34428) );
  or2s1 U26836 ( .DIN1(n34435), .DIN2(n34436), .Q(n9350) );
  and2s1 U26837 ( .DIN1(n15504), .DIN2(n34437), .Q(n34436) );
  and2s1 U26838 ( .DIN1(n34373), .DIN2(n32721), .Q(n34435) );
  hi1s1 U26839 ( .DIN1(n15504), .Q(n34373) );
  or2s1 U26840 ( .DIN1(n34438), .DIN2(n34439), .Q(n9349) );
  or2s1 U26841 ( .DIN1(n34440), .DIN2(n34441), .Q(n34439) );
  and2s1 U26842 ( .DIN1(n33674), .DIN2(n9067), .Q(n34441) );
  and2s1 U26843 ( .DIN1(n33675), .DIN2(n9052), .Q(n34440) );
  or2s1 U26844 ( .DIN1(n34442), .DIN2(n34443), .Q(n34438) );
  and2s1 U26845 ( .DIN1(n33682), .DIN2(n32721), .Q(n34443) );
  and2s1 U26846 ( .DIN1(n34380), .DIN2(n34437), .Q(n34442) );
  hi1s1 U26847 ( .DIN1(n36619), .Q(n34437) );
  and2s1 U26848 ( .DIN1(n34247), .DIN2(n34100), .Q(n9348) );
  or2s1 U26849 ( .DIN1(n34444), .DIN2(n34445), .Q(n9347) );
  and2s1 U26850 ( .DIN1(n15503), .DIN2(n34446), .Q(n34445) );
  and2s1 U26851 ( .DIN1(n34447), .DIN2(n32837), .Q(n34444) );
  or2s1 U26852 ( .DIN1(n34448), .DIN2(n34449), .Q(n9346) );
  or2s1 U26853 ( .DIN1(n34450), .DIN2(n34451), .Q(n34449) );
  and2s1 U26854 ( .DIN1(n33674), .DIN2(n9076), .Q(n34451) );
  and2s1 U26855 ( .DIN1(n33675), .DIN2(n9043), .Q(n34450) );
  or2s1 U26856 ( .DIN1(n34452), .DIN2(n34453), .Q(n34448) );
  or2s1 U26857 ( .DIN1(n34454), .DIN2(n34455), .Q(n34453) );
  and2s1 U26858 ( .DIN1(n33680), .DIN2(n34446), .Q(n34455) );
  hi1s1 U26859 ( .DIN1(n36621), .Q(n34446) );
  and2s1 U26860 ( .DIN1(n33681), .DIN2(n32837), .Q(n34454) );
  and2s1 U26861 ( .DIN1(n33682), .DIN2(n32694), .Q(n34452) );
  hi1s1 U26862 ( .DIN1(n36620), .Q(n32694) );
  or2s1 U26863 ( .DIN1(n34456), .DIN2(n34457), .Q(n9345) );
  and2s1 U26864 ( .DIN1(n15503), .DIN2(n34458), .Q(n34457) );
  and2s1 U26865 ( .DIN1(n34447), .DIN2(n32829), .Q(n34456) );
  or2s1 U26866 ( .DIN1(n34459), .DIN2(n34460), .Q(n9344) );
  or2s1 U26867 ( .DIN1(n34461), .DIN2(n34462), .Q(n34460) );
  and2s1 U26868 ( .DIN1(n33674), .DIN2(n9077), .Q(n34462) );
  and2s1 U26869 ( .DIN1(n33675), .DIN2(n9042), .Q(n34461) );
  or2s1 U26870 ( .DIN1(n34463), .DIN2(n34464), .Q(n34459) );
  or2s1 U26871 ( .DIN1(n34465), .DIN2(n34466), .Q(n34464) );
  and2s1 U26872 ( .DIN1(n33680), .DIN2(n34458), .Q(n34466) );
  hi1s1 U26873 ( .DIN1(n36623), .Q(n34458) );
  and2s1 U26874 ( .DIN1(n33681), .DIN2(n32829), .Q(n34465) );
  and2s1 U26875 ( .DIN1(n33682), .DIN2(n32691), .Q(n34463) );
  hi1s1 U26876 ( .DIN1(n36622), .Q(n32691) );
  or2s1 U26877 ( .DIN1(n34467), .DIN2(n34468), .Q(n9343) );
  and2s1 U26878 ( .DIN1(n15503), .DIN2(n34469), .Q(n34468) );
  and2s1 U26879 ( .DIN1(n34447), .DIN2(n32740), .Q(n34467) );
  or2s1 U26880 ( .DIN1(n34470), .DIN2(n34471), .Q(n9342) );
  or2s1 U26881 ( .DIN1(n34472), .DIN2(n34473), .Q(n34471) );
  and2s1 U26882 ( .DIN1(n33674), .DIN2(n9078), .Q(n34473) );
  and2s1 U26883 ( .DIN1(n33675), .DIN2(n9041), .Q(n34472) );
  or2s1 U26884 ( .DIN1(n34474), .DIN2(n34475), .Q(n34470) );
  or2s1 U26885 ( .DIN1(n34476), .DIN2(n34477), .Q(n34475) );
  and2s1 U26886 ( .DIN1(n33680), .DIN2(n34469), .Q(n34477) );
  hi1s1 U26887 ( .DIN1(n36625), .Q(n34469) );
  and2s1 U26888 ( .DIN1(n33681), .DIN2(n32740), .Q(n34476) );
  and2s1 U26889 ( .DIN1(n33682), .DIN2(n32688), .Q(n34474) );
  hi1s1 U26890 ( .DIN1(n36624), .Q(n32688) );
  or2s1 U26891 ( .DIN1(n34478), .DIN2(n34479), .Q(n9341) );
  and2s1 U26892 ( .DIN1(n15503), .DIN2(n34480), .Q(n34479) );
  and2s1 U26893 ( .DIN1(n34447), .DIN2(n32733), .Q(n34478) );
  or2s1 U26894 ( .DIN1(n34481), .DIN2(n34482), .Q(n9340) );
  or2s1 U26895 ( .DIN1(n34483), .DIN2(n34484), .Q(n34482) );
  and2s1 U26896 ( .DIN1(n33674), .DIN2(n9079), .Q(n34484) );
  and2s1 U26897 ( .DIN1(n33675), .DIN2(n9040), .Q(n34483) );
  or2s1 U26898 ( .DIN1(n34485), .DIN2(n34486), .Q(n34481) );
  or2s1 U26899 ( .DIN1(n34487), .DIN2(n34488), .Q(n34486) );
  and2s1 U26900 ( .DIN1(n33680), .DIN2(n34480), .Q(n34488) );
  hi1s1 U26901 ( .DIN1(n36627), .Q(n34480) );
  and2s1 U26902 ( .DIN1(n33681), .DIN2(n32733), .Q(n34487) );
  and2s1 U26903 ( .DIN1(n33682), .DIN2(n32685), .Q(n34485) );
  hi1s1 U26904 ( .DIN1(n36626), .Q(n32685) );
  or2s1 U26905 ( .DIN1(n34489), .DIN2(n34490), .Q(n9339) );
  and2s1 U26906 ( .DIN1(n15503), .DIN2(n34491), .Q(n34490) );
  and2s1 U26907 ( .DIN1(n34447), .DIN2(n32730), .Q(n34489) );
  or2s1 U26908 ( .DIN1(n34492), .DIN2(n34493), .Q(n9338) );
  or2s1 U26909 ( .DIN1(n34494), .DIN2(n34495), .Q(n34493) );
  and2s1 U26910 ( .DIN1(n33674), .DIN2(n9080), .Q(n34495) );
  and2s1 U26911 ( .DIN1(n33675), .DIN2(n9039), .Q(n34494) );
  or2s1 U26912 ( .DIN1(n34496), .DIN2(n34497), .Q(n34492) );
  or2s1 U26913 ( .DIN1(n34498), .DIN2(n34499), .Q(n34497) );
  and2s1 U26914 ( .DIN1(n33680), .DIN2(n34491), .Q(n34499) );
  hi1s1 U26915 ( .DIN1(n36629), .Q(n34491) );
  and2s1 U26916 ( .DIN1(n33681), .DIN2(n32730), .Q(n34498) );
  and2s1 U26917 ( .DIN1(n33682), .DIN2(n32682), .Q(n34496) );
  hi1s1 U26918 ( .DIN1(n36628), .Q(n32682) );
  or2s1 U26919 ( .DIN1(n34500), .DIN2(n34501), .Q(n9337) );
  and2s1 U26920 ( .DIN1(n15503), .DIN2(n34502), .Q(n34501) );
  and2s1 U26921 ( .DIN1(n34447), .DIN2(n32727), .Q(n34500) );
  or2s1 U26922 ( .DIN1(n34503), .DIN2(n34504), .Q(n9336) );
  or2s1 U26923 ( .DIN1(n34505), .DIN2(n34506), .Q(n34504) );
  and2s1 U26924 ( .DIN1(n33674), .DIN2(n9081), .Q(n34506) );
  and2s1 U26925 ( .DIN1(n33675), .DIN2(n9038), .Q(n34505) );
  or2s1 U26926 ( .DIN1(n34507), .DIN2(n34508), .Q(n34503) );
  or2s1 U26927 ( .DIN1(n34509), .DIN2(n34510), .Q(n34508) );
  and2s1 U26928 ( .DIN1(n33680), .DIN2(n34502), .Q(n34510) );
  hi1s1 U26929 ( .DIN1(n36631), .Q(n34502) );
  and2s1 U26930 ( .DIN1(n33681), .DIN2(n32727), .Q(n34509) );
  and2s1 U26931 ( .DIN1(n33682), .DIN2(n32679), .Q(n34507) );
  hi1s1 U26932 ( .DIN1(n36630), .Q(n32679) );
  or2s1 U26933 ( .DIN1(n34511), .DIN2(n34512), .Q(n9335) );
  and2s1 U26934 ( .DIN1(n15503), .DIN2(n34513), .Q(n34512) );
  and2s1 U26935 ( .DIN1(n34447), .DIN2(n32724), .Q(n34511) );
  or2s1 U26936 ( .DIN1(n34514), .DIN2(n34515), .Q(n9334) );
  or2s1 U26937 ( .DIN1(n34516), .DIN2(n34517), .Q(n34515) );
  and2s1 U26938 ( .DIN1(n33674), .DIN2(n9082), .Q(n34517) );
  and2s1 U26939 ( .DIN1(n33675), .DIN2(n9037), .Q(n34516) );
  or2s1 U26940 ( .DIN1(n34518), .DIN2(n34519), .Q(n34514) );
  or2s1 U26941 ( .DIN1(n34520), .DIN2(n34521), .Q(n34519) );
  and2s1 U26942 ( .DIN1(n33680), .DIN2(n34513), .Q(n34521) );
  hi1s1 U26943 ( .DIN1(n36633), .Q(n34513) );
  and2s1 U26944 ( .DIN1(n33681), .DIN2(n32724), .Q(n34520) );
  and2s1 U26945 ( .DIN1(n33682), .DIN2(n32676), .Q(n34518) );
  hi1s1 U26946 ( .DIN1(n36632), .Q(n32676) );
  or2s1 U26947 ( .DIN1(n34522), .DIN2(n34523), .Q(n9333) );
  and2s1 U26948 ( .DIN1(n15503), .DIN2(n34524), .Q(n34523) );
  and2s1 U26949 ( .DIN1(n34447), .DIN2(n32721), .Q(n34522) );
  hi1s1 U26950 ( .DIN1(n15503), .Q(n34447) );
  or2s1 U26951 ( .DIN1(n34525), .DIN2(n34526), .Q(n9332) );
  or2s1 U26952 ( .DIN1(n34527), .DIN2(n34528), .Q(n34526) );
  and2s1 U26953 ( .DIN1(n33674), .DIN2(n9083), .Q(n34528) );
  and2s1 U26954 ( .DIN1(n33675), .DIN2(n9036), .Q(n34527) );
  or2s1 U26955 ( .DIN1(n34529), .DIN2(n34530), .Q(n34525) );
  or2s1 U26956 ( .DIN1(n34531), .DIN2(n34532), .Q(n34530) );
  and2s1 U26957 ( .DIN1(n33680), .DIN2(n34524), .Q(n34532) );
  hi1s1 U26958 ( .DIN1(n36635), .Q(n34524) );
  and2s1 U26959 ( .DIN1(n34533), .DIN2(n34380), .Q(n33680) );
  and2s1 U26960 ( .DIN1(n33681), .DIN2(n32721), .Q(n34531) );
  and2s1 U26961 ( .DIN1(u0_csc[4]), .DIN2(n34380), .Q(n33681) );
  and2s1 U26962 ( .DIN1(n33682), .DIN2(n32673), .Q(n34529) );
  hi1s1 U26963 ( .DIN1(n36634), .Q(n32673) );
  or2s1 U26964 ( .DIN1(n34534), .DIN2(n34535), .Q(n9331) );
  and2s1 U26965 ( .DIN1(n34536), .DIN2(n32921), .Q(n34535) );
  hi1s1 U26966 ( .DIN1(n15512), .Q(n32921) );
  and2s1 U26967 ( .DIN1(u5_state[7]), .DIN2(n34259), .Q(n34534) );
  or2s1 U26968 ( .DIN1(n34339), .DIN2(n34336), .Q(n34259) );
  or2s1 U26969 ( .DIN1(n34537), .DIN2(n34538), .Q(n34336) );
  or2s1 U26970 ( .DIN1(n34539), .DIN2(n34540), .Q(n34538) );
  and2s1 U26971 ( .DIN1(n33894), .DIN2(n34541), .Q(n34540) );
  hi1s1 U26972 ( .DIN1(n33895), .Q(n34541) );
  or2s1 U26973 ( .DIN1(n32938), .DIN2(n4625), .Q(n33895) );
  and2s1 U26974 ( .DIN1(u5_wb_wait_r), .DIN2(n34542), .Q(n34539) );
  or2s1 U26975 ( .DIN1(n34543), .DIN2(n33911), .Q(n34542) );
  and2s1 U26976 ( .DIN1(n33910), .DIN2(n33902), .Q(n34543) );
  and2s1 U26977 ( .DIN1(n33900), .DIN2(n34363), .Q(n34537) );
  or2s1 U26978 ( .DIN1(n34544), .DIN2(n34545), .Q(n33900) );
  or2s1 U26979 ( .DIN1(n34546), .DIN2(n34547), .Q(n34339) );
  or2s1 U26980 ( .DIN1(n34548), .DIN2(n34549), .Q(n34547) );
  or2s1 U26981 ( .DIN1(n34550), .DIN2(n34551), .Q(n34549) );
  and2s1 U26982 ( .DIN1(n15512), .DIN2(n32940), .Q(n34551) );
  and2s1 U26983 ( .DIN1(n34552), .DIN2(n34363), .Q(n34550) );
  or2s1 U26984 ( .DIN1(n34553), .DIN2(n34554), .Q(n34552) );
  or2s1 U26985 ( .DIN1(n33911), .DIN2(n34125), .Q(n34554) );
  or2s1 U26986 ( .DIN1(n34274), .DIN2(n33901), .Q(n34553) );
  or2s1 U26987 ( .DIN1(n34555), .DIN2(n34556), .Q(n34548) );
  and2s1 U26988 ( .DIN1(n34557), .DIN2(n34350), .Q(n34556) );
  or2s1 U26989 ( .DIN1(n34558), .DIN2(n34559), .Q(n34557) );
  or2s1 U26990 ( .DIN1(n34297), .DIN2(n34560), .Q(n34559) );
  and2s1 U26991 ( .DIN1(n15513), .DIN2(n33875), .Q(n34558) );
  and2s1 U26992 ( .DIN1(n33017), .DIN2(n32869), .Q(n34555) );
  or2s1 U26993 ( .DIN1(n34561), .DIN2(n34562), .Q(n34546) );
  or2s1 U26994 ( .DIN1(n34563), .DIN2(n34564), .Q(n34562) );
  and2s1 U26995 ( .DIN1(n32943), .DIN2(n34565), .Q(n34564) );
  or2s1 U26996 ( .DIN1(n34566), .DIN2(n34567), .Q(n34565) );
  and2s1 U26997 ( .DIN1(n32958), .DIN2(n32934), .Q(n34566) );
  and2s1 U26998 ( .DIN1(n34568), .DIN2(n34569), .Q(n32958) );
  hi1s1 U26999 ( .DIN1(n33001), .Q(n34568) );
  and2s1 U27000 ( .DIN1(n34570), .DIN2(n32938), .Q(n33001) );
  and2s1 U27001 ( .DIN1(n32960), .DIN2(n34571), .Q(n34563) );
  or2s1 U27002 ( .DIN1(n34572), .DIN2(n33473), .Q(n34571) );
  or2s1 U27003 ( .DIN1(n33466), .DIN2(n34573), .Q(n33473) );
  or2s1 U27004 ( .DIN1(u5_ack_cnt[3]), .DIN2(u5_ack_cnt[2]), .Q(n34573) );
  or2s1 U27005 ( .DIN1(u5_ack_cnt[0]), .DIN2(u5_ack_cnt[1]), .Q(n33466) );
  and2s1 U27006 ( .DIN1(u5_mem_ack_r), .DIN2(n33004), .Q(n34572) );
  or2s1 U27007 ( .DIN1(u5_ap_en), .DIN2(n33902), .Q(n33004) );
  or2s1 U27008 ( .DIN1(n34574), .DIN2(n34575), .Q(n34561) );
  and2s1 U27009 ( .DIN1(n34576), .DIN2(n34318), .Q(n34575) );
  and2s1 U27010 ( .DIN1(n34577), .DIN2(n34578), .Q(n34318) );
  and2s1 U27011 ( .DIN1(n34579), .DIN2(n34580), .Q(n34578) );
  and2s1 U27012 ( .DIN1(n32870), .DIN2(n32979), .Q(n34576) );
  hi1s1 U27013 ( .DIN1(u7_mc_br_r), .Q(n32979) );
  or2s1 U27014 ( .DIN1(n34581), .DIN2(n34582), .Q(n9330) );
  and2s1 U27015 ( .DIN1(n32970), .DIN2(n34583), .Q(n34582) );
  and2s1 U27016 ( .DIN1(n9764), .DIN2(n34584), .Q(n34581) );
  or2s1 U27017 ( .DIN1(n34585), .DIN2(n34586), .Q(n9329) );
  and2s1 U27018 ( .DIN1(n9764), .DIN2(n34583), .Q(n34586) );
  hi1s1 U27019 ( .DIN1(n36636), .Q(n34583) );
  and2s1 U27020 ( .DIN1(n32970), .DIN2(n34587), .Q(n34585) );
  or2s1 U27021 ( .DIN1(n34588), .DIN2(n34589), .Q(n9327) );
  or2s1 U27022 ( .DIN1(n34590), .DIN2(n34591), .Q(n34589) );
  and2s1 U27023 ( .DIN1(n34592), .DIN2(n32837), .Q(n34591) );
  hi1s1 U27024 ( .DIN1(n36637), .Q(n32837) );
  and2s1 U27025 ( .DIN1(n34593), .DIN2(n32718), .Q(n34590) );
  and2s1 U27026 ( .DIN1(n34594), .DIN2(n34595), .Q(n34588) );
  or2s1 U27027 ( .DIN1(n34596), .DIN2(n34597), .Q(n9326) );
  or2s1 U27028 ( .DIN1(n34598), .DIN2(n34599), .Q(n34597) );
  and2s1 U27029 ( .DIN1(n33674), .DIN2(n9068), .Q(n34599) );
  and2s1 U27030 ( .DIN1(n33675), .DIN2(n9051), .Q(n34598) );
  or2s1 U27031 ( .DIN1(n34600), .DIN2(n34601), .Q(n34596) );
  and2s1 U27032 ( .DIN1(n33682), .DIN2(n32718), .Q(n34601) );
  hi1s1 U27033 ( .DIN1(n36639), .Q(n32718) );
  and2s1 U27034 ( .DIN1(n34380), .DIN2(n34595), .Q(n34600) );
  hi1s1 U27035 ( .DIN1(n36638), .Q(n34595) );
  or2s1 U27036 ( .DIN1(n34602), .DIN2(n34603), .Q(n9325) );
  or2s1 U27037 ( .DIN1(n34604), .DIN2(n34605), .Q(n34603) );
  and2s1 U27038 ( .DIN1(n34592), .DIN2(n32829), .Q(n34605) );
  hi1s1 U27039 ( .DIN1(n36640), .Q(n32829) );
  and2s1 U27040 ( .DIN1(n34593), .DIN2(n32715), .Q(n34604) );
  and2s1 U27041 ( .DIN1(n34594), .DIN2(n34606), .Q(n34602) );
  or2s1 U27042 ( .DIN1(n34607), .DIN2(n34608), .Q(n9324) );
  or2s1 U27043 ( .DIN1(n34609), .DIN2(n34610), .Q(n34608) );
  and2s1 U27044 ( .DIN1(n33674), .DIN2(n9069), .Q(n34610) );
  and2s1 U27045 ( .DIN1(n33675), .DIN2(n9050), .Q(n34609) );
  or2s1 U27046 ( .DIN1(n34611), .DIN2(n34612), .Q(n34607) );
  and2s1 U27047 ( .DIN1(n33682), .DIN2(n32715), .Q(n34612) );
  hi1s1 U27048 ( .DIN1(n36642), .Q(n32715) );
  and2s1 U27049 ( .DIN1(n34380), .DIN2(n34606), .Q(n34611) );
  hi1s1 U27050 ( .DIN1(n36641), .Q(n34606) );
  or2s1 U27051 ( .DIN1(n34613), .DIN2(n34614), .Q(n9323) );
  or2s1 U27052 ( .DIN1(n34615), .DIN2(n34616), .Q(n34614) );
  and2s1 U27053 ( .DIN1(n34592), .DIN2(n32740), .Q(n34616) );
  hi1s1 U27054 ( .DIN1(n36643), .Q(n32740) );
  and2s1 U27055 ( .DIN1(n34593), .DIN2(n32712), .Q(n34615) );
  and2s1 U27056 ( .DIN1(n34594), .DIN2(n34617), .Q(n34613) );
  or2s1 U27057 ( .DIN1(n34618), .DIN2(n34619), .Q(n9322) );
  or2s1 U27058 ( .DIN1(n34620), .DIN2(n34621), .Q(n34619) );
  and2s1 U27059 ( .DIN1(n33674), .DIN2(n9070), .Q(n34621) );
  and2s1 U27060 ( .DIN1(n33675), .DIN2(n9049), .Q(n34620) );
  or2s1 U27061 ( .DIN1(n34622), .DIN2(n34623), .Q(n34618) );
  and2s1 U27062 ( .DIN1(n33682), .DIN2(n32712), .Q(n34623) );
  hi1s1 U27063 ( .DIN1(n36645), .Q(n32712) );
  and2s1 U27064 ( .DIN1(n34380), .DIN2(n34617), .Q(n34622) );
  hi1s1 U27065 ( .DIN1(n36644), .Q(n34617) );
  or2s1 U27066 ( .DIN1(n34624), .DIN2(n34625), .Q(n9321) );
  or2s1 U27067 ( .DIN1(n34626), .DIN2(n34627), .Q(n34625) );
  and2s1 U27068 ( .DIN1(n34592), .DIN2(n32733), .Q(n34627) );
  hi1s1 U27069 ( .DIN1(n36646), .Q(n32733) );
  and2s1 U27070 ( .DIN1(n34593), .DIN2(n32709), .Q(n34626) );
  and2s1 U27071 ( .DIN1(n34594), .DIN2(n34628), .Q(n34624) );
  or2s1 U27072 ( .DIN1(n34629), .DIN2(n34630), .Q(n9320) );
  or2s1 U27073 ( .DIN1(n34631), .DIN2(n34632), .Q(n34630) );
  and2s1 U27074 ( .DIN1(n33674), .DIN2(n9071), .Q(n34632) );
  and2s1 U27075 ( .DIN1(n33675), .DIN2(n9048), .Q(n34631) );
  or2s1 U27076 ( .DIN1(n34633), .DIN2(n34634), .Q(n34629) );
  and2s1 U27077 ( .DIN1(n33682), .DIN2(n32709), .Q(n34634) );
  hi1s1 U27078 ( .DIN1(n36648), .Q(n32709) );
  and2s1 U27079 ( .DIN1(n34380), .DIN2(n34628), .Q(n34633) );
  hi1s1 U27080 ( .DIN1(n36647), .Q(n34628) );
  or2s1 U27081 ( .DIN1(n34635), .DIN2(n34636), .Q(n9319) );
  or2s1 U27082 ( .DIN1(n34637), .DIN2(n34638), .Q(n34636) );
  and2s1 U27083 ( .DIN1(n34592), .DIN2(n32730), .Q(n34638) );
  hi1s1 U27084 ( .DIN1(n36649), .Q(n32730) );
  and2s1 U27085 ( .DIN1(n34593), .DIN2(n32706), .Q(n34637) );
  and2s1 U27086 ( .DIN1(n34594), .DIN2(n34639), .Q(n34635) );
  or2s1 U27087 ( .DIN1(n34640), .DIN2(n34641), .Q(n9318) );
  or2s1 U27088 ( .DIN1(n34642), .DIN2(n34643), .Q(n34641) );
  and2s1 U27089 ( .DIN1(n33674), .DIN2(n9072), .Q(n34643) );
  and2s1 U27090 ( .DIN1(n33675), .DIN2(n9047), .Q(n34642) );
  or2s1 U27091 ( .DIN1(n34644), .DIN2(n34645), .Q(n34640) );
  and2s1 U27092 ( .DIN1(n33682), .DIN2(n32706), .Q(n34645) );
  hi1s1 U27093 ( .DIN1(n36651), .Q(n32706) );
  and2s1 U27094 ( .DIN1(n34380), .DIN2(n34639), .Q(n34644) );
  hi1s1 U27095 ( .DIN1(n36650), .Q(n34639) );
  or2s1 U27096 ( .DIN1(n34646), .DIN2(n34647), .Q(n9317) );
  or2s1 U27097 ( .DIN1(n34648), .DIN2(n34649), .Q(n34647) );
  and2s1 U27098 ( .DIN1(n34592), .DIN2(n32727), .Q(n34649) );
  hi1s1 U27099 ( .DIN1(n36652), .Q(n32727) );
  and2s1 U27100 ( .DIN1(n34593), .DIN2(n32703), .Q(n34648) );
  and2s1 U27101 ( .DIN1(n34594), .DIN2(n34650), .Q(n34646) );
  or2s1 U27102 ( .DIN1(n34651), .DIN2(n34652), .Q(n9316) );
  or2s1 U27103 ( .DIN1(n34653), .DIN2(n34654), .Q(n34652) );
  and2s1 U27104 ( .DIN1(n33674), .DIN2(n9073), .Q(n34654) );
  and2s1 U27105 ( .DIN1(n33675), .DIN2(n9046), .Q(n34653) );
  or2s1 U27106 ( .DIN1(n34655), .DIN2(n34656), .Q(n34651) );
  and2s1 U27107 ( .DIN1(n33682), .DIN2(n32703), .Q(n34656) );
  hi1s1 U27108 ( .DIN1(n36654), .Q(n32703) );
  and2s1 U27109 ( .DIN1(n34380), .DIN2(n34650), .Q(n34655) );
  hi1s1 U27110 ( .DIN1(n36653), .Q(n34650) );
  or2s1 U27111 ( .DIN1(n34657), .DIN2(n34658), .Q(n9315) );
  or2s1 U27112 ( .DIN1(n34659), .DIN2(n34660), .Q(n34658) );
  and2s1 U27113 ( .DIN1(n34592), .DIN2(n32724), .Q(n34660) );
  hi1s1 U27114 ( .DIN1(n36655), .Q(n32724) );
  and2s1 U27115 ( .DIN1(n34593), .DIN2(n32700), .Q(n34659) );
  and2s1 U27116 ( .DIN1(n34594), .DIN2(n34661), .Q(n34657) );
  or2s1 U27117 ( .DIN1(n34662), .DIN2(n34663), .Q(n9314) );
  or2s1 U27118 ( .DIN1(n34664), .DIN2(n34665), .Q(n34663) );
  and2s1 U27119 ( .DIN1(n33674), .DIN2(n9074), .Q(n34665) );
  and2s1 U27120 ( .DIN1(n33675), .DIN2(n9045), .Q(n34664) );
  or2s1 U27121 ( .DIN1(n34666), .DIN2(n34667), .Q(n34662) );
  and2s1 U27122 ( .DIN1(n33682), .DIN2(n32700), .Q(n34667) );
  hi1s1 U27123 ( .DIN1(n36657), .Q(n32700) );
  and2s1 U27124 ( .DIN1(n34380), .DIN2(n34661), .Q(n34666) );
  hi1s1 U27125 ( .DIN1(n36656), .Q(n34661) );
  or2s1 U27126 ( .DIN1(n34668), .DIN2(n34669), .Q(n9313) );
  or2s1 U27127 ( .DIN1(n34670), .DIN2(n34671), .Q(n34669) );
  and2s1 U27128 ( .DIN1(n34592), .DIN2(n32721), .Q(n34671) );
  hi1s1 U27129 ( .DIN1(n36658), .Q(n32721) );
  and2s1 U27130 ( .DIN1(n34533), .DIN2(n34672), .Q(n34592) );
  and2s1 U27131 ( .DIN1(n34593), .DIN2(n32697), .Q(n34670) );
  and2s1 U27132 ( .DIN1(u0_csc[4]), .DIN2(n34672), .Q(n34593) );
  hi1s1 U27133 ( .DIN1(n34594), .Q(n34672) );
  and2s1 U27134 ( .DIN1(n34594), .DIN2(n34673), .Q(n34668) );
  or2s1 U27135 ( .DIN1(n34674), .DIN2(n34675), .Q(n34594) );
  or2s1 U27136 ( .DIN1(u0_csc[5]), .DIN2(n34676), .Q(n34675) );
  and2s1 U27137 ( .DIN1(n15504), .DIN2(u0_csc[4]), .Q(n34676) );
  and2s1 U27138 ( .DIN1(n15481), .DIN2(n34533), .Q(n34674) );
  hi1s1 U27139 ( .DIN1(u0_csc[4]), .Q(n34533) );
  or2s1 U27140 ( .DIN1(n34677), .DIN2(n34678), .Q(n9312) );
  or2s1 U27141 ( .DIN1(n34679), .DIN2(n34680), .Q(n34678) );
  and2s1 U27142 ( .DIN1(n33674), .DIN2(n9075), .Q(n34680) );
  and2s1 U27143 ( .DIN1(n33675), .DIN2(n9044), .Q(n34679) );
  and2s1 U27144 ( .DIN1(n32614), .DIN2(n34681), .Q(n33675) );
  or2s1 U27145 ( .DIN1(n34682), .DIN2(n34683), .Q(n34677) );
  and2s1 U27146 ( .DIN1(n33682), .DIN2(n32697), .Q(n34683) );
  hi1s1 U27147 ( .DIN1(n36660), .Q(n32697) );
  and2s1 U27148 ( .DIN1(u0_csc[5]), .DIN2(n34684), .Q(n33682) );
  and2s1 U27149 ( .DIN1(n34685), .DIN2(n32614), .Q(n34684) );
  and2s1 U27150 ( .DIN1(n34380), .DIN2(n34673), .Q(n34682) );
  hi1s1 U27151 ( .DIN1(n36659), .Q(n34673) );
  and2s1 U27152 ( .DIN1(n32614), .DIN2(n34686), .Q(n34380) );
  and2s1 U27153 ( .DIN1(n34687), .DIN2(n34685), .Q(n34686) );
  hi1s1 U27154 ( .DIN1(u0_csc[5]), .Q(n34687) );
  hi1s1 U27155 ( .DIN1(n33674), .Q(n32614) );
  or2s1 U27156 ( .DIN1(wb_addr_i[29]), .DIN2(n34688), .Q(n33674) );
  or2s1 U27157 ( .DIN1(wb_addr_i[31]), .DIN2(wb_addr_i[30]), .Q(n34688) );
  or2s1 U27158 ( .DIN1(n34689), .DIN2(n34690), .Q(n9310) );
  or2s1 U27159 ( .DIN1(n34691), .DIN2(n34692), .Q(n34690) );
  and2s1 U27160 ( .DIN1(n34693), .DIN2(wb_addr_i[11]), .Q(n34692) );
  and2s1 U27161 ( .DIN1(n34694), .DIN2(wb_addr_i[12]), .Q(n34691) );
  or2s1 U27162 ( .DIN1(n34695), .DIN2(n34696), .Q(n34689) );
  or2s1 U27163 ( .DIN1(n34697), .DIN2(n34698), .Q(n34696) );
  and2s1 U27164 ( .DIN1(n34699), .DIN2(wb_addr_i[13]), .Q(n34698) );
  and2s1 U27165 ( .DIN1(u1_u0_inc_in[11]), .DIN2(n34700), .Q(n34697) );
  and2s1 U27166 ( .DIN1(n34701), .DIN2(n4581), .Q(n34695) );
  or2s1 U27167 ( .DIN1(n34702), .DIN2(n34703), .Q(n9309) );
  or2s1 U27168 ( .DIN1(n34704), .DIN2(n34705), .Q(n34703) );
  and2s1 U27169 ( .DIN1(wb_addr_i[0]), .DIN2(n34693), .Q(n34705) );
  and2s1 U27170 ( .DIN1(wb_addr_i[1]), .DIN2(n34694), .Q(n34704) );
  or2s1 U27171 ( .DIN1(n34706), .DIN2(n34707), .Q(n34702) );
  or2s1 U27172 ( .DIN1(n34708), .DIN2(n34709), .Q(n34707) );
  and2s1 U27173 ( .DIN1(n34699), .DIN2(wb_addr_i[2]), .Q(n34709) );
  and2s1 U27174 ( .DIN1(n34700), .DIN2(u1_u0_inc_in[0]), .Q(n34708) );
  and2s1 U27175 ( .DIN1(n34701), .DIN2(n4580), .Q(n34706) );
  or2s1 U27176 ( .DIN1(n34710), .DIN2(n34711), .Q(n9308) );
  or2s1 U27177 ( .DIN1(n34712), .DIN2(n34713), .Q(n34711) );
  and2s1 U27178 ( .DIN1(wb_addr_i[1]), .DIN2(n34693), .Q(n34713) );
  and2s1 U27179 ( .DIN1(n34694), .DIN2(wb_addr_i[2]), .Q(n34712) );
  or2s1 U27180 ( .DIN1(n34714), .DIN2(n34715), .Q(n34710) );
  or2s1 U27181 ( .DIN1(n34716), .DIN2(n34717), .Q(n34715) );
  and2s1 U27182 ( .DIN1(n34699), .DIN2(wb_addr_i[3]), .Q(n34717) );
  and2s1 U27183 ( .DIN1(u1_u0_inc_in[1]), .DIN2(n34700), .Q(n34716) );
  and2s1 U27184 ( .DIN1(n34701), .DIN2(n4579), .Q(n34714) );
  or2s1 U27185 ( .DIN1(n34718), .DIN2(n34719), .Q(n9307) );
  or2s1 U27186 ( .DIN1(n34720), .DIN2(n34721), .Q(n34719) );
  and2s1 U27187 ( .DIN1(n34693), .DIN2(wb_addr_i[2]), .Q(n34721) );
  and2s1 U27188 ( .DIN1(n34694), .DIN2(wb_addr_i[3]), .Q(n34720) );
  or2s1 U27189 ( .DIN1(n34722), .DIN2(n34723), .Q(n34718) );
  or2s1 U27190 ( .DIN1(n34724), .DIN2(n34725), .Q(n34723) );
  and2s1 U27191 ( .DIN1(n34699), .DIN2(wb_addr_i[4]), .Q(n34725) );
  and2s1 U27192 ( .DIN1(u1_u0_inc_in[2]), .DIN2(n34700), .Q(n34724) );
  and2s1 U27193 ( .DIN1(n34701), .DIN2(n4578), .Q(n34722) );
  or2s1 U27194 ( .DIN1(n34726), .DIN2(n34727), .Q(n9306) );
  or2s1 U27195 ( .DIN1(n34728), .DIN2(n34729), .Q(n34727) );
  and2s1 U27196 ( .DIN1(n34693), .DIN2(wb_addr_i[3]), .Q(n34729) );
  and2s1 U27197 ( .DIN1(n34694), .DIN2(wb_addr_i[4]), .Q(n34728) );
  or2s1 U27198 ( .DIN1(n34730), .DIN2(n34731), .Q(n34726) );
  or2s1 U27199 ( .DIN1(n34732), .DIN2(n34733), .Q(n34731) );
  and2s1 U27200 ( .DIN1(n34699), .DIN2(wb_addr_i[5]), .Q(n34733) );
  and2s1 U27201 ( .DIN1(u1_u0_inc_in[3]), .DIN2(n34700), .Q(n34732) );
  and2s1 U27202 ( .DIN1(n34701), .DIN2(n4577), .Q(n34730) );
  or2s1 U27203 ( .DIN1(n34734), .DIN2(n34735), .Q(n9305) );
  or2s1 U27204 ( .DIN1(n34736), .DIN2(n34737), .Q(n34735) );
  and2s1 U27205 ( .DIN1(n34693), .DIN2(wb_addr_i[4]), .Q(n34737) );
  and2s1 U27206 ( .DIN1(n34694), .DIN2(wb_addr_i[5]), .Q(n34736) );
  or2s1 U27207 ( .DIN1(n34738), .DIN2(n34739), .Q(n34734) );
  or2s1 U27208 ( .DIN1(n34740), .DIN2(n34741), .Q(n34739) );
  and2s1 U27209 ( .DIN1(n34699), .DIN2(wb_addr_i[6]), .Q(n34741) );
  and2s1 U27210 ( .DIN1(u1_u0_inc_in[4]), .DIN2(n34700), .Q(n34740) );
  and2s1 U27211 ( .DIN1(n34701), .DIN2(n4576), .Q(n34738) );
  or2s1 U27212 ( .DIN1(n34742), .DIN2(n34743), .Q(n9304) );
  or2s1 U27213 ( .DIN1(n34744), .DIN2(n34745), .Q(n34743) );
  and2s1 U27214 ( .DIN1(n34693), .DIN2(wb_addr_i[5]), .Q(n34745) );
  and2s1 U27215 ( .DIN1(n34694), .DIN2(wb_addr_i[6]), .Q(n34744) );
  or2s1 U27216 ( .DIN1(n34746), .DIN2(n34747), .Q(n34742) );
  or2s1 U27217 ( .DIN1(n34748), .DIN2(n34749), .Q(n34747) );
  and2s1 U27218 ( .DIN1(n34699), .DIN2(wb_addr_i[7]), .Q(n34749) );
  and2s1 U27219 ( .DIN1(u1_u0_inc_in[5]), .DIN2(n34700), .Q(n34748) );
  and2s1 U27220 ( .DIN1(n34701), .DIN2(n4575), .Q(n34746) );
  or2s1 U27221 ( .DIN1(n34750), .DIN2(n34751), .Q(n9303) );
  or2s1 U27222 ( .DIN1(n34752), .DIN2(n34753), .Q(n34751) );
  and2s1 U27223 ( .DIN1(n34693), .DIN2(wb_addr_i[6]), .Q(n34753) );
  and2s1 U27224 ( .DIN1(n34694), .DIN2(wb_addr_i[7]), .Q(n34752) );
  or2s1 U27225 ( .DIN1(n34754), .DIN2(n34755), .Q(n34750) );
  or2s1 U27226 ( .DIN1(n34756), .DIN2(n34757), .Q(n34755) );
  and2s1 U27227 ( .DIN1(n34699), .DIN2(wb_addr_i[8]), .Q(n34757) );
  and2s1 U27228 ( .DIN1(u1_u0_inc_in[6]), .DIN2(n34700), .Q(n34756) );
  and2s1 U27229 ( .DIN1(n34701), .DIN2(n4574), .Q(n34754) );
  or2s1 U27230 ( .DIN1(n34758), .DIN2(n34759), .Q(n9302) );
  or2s1 U27231 ( .DIN1(n34760), .DIN2(n34761), .Q(n34759) );
  and2s1 U27232 ( .DIN1(n34693), .DIN2(wb_addr_i[7]), .Q(n34761) );
  and2s1 U27233 ( .DIN1(n34694), .DIN2(wb_addr_i[8]), .Q(n34760) );
  or2s1 U27234 ( .DIN1(n34762), .DIN2(n34763), .Q(n34758) );
  or2s1 U27235 ( .DIN1(n34764), .DIN2(n34765), .Q(n34763) );
  and2s1 U27236 ( .DIN1(n34699), .DIN2(wb_addr_i[9]), .Q(n34765) );
  and2s1 U27237 ( .DIN1(u1_u0_inc_in[7]), .DIN2(n34700), .Q(n34764) );
  and2s1 U27238 ( .DIN1(n34701), .DIN2(n4573), .Q(n34762) );
  or2s1 U27239 ( .DIN1(n34766), .DIN2(n34767), .Q(n9301) );
  or2s1 U27240 ( .DIN1(n34768), .DIN2(n34769), .Q(n34767) );
  and2s1 U27241 ( .DIN1(n34693), .DIN2(wb_addr_i[8]), .Q(n34769) );
  and2s1 U27242 ( .DIN1(n34694), .DIN2(wb_addr_i[9]), .Q(n34768) );
  or2s1 U27243 ( .DIN1(n34770), .DIN2(n34771), .Q(n34766) );
  or2s1 U27244 ( .DIN1(n34772), .DIN2(n34773), .Q(n34771) );
  and2s1 U27245 ( .DIN1(n34699), .DIN2(wb_addr_i[10]), .Q(n34773) );
  and2s1 U27246 ( .DIN1(u1_u0_inc_in[8]), .DIN2(n34700), .Q(n34772) );
  and2s1 U27247 ( .DIN1(n34701), .DIN2(n4572), .Q(n34770) );
  or2s1 U27248 ( .DIN1(n34774), .DIN2(n34775), .Q(n9300) );
  or2s1 U27249 ( .DIN1(n34776), .DIN2(n34777), .Q(n34775) );
  and2s1 U27250 ( .DIN1(n34693), .DIN2(wb_addr_i[9]), .Q(n34777) );
  and2s1 U27251 ( .DIN1(n34694), .DIN2(wb_addr_i[10]), .Q(n34776) );
  or2s1 U27252 ( .DIN1(n34778), .DIN2(n34779), .Q(n34774) );
  or2s1 U27253 ( .DIN1(n34780), .DIN2(n34781), .Q(n34779) );
  and2s1 U27254 ( .DIN1(n34699), .DIN2(wb_addr_i[11]), .Q(n34781) );
  and2s1 U27255 ( .DIN1(u1_u0_inc_in[9]), .DIN2(n34700), .Q(n34780) );
  and2s1 U27256 ( .DIN1(n34701), .DIN2(n4571), .Q(n34778) );
  or2s1 U27257 ( .DIN1(n34782), .DIN2(n34783), .Q(n9299) );
  or2s1 U27258 ( .DIN1(n34784), .DIN2(n34785), .Q(n34783) );
  and2s1 U27259 ( .DIN1(n34693), .DIN2(wb_addr_i[10]), .Q(n34785) );
  and2s1 U27260 ( .DIN1(n34694), .DIN2(wb_addr_i[11]), .Q(n34784) );
  or2s1 U27261 ( .DIN1(n34786), .DIN2(n34787), .Q(n34782) );
  or2s1 U27262 ( .DIN1(n34788), .DIN2(n34789), .Q(n34787) );
  and2s1 U27263 ( .DIN1(n34699), .DIN2(wb_addr_i[12]), .Q(n34789) );
  and2s1 U27264 ( .DIN1(u1_u0_inc_in[10]), .DIN2(n34700), .Q(n34788) );
  and2s1 U27265 ( .DIN1(n34701), .DIN2(n4570), .Q(n34786) );
  or2s1 U27266 ( .DIN1(n34790), .DIN2(n34791), .Q(n9298) );
  or2s1 U27267 ( .DIN1(n34792), .DIN2(n34793), .Q(n34791) );
  and2s1 U27268 ( .DIN1(n34693), .DIN2(wb_addr_i[12]), .Q(n34793) );
  and2s1 U27269 ( .DIN1(n34694), .DIN2(wb_addr_i[13]), .Q(n34792) );
  or2s1 U27270 ( .DIN1(n34794), .DIN2(n34795), .Q(n34790) );
  or2s1 U27271 ( .DIN1(n34796), .DIN2(n34797), .Q(n34795) );
  and2s1 U27272 ( .DIN1(n34699), .DIN2(wb_addr_i[14]), .Q(n34797) );
  and2s1 U27273 ( .DIN1(u1_u0_inc_in[12]), .DIN2(n34700), .Q(n34796) );
  and2s1 U27274 ( .DIN1(\u1_u0_out_r[12] ), .DIN2(n34701), .Q(n34794) );
  or2s1 U27275 ( .DIN1(n34798), .DIN2(n34799), .Q(n9297) );
  or2s1 U27276 ( .DIN1(n34800), .DIN2(n34801), .Q(n34799) );
  and2s1 U27277 ( .DIN1(n34693), .DIN2(wb_addr_i[22]), .Q(n34801) );
  and2s1 U27278 ( .DIN1(n34694), .DIN2(wb_addr_i[23]), .Q(n34800) );
  or2s1 U27279 ( .DIN1(n34802), .DIN2(n34803), .Q(n34798) );
  or2s1 U27280 ( .DIN1(n34804), .DIN2(n34805), .Q(n34803) );
  and2s1 U27281 ( .DIN1(u1_u0_inc_in[22]), .DIN2(n34700), .Q(n34805) );
  and2s1 U27282 ( .DIN1(n34701), .DIN2(n34806), .Q(n34804) );
  or2s1 U27283 ( .DIN1(n34807), .DIN2(n34808), .Q(n34806) );
  and2s1 U27284 ( .DIN1(n34809), .DIN2(n34810), .Q(n34808) );
  and2s1 U27285 ( .DIN1(u1_u0_inc_in[21]), .DIN2(n34811), .Q(n34807) );
  and2s1 U27286 ( .DIN1(n34699), .DIN2(wb_addr_i[24]), .Q(n34802) );
  or2s1 U27287 ( .DIN1(n34812), .DIN2(n34813), .Q(n9296) );
  or2s1 U27288 ( .DIN1(n34814), .DIN2(n34815), .Q(n34813) );
  and2s1 U27289 ( .DIN1(n34693), .DIN2(wb_addr_i[13]), .Q(n34815) );
  and2s1 U27290 ( .DIN1(n34694), .DIN2(wb_addr_i[14]), .Q(n34814) );
  or2s1 U27291 ( .DIN1(n34816), .DIN2(n34817), .Q(n34812) );
  or2s1 U27292 ( .DIN1(n34818), .DIN2(n34819), .Q(n34817) );
  and2s1 U27293 ( .DIN1(u1_u0_inc_in[13]), .DIN2(n34700), .Q(n34819) );
  and2s1 U27294 ( .DIN1(n34820), .DIN2(n34701), .Q(n34818) );
  and2s1 U27295 ( .DIN1(n34821), .DIN2(n34822), .Q(n34820) );
  or2s1 U27296 ( .DIN1(u1_u0_inc_in[12]), .DIN2(\u1_u0_out_r[12] ), .Q(n34821) );
  and2s1 U27297 ( .DIN1(n34699), .DIN2(wb_addr_i[15]), .Q(n34816) );
  or2s1 U27298 ( .DIN1(n34823), .DIN2(n34824), .Q(n9295) );
  or2s1 U27299 ( .DIN1(n34825), .DIN2(n34826), .Q(n34824) );
  and2s1 U27300 ( .DIN1(n34693), .DIN2(wb_addr_i[14]), .Q(n34826) );
  and2s1 U27301 ( .DIN1(n34694), .DIN2(wb_addr_i[15]), .Q(n34825) );
  or2s1 U27302 ( .DIN1(n34827), .DIN2(n34828), .Q(n34823) );
  or2s1 U27303 ( .DIN1(n34829), .DIN2(n34830), .Q(n34828) );
  and2s1 U27304 ( .DIN1(u1_u0_inc_in[14]), .DIN2(n34700), .Q(n34830) );
  and2s1 U27305 ( .DIN1(n34701), .DIN2(n34831), .Q(n34829) );
  or2s1 U27306 ( .DIN1(n34832), .DIN2(n34833), .Q(n34831) );
  and2s1 U27307 ( .DIN1(n34834), .DIN2(n34835), .Q(n34833) );
  and2s1 U27308 ( .DIN1(u1_u0_inc_in[13]), .DIN2(n34822), .Q(n34832) );
  and2s1 U27309 ( .DIN1(n34699), .DIN2(wb_addr_i[16]), .Q(n34827) );
  or2s1 U27310 ( .DIN1(n34836), .DIN2(n34837), .Q(n9294) );
  or2s1 U27311 ( .DIN1(n34838), .DIN2(n34839), .Q(n34837) );
  and2s1 U27312 ( .DIN1(n34693), .DIN2(wb_addr_i[15]), .Q(n34839) );
  and2s1 U27313 ( .DIN1(n34694), .DIN2(wb_addr_i[16]), .Q(n34838) );
  or2s1 U27314 ( .DIN1(n34840), .DIN2(n34841), .Q(n34836) );
  or2s1 U27315 ( .DIN1(n34842), .DIN2(n34843), .Q(n34841) );
  and2s1 U27316 ( .DIN1(u1_u0_inc_in[15]), .DIN2(n34700), .Q(n34843) );
  and2s1 U27317 ( .DIN1(n34701), .DIN2(n34844), .Q(n34842) );
  or2s1 U27318 ( .DIN1(n34845), .DIN2(n34846), .Q(n34844) );
  and2s1 U27319 ( .DIN1(n34847), .DIN2(n34848), .Q(n34846) );
  hi1s1 U27320 ( .DIN1(n34849), .Q(n34847) );
  and2s1 U27321 ( .DIN1(u1_u0_inc_in[14]), .DIN2(n34849), .Q(n34845) );
  and2s1 U27322 ( .DIN1(n34699), .DIN2(wb_addr_i[17]), .Q(n34840) );
  or2s1 U27323 ( .DIN1(n34850), .DIN2(n34851), .Q(n9293) );
  or2s1 U27324 ( .DIN1(n34852), .DIN2(n34853), .Q(n34851) );
  and2s1 U27325 ( .DIN1(n34693), .DIN2(wb_addr_i[16]), .Q(n34853) );
  and2s1 U27326 ( .DIN1(n34694), .DIN2(wb_addr_i[17]), .Q(n34852) );
  or2s1 U27327 ( .DIN1(n34854), .DIN2(n34855), .Q(n34850) );
  or2s1 U27328 ( .DIN1(n34856), .DIN2(n34857), .Q(n34855) );
  and2s1 U27329 ( .DIN1(u1_u0_inc_in[16]), .DIN2(n34700), .Q(n34857) );
  and2s1 U27330 ( .DIN1(n34701), .DIN2(n34858), .Q(n34856) );
  or2s1 U27331 ( .DIN1(n34859), .DIN2(n34860), .Q(n34858) );
  and2s1 U27332 ( .DIN1(n34861), .DIN2(n34862), .Q(n34860) );
  hi1s1 U27333 ( .DIN1(n34863), .Q(n34861) );
  and2s1 U27334 ( .DIN1(u1_u0_inc_in[15]), .DIN2(n34863), .Q(n34859) );
  and2s1 U27335 ( .DIN1(n34699), .DIN2(wb_addr_i[18]), .Q(n34854) );
  or2s1 U27336 ( .DIN1(n34864), .DIN2(n34865), .Q(n9292) );
  or2s1 U27337 ( .DIN1(n34866), .DIN2(n34867), .Q(n34865) );
  and2s1 U27338 ( .DIN1(n34693), .DIN2(wb_addr_i[17]), .Q(n34867) );
  and2s1 U27339 ( .DIN1(n34694), .DIN2(wb_addr_i[18]), .Q(n34866) );
  or2s1 U27340 ( .DIN1(n34868), .DIN2(n34869), .Q(n34864) );
  or2s1 U27341 ( .DIN1(n34870), .DIN2(n34871), .Q(n34869) );
  and2s1 U27342 ( .DIN1(u1_u0_inc_in[17]), .DIN2(n34700), .Q(n34871) );
  and2s1 U27343 ( .DIN1(n34701), .DIN2(n34872), .Q(n34870) );
  or2s1 U27344 ( .DIN1(n34873), .DIN2(n34874), .Q(n34872) );
  and2s1 U27345 ( .DIN1(n34875), .DIN2(n34876), .Q(n34874) );
  hi1s1 U27346 ( .DIN1(n34877), .Q(n34875) );
  and2s1 U27347 ( .DIN1(u1_u0_inc_in[16]), .DIN2(n34877), .Q(n34873) );
  and2s1 U27348 ( .DIN1(n34699), .DIN2(wb_addr_i[19]), .Q(n34868) );
  or2s1 U27349 ( .DIN1(n34878), .DIN2(n34879), .Q(n9291) );
  or2s1 U27350 ( .DIN1(n34880), .DIN2(n34881), .Q(n34879) );
  and2s1 U27351 ( .DIN1(n34693), .DIN2(wb_addr_i[18]), .Q(n34881) );
  and2s1 U27352 ( .DIN1(n34694), .DIN2(wb_addr_i[19]), .Q(n34880) );
  or2s1 U27353 ( .DIN1(n34882), .DIN2(n34883), .Q(n34878) );
  or2s1 U27354 ( .DIN1(n34884), .DIN2(n34885), .Q(n34883) );
  and2s1 U27355 ( .DIN1(u1_u0_inc_in[18]), .DIN2(n34700), .Q(n34885) );
  and2s1 U27356 ( .DIN1(n34701), .DIN2(n34886), .Q(n34884) );
  or2s1 U27357 ( .DIN1(n34887), .DIN2(n34888), .Q(n34886) );
  and2s1 U27358 ( .DIN1(n34889), .DIN2(n34890), .Q(n34888) );
  hi1s1 U27359 ( .DIN1(n34891), .Q(n34889) );
  and2s1 U27360 ( .DIN1(u1_u0_inc_in[17]), .DIN2(n34891), .Q(n34887) );
  and2s1 U27361 ( .DIN1(n34699), .DIN2(wb_addr_i[20]), .Q(n34882) );
  or2s1 U27362 ( .DIN1(n34892), .DIN2(n34893), .Q(n9290) );
  or2s1 U27363 ( .DIN1(n34894), .DIN2(n34895), .Q(n34893) );
  and2s1 U27364 ( .DIN1(n34693), .DIN2(wb_addr_i[19]), .Q(n34895) );
  and2s1 U27365 ( .DIN1(n34694), .DIN2(wb_addr_i[20]), .Q(n34894) );
  or2s1 U27366 ( .DIN1(n34896), .DIN2(n34897), .Q(n34892) );
  or2s1 U27367 ( .DIN1(n34898), .DIN2(n34899), .Q(n34897) );
  and2s1 U27368 ( .DIN1(u1_u0_inc_in[19]), .DIN2(n34700), .Q(n34899) );
  and2s1 U27369 ( .DIN1(n34701), .DIN2(n34900), .Q(n34898) );
  or2s1 U27370 ( .DIN1(n34901), .DIN2(n34902), .Q(n34900) );
  and2s1 U27371 ( .DIN1(n34903), .DIN2(n34904), .Q(n34902) );
  hi1s1 U27372 ( .DIN1(u1_u0_inc_in[18]), .Q(n34904) );
  and2s1 U27373 ( .DIN1(u1_u0_inc_in[18]), .DIN2(n34905), .Q(n34901) );
  and2s1 U27374 ( .DIN1(n34699), .DIN2(wb_addr_i[21]), .Q(n34896) );
  or2s1 U27375 ( .DIN1(n34906), .DIN2(n34907), .Q(n9289) );
  or2s1 U27376 ( .DIN1(n34908), .DIN2(n34909), .Q(n34907) );
  and2s1 U27377 ( .DIN1(n34693), .DIN2(wb_addr_i[20]), .Q(n34909) );
  and2s1 U27378 ( .DIN1(n34694), .DIN2(wb_addr_i[21]), .Q(n34908) );
  or2s1 U27379 ( .DIN1(n34910), .DIN2(n34911), .Q(n34906) );
  or2s1 U27380 ( .DIN1(n34912), .DIN2(n34913), .Q(n34911) );
  and2s1 U27381 ( .DIN1(u1_u0_inc_in[20]), .DIN2(n34700), .Q(n34913) );
  and2s1 U27382 ( .DIN1(n34701), .DIN2(n34914), .Q(n34912) );
  or2s1 U27383 ( .DIN1(n34915), .DIN2(n34916), .Q(n34914) );
  hi1s1 U27384 ( .DIN1(n34917), .Q(n34916) );
  or2s1 U27385 ( .DIN1(n34918), .DIN2(u1_u0_inc_in[19]), .Q(n34917) );
  and2s1 U27386 ( .DIN1(u1_u0_inc_in[19]), .DIN2(n34918), .Q(n34915) );
  hi1s1 U27387 ( .DIN1(n34919), .Q(n34918) );
  and2s1 U27388 ( .DIN1(n34699), .DIN2(wb_addr_i[22]), .Q(n34910) );
  or2s1 U27389 ( .DIN1(n34920), .DIN2(n34921), .Q(n9288) );
  or2s1 U27390 ( .DIN1(n34922), .DIN2(n34923), .Q(n34921) );
  and2s1 U27391 ( .DIN1(n34693), .DIN2(wb_addr_i[21]), .Q(n34923) );
  and2s1 U27392 ( .DIN1(n34694), .DIN2(wb_addr_i[22]), .Q(n34922) );
  or2s1 U27393 ( .DIN1(n34924), .DIN2(n34925), .Q(n34920) );
  or2s1 U27394 ( .DIN1(n34926), .DIN2(n34927), .Q(n34925) );
  and2s1 U27395 ( .DIN1(u1_u0_inc_in[21]), .DIN2(n34700), .Q(n34927) );
  and2s1 U27396 ( .DIN1(n34701), .DIN2(n34928), .Q(n34926) );
  or2s1 U27397 ( .DIN1(n34929), .DIN2(n34930), .Q(n34928) );
  and2s1 U27398 ( .DIN1(n34931), .DIN2(n34932), .Q(n34930) );
  hi1s1 U27399 ( .DIN1(n34933), .Q(n34929) );
  or2s1 U27400 ( .DIN1(n34932), .DIN2(n34931), .Q(n34933) );
  hi1s1 U27401 ( .DIN1(u1_u0_inc_in[20]), .Q(n34932) );
  and2s1 U27402 ( .DIN1(n34699), .DIN2(wb_addr_i[23]), .Q(n34924) );
  or2s1 U27403 ( .DIN1(n34934), .DIN2(n34935), .Q(n9287) );
  or2s1 U27404 ( .DIN1(n34936), .DIN2(n34937), .Q(n34935) );
  and2s1 U27405 ( .DIN1(n34693), .DIN2(wb_addr_i[23]), .Q(n34937) );
  and2s1 U27406 ( .DIN1(n34694), .DIN2(wb_addr_i[24]), .Q(n34936) );
  or2s1 U27407 ( .DIN1(n34938), .DIN2(n34939), .Q(n34934) );
  or2s1 U27408 ( .DIN1(n34940), .DIN2(n34941), .Q(n34939) );
  and2s1 U27409 ( .DIN1(n34700), .DIN2(n34942), .Q(n34941) );
  hi1s1 U27410 ( .DIN1(n34943), .Q(n34700) );
  or2s1 U27411 ( .DIN1(n34944), .DIN2(n34945), .Q(n34943) );
  or2s1 U27412 ( .DIN1(n34701), .DIN2(n34699), .Q(n34945) );
  or2s1 U27413 ( .DIN1(n34693), .DIN2(n34694), .Q(n34944) );
  and2s1 U27414 ( .DIN1(n34946), .DIN2(n34296), .Q(n34694) );
  and2s1 U27415 ( .DIN1(n34946), .DIN2(n34100), .Q(n34693) );
  and2s1 U27416 ( .DIN1(n34701), .DIN2(n34947), .Q(n34940) );
  or2s1 U27417 ( .DIN1(n34948), .DIN2(n34949), .Q(n34947) );
  hi1s1 U27418 ( .DIN1(n34950), .Q(n34949) );
  or2s1 U27419 ( .DIN1(n34951), .DIN2(u1_u0_inc_in[22]), .Q(n34950) );
  and2s1 U27420 ( .DIN1(u1_u0_inc_in[22]), .DIN2(n34951), .Q(n34948) );
  or2s1 U27421 ( .DIN1(n34810), .DIN2(n34811), .Q(n34951) );
  hi1s1 U27422 ( .DIN1(n34809), .Q(n34811) );
  and2s1 U27423 ( .DIN1(n34931), .DIN2(u1_u0_inc_in[20]), .Q(n34809) );
  and2s1 U27424 ( .DIN1(n34919), .DIN2(u1_u0_inc_in[19]), .Q(n34931) );
  and2s1 U27425 ( .DIN1(n34903), .DIN2(u1_u0_inc_in[18]), .Q(n34919) );
  hi1s1 U27426 ( .DIN1(n34905), .Q(n34903) );
  or2s1 U27427 ( .DIN1(n34891), .DIN2(n34890), .Q(n34905) );
  hi1s1 U27428 ( .DIN1(u1_u0_inc_in[17]), .Q(n34890) );
  or2s1 U27429 ( .DIN1(n34877), .DIN2(n34876), .Q(n34891) );
  hi1s1 U27430 ( .DIN1(u1_u0_inc_in[16]), .Q(n34876) );
  or2s1 U27431 ( .DIN1(n34863), .DIN2(n34862), .Q(n34877) );
  hi1s1 U27432 ( .DIN1(u1_u0_inc_in[15]), .Q(n34862) );
  or2s1 U27433 ( .DIN1(n34849), .DIN2(n34848), .Q(n34863) );
  hi1s1 U27434 ( .DIN1(u1_u0_inc_in[14]), .Q(n34848) );
  or2s1 U27435 ( .DIN1(n34822), .DIN2(n34835), .Q(n34849) );
  hi1s1 U27436 ( .DIN1(u1_u0_inc_in[13]), .Q(n34835) );
  hi1s1 U27437 ( .DIN1(n34834), .Q(n34822) );
  and2s1 U27438 ( .DIN1(u1_u0_inc_in[12]), .DIN2(\u1_u0_out_r[12] ), .Q(n34834) );
  hi1s1 U27439 ( .DIN1(u1_u0_inc_in[21]), .Q(n34810) );
  and2s1 U27440 ( .DIN1(n34952), .DIN2(n34953), .Q(n34701) );
  and2s1 U27441 ( .DIN1(n34954), .DIN2(u5_tmr2_done), .Q(n34953) );
  or2s1 U27442 ( .DIN1(n34955), .DIN2(n34956), .Q(n34954) );
  and2s1 U27443 ( .DIN1(n34297), .DIN2(n34957), .Q(n34956) );
  and2s1 U27444 ( .DIN1(n34699), .DIN2(wb_addr_i[25]), .Q(n34938) );
  and2s1 U27445 ( .DIN1(n34958), .DIN2(n34959), .Q(n34699) );
  and2s1 U27446 ( .DIN1(n32850), .DIN2(n34946), .Q(n34959) );
  hi1s1 U27447 ( .DIN1(n34952), .Q(n34946) );
  and2s1 U27448 ( .DIN1(n33495), .DIN2(n32639), .Q(n34952) );
  hi1s1 U27449 ( .DIN1(wb_we_i), .Q(n32639) );
  or2s1 U27450 ( .DIN1(n34960), .DIN2(n34961), .Q(n9286) );
  or2s1 U27451 ( .DIN1(n34962), .DIN2(n34963), .Q(n34961) );
  and2s1 U27452 ( .DIN1(u5_burst_cnt[9]), .DIN2(n33483), .Q(n34963) );
  or2s1 U27453 ( .DIN1(n34964), .DIN2(n34965), .Q(n33483) );
  and2s1 U27454 ( .DIN1(n33479), .DIN2(n34966), .Q(n34964) );
  and2s1 U27455 ( .DIN1(n34967), .DIN2(n33479), .Q(n34962) );
  hi1s1 U27456 ( .DIN1(n34968), .Q(n34967) );
  or2s1 U27457 ( .DIN1(n34966), .DIN2(u5_burst_cnt[9]), .Q(n34968) );
  and2s1 U27458 ( .DIN1(n32870), .DIN2(n9018), .Q(n34960) );
  or2s1 U27459 ( .DIN1(n34969), .DIN2(n34970), .Q(n9285) );
  or2s1 U27460 ( .DIN1(n34971), .DIN2(n34972), .Q(n34970) );
  and2s1 U27461 ( .DIN1(u5_burst_cnt[0]), .DIN2(n34965), .Q(n34972) );
  and2s1 U27462 ( .DIN1(n33479), .DIN2(n34973), .Q(n34971) );
  hi1s1 U27463 ( .DIN1(u5_burst_cnt[0]), .Q(n34973) );
  and2s1 U27464 ( .DIN1(n32870), .DIN2(n9027), .Q(n34969) );
  or2s1 U27465 ( .DIN1(n34974), .DIN2(n34975), .Q(n9284) );
  or2s1 U27466 ( .DIN1(n34976), .DIN2(n34977), .Q(n34975) );
  and2s1 U27467 ( .DIN1(n33479), .DIN2(n34978), .Q(n34977) );
  hi1s1 U27468 ( .DIN1(n34979), .Q(n34978) );
  and2s1 U27469 ( .DIN1(u5_burst_cnt[1]), .DIN2(n34980), .Q(n34976) );
  or2s1 U27470 ( .DIN1(n34981), .DIN2(n34965), .Q(n34980) );
  and2s1 U27471 ( .DIN1(u5_burst_cnt[0]), .DIN2(n33479), .Q(n34981) );
  and2s1 U27472 ( .DIN1(n32870), .DIN2(n9026), .Q(n34974) );
  or2s1 U27473 ( .DIN1(n34982), .DIN2(n34983), .Q(n9283) );
  and2s1 U27474 ( .DIN1(n34984), .DIN2(n34985), .Q(n34983) );
  or2s1 U27475 ( .DIN1(n34986), .DIN2(n34987), .Q(n34984) );
  or2s1 U27476 ( .DIN1(n34111), .DIN2(n34988), .Q(n34987) );
  and2s1 U27477 ( .DIN1(n34989), .DIN2(n34315), .Q(n34988) );
  hi1s1 U27478 ( .DIN1(n34990), .Q(n34989) );
  and2s1 U27479 ( .DIN1(n32870), .DIN2(n9025), .Q(n34986) );
  and2s1 U27480 ( .DIN1(u5_burst_cnt[2]), .DIN2(n34991), .Q(n34982) );
  or2s1 U27481 ( .DIN1(n34992), .DIN2(n34965), .Q(n34991) );
  and2s1 U27482 ( .DIN1(n34979), .DIN2(n34315), .Q(n34992) );
  or2s1 U27483 ( .DIN1(n34993), .DIN2(n34994), .Q(n9282) );
  or2s1 U27484 ( .DIN1(n34995), .DIN2(n34996), .Q(n34994) );
  and2s1 U27485 ( .DIN1(u5_burst_cnt[3]), .DIN2(n34997), .Q(n34996) );
  and2s1 U27486 ( .DIN1(n34998), .DIN2(n33479), .Q(n34995) );
  hi1s1 U27487 ( .DIN1(n34999), .Q(n34998) );
  or2s1 U27488 ( .DIN1(n34990), .DIN2(u5_burst_cnt[3]), .Q(n34999) );
  and2s1 U27489 ( .DIN1(n32870), .DIN2(n9024), .Q(n34993) );
  or2s1 U27490 ( .DIN1(n35000), .DIN2(n35001), .Q(n9281) );
  or2s1 U27491 ( .DIN1(n35002), .DIN2(n35003), .Q(n35001) );
  and2s1 U27492 ( .DIN1(n33479), .DIN2(n35004), .Q(n35003) );
  hi1s1 U27493 ( .DIN1(n35005), .Q(n35004) );
  and2s1 U27494 ( .DIN1(u5_burst_cnt[4]), .DIN2(n35006), .Q(n35002) );
  or2s1 U27495 ( .DIN1(n35007), .DIN2(n34997), .Q(n35006) );
  or2s1 U27496 ( .DIN1(n35008), .DIN2(n34965), .Q(n34997) );
  and2s1 U27497 ( .DIN1(n33479), .DIN2(n34990), .Q(n35008) );
  and2s1 U27498 ( .DIN1(u5_burst_cnt[3]), .DIN2(n33479), .Q(n35007) );
  and2s1 U27499 ( .DIN1(n32870), .DIN2(n9023), .Q(n35000) );
  or2s1 U27500 ( .DIN1(n35009), .DIN2(n35010), .Q(n9280) );
  or2s1 U27501 ( .DIN1(n35011), .DIN2(n35012), .Q(n35010) );
  and2s1 U27502 ( .DIN1(u5_burst_cnt[5]), .DIN2(n35013), .Q(n35012) );
  and2s1 U27503 ( .DIN1(n35014), .DIN2(n33479), .Q(n35011) );
  hi1s1 U27504 ( .DIN1(n35015), .Q(n35014) );
  or2s1 U27505 ( .DIN1(n35005), .DIN2(u5_burst_cnt[5]), .Q(n35015) );
  and2s1 U27506 ( .DIN1(n32870), .DIN2(n9022), .Q(n35009) );
  or2s1 U27507 ( .DIN1(n35016), .DIN2(n35017), .Q(n9279) );
  or2s1 U27508 ( .DIN1(n35018), .DIN2(n35019), .Q(n35017) );
  and2s1 U27509 ( .DIN1(n33479), .DIN2(n35020), .Q(n35019) );
  hi1s1 U27510 ( .DIN1(n35021), .Q(n35020) );
  and2s1 U27511 ( .DIN1(u5_burst_cnt[6]), .DIN2(n35022), .Q(n35018) );
  or2s1 U27512 ( .DIN1(n35023), .DIN2(n35013), .Q(n35022) );
  or2s1 U27513 ( .DIN1(n35024), .DIN2(n34965), .Q(n35013) );
  and2s1 U27514 ( .DIN1(n33479), .DIN2(n35005), .Q(n35024) );
  and2s1 U27515 ( .DIN1(u5_burst_cnt[5]), .DIN2(n33479), .Q(n35023) );
  and2s1 U27516 ( .DIN1(n32870), .DIN2(n9021), .Q(n35016) );
  or2s1 U27517 ( .DIN1(n35025), .DIN2(n35026), .Q(n9278) );
  or2s1 U27518 ( .DIN1(n35027), .DIN2(n35028), .Q(n35026) );
  and2s1 U27519 ( .DIN1(u5_burst_cnt[7]), .DIN2(n35029), .Q(n35028) );
  and2s1 U27520 ( .DIN1(n35030), .DIN2(n33479), .Q(n35027) );
  hi1s1 U27521 ( .DIN1(n35031), .Q(n35030) );
  or2s1 U27522 ( .DIN1(n35021), .DIN2(u5_burst_cnt[7]), .Q(n35031) );
  and2s1 U27523 ( .DIN1(n32870), .DIN2(n9020), .Q(n35025) );
  or2s1 U27524 ( .DIN1(n35032), .DIN2(n35033), .Q(n9277) );
  or2s1 U27525 ( .DIN1(n35034), .DIN2(n35035), .Q(n35033) );
  and2s1 U27526 ( .DIN1(n33479), .DIN2(n35036), .Q(n35035) );
  hi1s1 U27527 ( .DIN1(n34966), .Q(n35036) );
  and2s1 U27528 ( .DIN1(u5_burst_cnt[8]), .DIN2(n35037), .Q(n35034) );
  or2s1 U27529 ( .DIN1(n35038), .DIN2(n35029), .Q(n35037) );
  or2s1 U27530 ( .DIN1(n35039), .DIN2(n34965), .Q(n35029) );
  hi1s1 U27531 ( .DIN1(n34985), .Q(n34965) );
  and2s1 U27532 ( .DIN1(n33479), .DIN2(n35021), .Q(n35039) );
  and2s1 U27533 ( .DIN1(u5_burst_cnt[7]), .DIN2(n33479), .Q(n35038) );
  and2s1 U27534 ( .DIN1(n34985), .DIN2(n35040), .Q(n33479) );
  and2s1 U27535 ( .DIN1(n35041), .DIN2(n34315), .Q(n35040) );
  or2s1 U27536 ( .DIN1(n35042), .DIN2(n35043), .Q(n34985) );
  or2s1 U27537 ( .DIN1(n35044), .DIN2(n35045), .Q(n35043) );
  and2s1 U27538 ( .DIN1(n15502), .DIN2(u5_dv), .Q(n35045) );
  or2s1 U27539 ( .DIN1(n35046), .DIN2(n35047), .Q(u5_dv) );
  and2s1 U27540 ( .DIN1(n35048), .DIN2(n34116), .Q(n35047) );
  and2s1 U27541 ( .DIN1(n34587), .DIN2(n4987), .Q(n35048) );
  hi1s1 U27542 ( .DIN1(n36661), .Q(n34587) );
  and2s1 U27543 ( .DIN1(n35049), .DIN2(n35050), .Q(n35046) );
  and2s1 U27544 ( .DIN1(n35051), .DIN2(n4771), .Q(n35050) );
  and2s1 U27545 ( .DIN1(n4770), .DIN2(n35052), .Q(n35051) );
  and2s1 U27546 ( .DIN1(n32869), .DIN2(u5_wb_cycle), .Q(n35049) );
  and2s1 U27547 ( .DIN1(n35053), .DIN2(n35054), .Q(n35044) );
  or2s1 U27548 ( .DIN1(n33889), .DIN2(n35055), .Q(n35053) );
  or2s1 U27549 ( .DIN1(n33006), .DIN2(n34333), .Q(n35055) );
  or2s1 U27550 ( .DIN1(n34111), .DIN2(n32870), .Q(n35042) );
  and2s1 U27551 ( .DIN1(n32870), .DIN2(n9019), .Q(n35032) );
  or2s1 U27552 ( .DIN1(n35056), .DIN2(n35057), .Q(n9276) );
  or2s1 U27553 ( .DIN1(n35058), .DIN2(n35059), .Q(n35057) );
  and2s1 U27554 ( .DIN1(n35060), .DIN2(n35061), .Q(n35059) );
  or2s1 U27555 ( .DIN1(n35062), .DIN2(n35063), .Q(n35061) );
  or2s1 U27556 ( .DIN1(n35064), .DIN2(n35065), .Q(n35063) );
  and2s1 U27557 ( .DIN1(n35066), .DIN2(n35067), .Q(n35065) );
  and2s1 U27558 ( .DIN1(n35068), .DIN2(n35069), .Q(n35064) );
  and2s1 U27559 ( .DIN1(n35070), .DIN2(n35071), .Q(n35062) );
  and2s1 U27560 ( .DIN1(n35072), .DIN2(n35073), .Q(n35058) );
  or2s1 U27561 ( .DIN1(n35074), .DIN2(n35075), .Q(n35073) );
  and2s1 U27562 ( .DIN1(wb_addr_i[10]), .DIN2(n35076), .Q(n35075) );
  and2s1 U27563 ( .DIN1(n35077), .DIN2(n35078), .Q(n35074) );
  or2s1 U27564 ( .DIN1(n35079), .DIN2(n35080), .Q(n35078) );
  and2s1 U27565 ( .DIN1(n35081), .DIN2(n35082), .Q(n35080) );
  and2s1 U27566 ( .DIN1(n35066), .DIN2(wb_addr_i[11]), .Q(n35079) );
  and2s1 U27567 ( .DIN1(n35083), .DIN2(n35084), .Q(n35056) );
  or2s1 U27568 ( .DIN1(n35085), .DIN2(n35086), .Q(n9275) );
  or2s1 U27569 ( .DIN1(n35087), .DIN2(n35088), .Q(n35086) );
  and2s1 U27570 ( .DIN1(n35072), .DIN2(n35089), .Q(n35088) );
  and2s1 U27571 ( .DIN1(n35060), .DIN2(n35090), .Q(n35087) );
  or2s1 U27572 ( .DIN1(n35091), .DIN2(n35092), .Q(n35090) );
  or2s1 U27573 ( .DIN1(n35093), .DIN2(n35094), .Q(n35092) );
  and2s1 U27574 ( .DIN1(n35095), .DIN2(n35071), .Q(n35094) );
  and2s1 U27575 ( .DIN1(n35070), .DIN2(n35069), .Q(n35093) );
  and2s1 U27576 ( .DIN1(n35066), .DIN2(n35068), .Q(n35091) );
  and2s1 U27577 ( .DIN1(n35083), .DIN2(n35096), .Q(n35085) );
  or2s1 U27578 ( .DIN1(n35097), .DIN2(n35098), .Q(n9274) );
  and2s1 U27579 ( .DIN1(n35083), .DIN2(n35099), .Q(n35098) );
  and2s1 U27580 ( .DIN1(n35100), .DIN2(n35071), .Q(n35097) );
  or2s1 U27581 ( .DIN1(n35101), .DIN2(n35102), .Q(n35100) );
  and2s1 U27582 ( .DIN1(n35060), .DIN2(n35068), .Q(n35102) );
  or2s1 U27583 ( .DIN1(n35103), .DIN2(n35104), .Q(n35068) );
  and2s1 U27584 ( .DIN1(n34957), .DIN2(n35105), .Q(n35103) );
  and2s1 U27585 ( .DIN1(n35072), .DIN2(n35095), .Q(n35101) );
  or2s1 U27586 ( .DIN1(n35106), .DIN2(n35107), .Q(n35095) );
  or2s1 U27587 ( .DIN1(n35108), .DIN2(n35109), .Q(n35107) );
  and2s1 U27588 ( .DIN1(n34100), .DIN2(wb_addr_i[26]), .Q(n35109) );
  and2s1 U27589 ( .DIN1(n34296), .DIN2(wb_addr_i[25]), .Q(n35108) );
  and2s1 U27590 ( .DIN1(wb_addr_i[24]), .DIN2(n32850), .Q(n35106) );
  or2s1 U27591 ( .DIN1(n35110), .DIN2(n35111), .Q(n9273) );
  or2s1 U27592 ( .DIN1(n35112), .DIN2(n35113), .Q(n35111) );
  and2s1 U27593 ( .DIN1(n35060), .DIN2(n35114), .Q(n35113) );
  or2s1 U27594 ( .DIN1(n35115), .DIN2(n35116), .Q(n35114) );
  and2s1 U27595 ( .DIN1(n35067), .DIN2(n35082), .Q(n35115) );
  or2s1 U27596 ( .DIN1(n35117), .DIN2(n35118), .Q(n35067) );
  and2s1 U27597 ( .DIN1(n34957), .DIN2(n35119), .Q(n35117) );
  and2s1 U27598 ( .DIN1(n35072), .DIN2(n35120), .Q(n35112) );
  or2s1 U27599 ( .DIN1(n35121), .DIN2(n35122), .Q(n35120) );
  and2s1 U27600 ( .DIN1(n35070), .DIN2(n35082), .Q(n35122) );
  or2s1 U27601 ( .DIN1(n35123), .DIN2(n35124), .Q(n35070) );
  or2s1 U27602 ( .DIN1(n35125), .DIN2(n35126), .Q(n35124) );
  and2s1 U27603 ( .DIN1(n34100), .DIN2(wb_addr_i[25]), .Q(n35126) );
  and2s1 U27604 ( .DIN1(n34296), .DIN2(wb_addr_i[24]), .Q(n35125) );
  and2s1 U27605 ( .DIN1(wb_addr_i[23]), .DIN2(n32850), .Q(n35123) );
  and2s1 U27606 ( .DIN1(n35127), .DIN2(n35105), .Q(n35121) );
  and2s1 U27607 ( .DIN1(n35083), .DIN2(n35128), .Q(n35110) );
  or2s1 U27608 ( .DIN1(n35129), .DIN2(n35130), .Q(n9272) );
  or2s1 U27609 ( .DIN1(n35131), .DIN2(n35132), .Q(n35130) );
  and2s1 U27610 ( .DIN1(n35060), .DIN2(n35133), .Q(n35132) );
  and2s1 U27611 ( .DIN1(n35072), .DIN2(n35134), .Q(n35131) );
  or2s1 U27612 ( .DIN1(n35135), .DIN2(n35104), .Q(n35134) );
  and2s1 U27613 ( .DIN1(wb_addr_i[22]), .DIN2(n32850), .Q(n35104) );
  and2s1 U27614 ( .DIN1(n34957), .DIN2(n35136), .Q(n35135) );
  or2s1 U27615 ( .DIN1(n35137), .DIN2(n35138), .Q(n35136) );
  and2s1 U27616 ( .DIN1(n35066), .DIN2(n35119), .Q(n35138) );
  and2s1 U27617 ( .DIN1(n35105), .DIN2(n35082), .Q(n35137) );
  or2s1 U27618 ( .DIN1(n35139), .DIN2(n35140), .Q(n35105) );
  and2s1 U27619 ( .DIN1(wb_addr_i[23]), .DIN2(n35141), .Q(n35140) );
  and2s1 U27620 ( .DIN1(n34958), .DIN2(wb_addr_i[24]), .Q(n35139) );
  and2s1 U27621 ( .DIN1(n35083), .DIN2(n35142), .Q(n35129) );
  or2s1 U27622 ( .DIN1(n35143), .DIN2(n35144), .Q(n9271) );
  or2s1 U27623 ( .DIN1(n35145), .DIN2(n35146), .Q(n35144) );
  and2s1 U27624 ( .DIN1(n35060), .DIN2(n35147), .Q(n35146) );
  and2s1 U27625 ( .DIN1(n35072), .DIN2(n35148), .Q(n35145) );
  or2s1 U27626 ( .DIN1(n35118), .DIN2(n35149), .Q(n35148) );
  or2s1 U27627 ( .DIN1(n35116), .DIN2(n35150), .Q(n35149) );
  and2s1 U27628 ( .DIN1(n35151), .DIN2(n35119), .Q(n35150) );
  or2s1 U27629 ( .DIN1(n35152), .DIN2(n35153), .Q(n35119) );
  and2s1 U27630 ( .DIN1(wb_addr_i[22]), .DIN2(n35141), .Q(n35153) );
  and2s1 U27631 ( .DIN1(n34958), .DIN2(wb_addr_i[23]), .Q(n35152) );
  and2s1 U27632 ( .DIN1(n35154), .DIN2(n35127), .Q(n35116) );
  and2s1 U27633 ( .DIN1(wb_addr_i[21]), .DIN2(n32850), .Q(n35118) );
  and2s1 U27634 ( .DIN1(n35083), .DIN2(n35155), .Q(n35143) );
  or2s1 U27635 ( .DIN1(n35156), .DIN2(n35157), .Q(n9270) );
  or2s1 U27636 ( .DIN1(n35158), .DIN2(n35159), .Q(n35157) );
  and2s1 U27637 ( .DIN1(n35060), .DIN2(n35160), .Q(n35159) );
  and2s1 U27638 ( .DIN1(n35072), .DIN2(n35133), .Q(n35158) );
  or2s1 U27639 ( .DIN1(n35161), .DIN2(n35162), .Q(n35133) );
  or2s1 U27640 ( .DIN1(n35163), .DIN2(n35164), .Q(n35162) );
  and2s1 U27641 ( .DIN1(n35151), .DIN2(n35154), .Q(n35164) );
  or2s1 U27642 ( .DIN1(n35165), .DIN2(n35166), .Q(n35154) );
  and2s1 U27643 ( .DIN1(wb_addr_i[21]), .DIN2(n35141), .Q(n35166) );
  and2s1 U27644 ( .DIN1(n34958), .DIN2(wb_addr_i[22]), .Q(n35165) );
  and2s1 U27645 ( .DIN1(n35167), .DIN2(wb_addr_i[21]), .Q(n35163) );
  and2s1 U27646 ( .DIN1(wb_addr_i[20]), .DIN2(n35076), .Q(n35161) );
  and2s1 U27647 ( .DIN1(n35083), .DIN2(n35168), .Q(n35156) );
  or2s1 U27648 ( .DIN1(n35169), .DIN2(n35170), .Q(n9269) );
  or2s1 U27649 ( .DIN1(n35171), .DIN2(n35172), .Q(n35170) );
  and2s1 U27650 ( .DIN1(n35060), .DIN2(n35173), .Q(n35172) );
  and2s1 U27651 ( .DIN1(n35072), .DIN2(n35147), .Q(n35171) );
  or2s1 U27652 ( .DIN1(n35174), .DIN2(n35175), .Q(n35147) );
  or2s1 U27653 ( .DIN1(n35176), .DIN2(n35177), .Q(n35175) );
  and2s1 U27654 ( .DIN1(wb_addr_i[20]), .DIN2(n35178), .Q(n35177) );
  and2s1 U27655 ( .DIN1(n35179), .DIN2(wb_addr_i[21]), .Q(n35176) );
  and2s1 U27656 ( .DIN1(wb_addr_i[19]), .DIN2(n35076), .Q(n35174) );
  and2s1 U27657 ( .DIN1(n35083), .DIN2(n35180), .Q(n35169) );
  or2s1 U27658 ( .DIN1(n35181), .DIN2(n35182), .Q(n9268) );
  or2s1 U27659 ( .DIN1(n35183), .DIN2(n35184), .Q(n35182) );
  and2s1 U27660 ( .DIN1(n35060), .DIN2(n35185), .Q(n35184) );
  and2s1 U27661 ( .DIN1(n35072), .DIN2(n35160), .Q(n35183) );
  or2s1 U27662 ( .DIN1(n35186), .DIN2(n35187), .Q(n35160) );
  or2s1 U27663 ( .DIN1(n35188), .DIN2(n35189), .Q(n35187) );
  and2s1 U27664 ( .DIN1(wb_addr_i[19]), .DIN2(n35178), .Q(n35189) );
  and2s1 U27665 ( .DIN1(n35179), .DIN2(wb_addr_i[20]), .Q(n35188) );
  and2s1 U27666 ( .DIN1(wb_addr_i[18]), .DIN2(n35076), .Q(n35186) );
  and2s1 U27667 ( .DIN1(n35083), .DIN2(n35190), .Q(n35181) );
  or2s1 U27668 ( .DIN1(n35191), .DIN2(n35192), .Q(n9267) );
  or2s1 U27669 ( .DIN1(n35193), .DIN2(n35194), .Q(n35192) );
  and2s1 U27670 ( .DIN1(n35060), .DIN2(n35195), .Q(n35194) );
  and2s1 U27671 ( .DIN1(n35072), .DIN2(n35173), .Q(n35193) );
  or2s1 U27672 ( .DIN1(n35196), .DIN2(n35197), .Q(n35173) );
  or2s1 U27673 ( .DIN1(n35198), .DIN2(n35199), .Q(n35197) );
  and2s1 U27674 ( .DIN1(wb_addr_i[18]), .DIN2(n35178), .Q(n35199) );
  and2s1 U27675 ( .DIN1(n35179), .DIN2(wb_addr_i[19]), .Q(n35198) );
  and2s1 U27676 ( .DIN1(wb_addr_i[17]), .DIN2(n35076), .Q(n35196) );
  and2s1 U27677 ( .DIN1(n35083), .DIN2(n35200), .Q(n35191) );
  or2s1 U27678 ( .DIN1(n35201), .DIN2(n35202), .Q(n9266) );
  or2s1 U27679 ( .DIN1(n35203), .DIN2(n35204), .Q(n35202) );
  and2s1 U27680 ( .DIN1(n35060), .DIN2(n35205), .Q(n35204) );
  and2s1 U27681 ( .DIN1(n35072), .DIN2(n35185), .Q(n35203) );
  or2s1 U27682 ( .DIN1(n35206), .DIN2(n35207), .Q(n35185) );
  or2s1 U27683 ( .DIN1(n35208), .DIN2(n35209), .Q(n35207) );
  and2s1 U27684 ( .DIN1(wb_addr_i[17]), .DIN2(n35178), .Q(n35209) );
  and2s1 U27685 ( .DIN1(n35179), .DIN2(wb_addr_i[18]), .Q(n35208) );
  and2s1 U27686 ( .DIN1(wb_addr_i[16]), .DIN2(n35076), .Q(n35206) );
  and2s1 U27687 ( .DIN1(n35083), .DIN2(n35210), .Q(n35201) );
  or2s1 U27688 ( .DIN1(n35211), .DIN2(n35212), .Q(n9265) );
  or2s1 U27689 ( .DIN1(n35213), .DIN2(n35214), .Q(n35212) );
  and2s1 U27690 ( .DIN1(n35060), .DIN2(n35215), .Q(n35214) );
  and2s1 U27691 ( .DIN1(n35072), .DIN2(n35195), .Q(n35213) );
  or2s1 U27692 ( .DIN1(n35216), .DIN2(n35217), .Q(n35195) );
  or2s1 U27693 ( .DIN1(n35218), .DIN2(n35219), .Q(n35217) );
  and2s1 U27694 ( .DIN1(wb_addr_i[16]), .DIN2(n35178), .Q(n35219) );
  and2s1 U27695 ( .DIN1(n35179), .DIN2(wb_addr_i[17]), .Q(n35218) );
  and2s1 U27696 ( .DIN1(wb_addr_i[15]), .DIN2(n35076), .Q(n35216) );
  and2s1 U27697 ( .DIN1(n35083), .DIN2(n35220), .Q(n35211) );
  or2s1 U27698 ( .DIN1(n35221), .DIN2(n35222), .Q(n9264) );
  or2s1 U27699 ( .DIN1(n35223), .DIN2(n35224), .Q(n35222) );
  and2s1 U27700 ( .DIN1(n35060), .DIN2(n35225), .Q(n35224) );
  and2s1 U27701 ( .DIN1(n35072), .DIN2(n35205), .Q(n35223) );
  or2s1 U27702 ( .DIN1(n35226), .DIN2(n35227), .Q(n35205) );
  or2s1 U27703 ( .DIN1(n35228), .DIN2(n35229), .Q(n35227) );
  and2s1 U27704 ( .DIN1(wb_addr_i[15]), .DIN2(n35178), .Q(n35229) );
  and2s1 U27705 ( .DIN1(n35179), .DIN2(wb_addr_i[16]), .Q(n35228) );
  and2s1 U27706 ( .DIN1(wb_addr_i[14]), .DIN2(n35076), .Q(n35226) );
  and2s1 U27707 ( .DIN1(n35083), .DIN2(n35230), .Q(n35221) );
  or2s1 U27708 ( .DIN1(n35231), .DIN2(n35232), .Q(n9263) );
  or2s1 U27709 ( .DIN1(n35233), .DIN2(n35234), .Q(n35232) );
  and2s1 U27710 ( .DIN1(n35060), .DIN2(n35089), .Q(n35234) );
  or2s1 U27711 ( .DIN1(n35235), .DIN2(n35236), .Q(n35089) );
  or2s1 U27712 ( .DIN1(n35237), .DIN2(n35238), .Q(n35236) );
  and2s1 U27713 ( .DIN1(wb_addr_i[11]), .DIN2(n32850), .Q(n35238) );
  and2s1 U27714 ( .DIN1(n35179), .DIN2(wb_addr_i[13]), .Q(n35237) );
  or2s1 U27715 ( .DIN1(n35239), .DIN2(n35240), .Q(n35235) );
  and2s1 U27716 ( .DIN1(n35127), .DIN2(n35081), .Q(n35240) );
  and2s1 U27717 ( .DIN1(n34957), .DIN2(n35066), .Q(n35127) );
  and2s1 U27718 ( .DIN1(n35241), .DIN2(n34296), .Q(n35239) );
  and2s1 U27719 ( .DIN1(wb_addr_i[12]), .DIN2(n35082), .Q(n35241) );
  and2s1 U27720 ( .DIN1(n35072), .DIN2(n35215), .Q(n35233) );
  or2s1 U27721 ( .DIN1(n35242), .DIN2(n35243), .Q(n35215) );
  or2s1 U27722 ( .DIN1(n35244), .DIN2(n35245), .Q(n35243) );
  and2s1 U27723 ( .DIN1(wb_addr_i[14]), .DIN2(n35178), .Q(n35245) );
  and2s1 U27724 ( .DIN1(n35179), .DIN2(wb_addr_i[15]), .Q(n35244) );
  and2s1 U27725 ( .DIN1(wb_addr_i[13]), .DIN2(n35076), .Q(n35242) );
  and2s1 U27726 ( .DIN1(n35083), .DIN2(n35246), .Q(n35231) );
  or2s1 U27727 ( .DIN1(n35247), .DIN2(n35248), .Q(n9262) );
  or2s1 U27728 ( .DIN1(n35249), .DIN2(n35250), .Q(n35248) );
  and2s1 U27729 ( .DIN1(n35072), .DIN2(n35225), .Q(n35250) );
  or2s1 U27730 ( .DIN1(n35251), .DIN2(n35252), .Q(n35225) );
  or2s1 U27731 ( .DIN1(n35253), .DIN2(n35254), .Q(n35252) );
  and2s1 U27732 ( .DIN1(wb_addr_i[13]), .DIN2(n35178), .Q(n35254) );
  or2s1 U27733 ( .DIN1(n35255), .DIN2(n35167), .Q(n35178) );
  and2s1 U27734 ( .DIN1(n34296), .DIN2(n35082), .Q(n35255) );
  and2s1 U27735 ( .DIN1(n35179), .DIN2(wb_addr_i[14]), .Q(n35253) );
  and2s1 U27736 ( .DIN1(n35082), .DIN2(n34100), .Q(n35179) );
  and2s1 U27737 ( .DIN1(wb_addr_i[12]), .DIN2(n35076), .Q(n35251) );
  or2s1 U27738 ( .DIN1(n35256), .DIN2(n32850), .Q(n35076) );
  and2s1 U27739 ( .DIN1(n35066), .DIN2(n35141), .Q(n35256) );
  and2s1 U27740 ( .DIN1(n35257), .DIN2(n35258), .Q(n35072) );
  hi1s1 U27741 ( .DIN1(n35259), .Q(n35257) );
  and2s1 U27742 ( .DIN1(n35060), .DIN2(n35260), .Q(n35249) );
  or2s1 U27743 ( .DIN1(n35261), .DIN2(n35262), .Q(n35260) );
  and2s1 U27744 ( .DIN1(wb_addr_i[10]), .DIN2(n32850), .Q(n35262) );
  and2s1 U27745 ( .DIN1(n34957), .DIN2(n35263), .Q(n35261) );
  or2s1 U27746 ( .DIN1(n35264), .DIN2(n35265), .Q(n35263) );
  or2s1 U27747 ( .DIN1(n35266), .DIN2(n35267), .Q(n35265) );
  and2s1 U27748 ( .DIN1(n35268), .DIN2(n35269), .Q(n35267) );
  or2s1 U27749 ( .DIN1(n35270), .DIN2(n35271), .Q(n35269) );
  and2s1 U27750 ( .DIN1(n35066), .DIN2(wb_addr_i[10]), .Q(n35271) );
  and2s1 U27751 ( .DIN1(wb_addr_i[12]), .DIN2(n35069), .Q(n35270) );
  hi1s1 U27752 ( .DIN1(n35272), .Q(n35268) );
  and2s1 U27753 ( .DIN1(n35273), .DIN2(n35272), .Q(n35266) );
  and2s1 U27754 ( .DIN1(n35274), .DIN2(n35275), .Q(n35272) );
  or2s1 U27755 ( .DIN1(n35069), .DIN2(n34958), .Q(n35275) );
  or2s1 U27756 ( .DIN1(n35141), .DIN2(n35276), .Q(n35274) );
  and2s1 U27757 ( .DIN1(n35277), .DIN2(wb_addr_i[11]), .Q(n35273) );
  and2s1 U27758 ( .DIN1(n35081), .DIN2(n35071), .Q(n35264) );
  or2s1 U27759 ( .DIN1(n35278), .DIN2(n35279), .Q(n35081) );
  and2s1 U27760 ( .DIN1(wb_addr_i[11]), .DIN2(n35141), .Q(n35279) );
  and2s1 U27761 ( .DIN1(n34958), .DIN2(wb_addr_i[12]), .Q(n35278) );
  and2s1 U27762 ( .DIN1(n35259), .DIN2(n35258), .Q(n35060) );
  hi1s1 U27763 ( .DIN1(n35083), .Q(n35258) );
  or2s1 U27764 ( .DIN1(n35280), .DIN2(n35281), .Q(n35259) );
  and2s1 U27765 ( .DIN1(u0_sp_csc_9), .DIN2(n35282), .Q(n35281) );
  and2s1 U27766 ( .DIN1(u0_csc_9), .DIN2(n35283), .Q(n35280) );
  and2s1 U27767 ( .DIN1(n35083), .DIN2(n35284), .Q(n35247) );
  or2s1 U27768 ( .DIN1(n33495), .DIN2(n35285), .Q(n35083) );
  hi1s1 U27769 ( .DIN1(u5_cs_le), .Q(n33495) );
  or2s1 U27770 ( .DIN1(n35286), .DIN2(n35287), .Q(n9261) );
  or2s1 U27771 ( .DIN1(n35288), .DIN2(n35289), .Q(n35287) );
  and2s1 U27772 ( .DIN1(n34075), .DIN2(u0_csc1[3]), .Q(n35289) );
  and2s1 U27773 ( .DIN1(n34076), .DIN2(u0_csc0[3]), .Q(n35288) );
  and2s1 U27774 ( .DIN1(u0_sp_csc[3]), .DIN2(n33641), .Q(n35286) );
  or2s1 U27775 ( .DIN1(n35290), .DIN2(n35291), .Q(n9260) );
  or2s1 U27776 ( .DIN1(n35292), .DIN2(n35293), .Q(n35291) );
  and2s1 U27777 ( .DIN1(n34075), .DIN2(u0_csc1[2]), .Q(n35293) );
  and2s1 U27778 ( .DIN1(n34076), .DIN2(u0_csc0[2]), .Q(n35292) );
  and2s1 U27779 ( .DIN1(u0_sp_csc[2]), .DIN2(n33641), .Q(n35290) );
  or2s1 U27780 ( .DIN1(n35294), .DIN2(n35295), .Q(n9259) );
  or2s1 U27781 ( .DIN1(n35296), .DIN2(n35297), .Q(n35295) );
  and2s1 U27782 ( .DIN1(n34075), .DIN2(n32426), .Q(n35297) );
  and2s1 U27783 ( .DIN1(u0_spec_req_cs[1]), .DIN2(n35298), .Q(n34075) );
  and2s1 U27784 ( .DIN1(n33952), .DIN2(n33743), .Q(n35298) );
  and2s1 U27785 ( .DIN1(n34076), .DIN2(n32750), .Q(n35296) );
  and2s1 U27786 ( .DIN1(n33743), .DIN2(u0_spec_req_cs[0]), .Q(n34076) );
  and2s1 U27787 ( .DIN1(u0_sp_csc[1]), .DIN2(n33641), .Q(n35294) );
  hi1s1 U27788 ( .DIN1(n33743), .Q(n33641) );
  and2s1 U27789 ( .DIN1(n9533), .DIN2(n32625), .Q(n33743) );
  or2s1 U27790 ( .DIN1(n35299), .DIN2(n35300), .Q(n9533) );
  or2s1 U27791 ( .DIN1(n35301), .DIN2(n35302), .Q(n35300) );
  or2s1 U27792 ( .DIN1(n35303), .DIN2(n35304), .Q(n35302) );
  and2s1 U27793 ( .DIN1(u5_wb_stb_first), .DIN2(n32870), .Q(n35304) );
  and2s1 U27794 ( .DIN1(u5_wb_cycle), .DIN2(n35305), .Q(n35303) );
  or2s1 U27795 ( .DIN1(n35306), .DIN2(n35307), .Q(n35305) );
  or2s1 U27796 ( .DIN1(n33894), .DIN2(n33896), .Q(n35307) );
  and2s1 U27797 ( .DIN1(n34560), .DIN2(u5_tmr2_done), .Q(n33894) );
  and2s1 U27798 ( .DIN1(n34545), .DIN2(u5_tmr_done), .Q(n35306) );
  or2s1 U27799 ( .DIN1(n32865), .DIN2(n34324), .Q(n35301) );
  or2s1 U27800 ( .DIN1(n35308), .DIN2(n35309), .Q(n35299) );
  or2s1 U27801 ( .DIN1(n34243), .DIN2(n34263), .Q(n35309) );
  or2s1 U27802 ( .DIN1(n34241), .DIN2(n35310), .Q(n35308) );
  or2s1 U27803 ( .DIN1(n34320), .DIN2(n34280), .Q(n35310) );
  hi1s1 U27804 ( .DIN1(n35311), .Q(n34280) );
  or2s1 U27805 ( .DIN1(n34580), .DIN2(n35312), .Q(n35311) );
  or2s1 U27806 ( .DIN1(n34315), .DIN2(n35313), .Q(n35312) );
  and2s1 U27807 ( .DIN1(n35314), .DIN2(n35315), .Q(n34320) );
  hi1s1 U27808 ( .DIN1(n35316), .Q(n35315) );
  or2s1 U27809 ( .DIN1(n35313), .DIN2(n34579), .Q(n35316) );
  or2s1 U27810 ( .DIN1(n15515), .DIN2(u5_wb_cycle), .Q(n34579) );
  and2s1 U27811 ( .DIN1(n34580), .DIN2(n32870), .Q(n35314) );
  or2s1 U27812 ( .DIN1(n33919), .DIN2(n4990), .Q(n34580) );
  and2s1 U27813 ( .DIN1(u0_init_req), .DIN2(n35317), .Q(n34241) );
  hi1s1 U27814 ( .DIN1(n35318), .Q(n35317) );
  or2s1 U27815 ( .DIN1(u4_rfr_req), .DIN2(n34315), .Q(n35318) );
  hi1s1 U27816 ( .DIN1(n35319), .Q(n9258) );
  or2s1 U27817 ( .DIN1(n33924), .DIN2(n15494), .Q(n35319) );
  hi1s1 U27818 ( .DIN1(n35320), .Q(n9257) );
  or2s1 U27819 ( .DIN1(n33924), .DIN2(n15493), .Q(n35320) );
  hi1s1 U27820 ( .DIN1(n35321), .Q(n9256) );
  or2s1 U27821 ( .DIN1(n33924), .DIN2(n15492), .Q(n35321) );
  hi1s1 U27822 ( .DIN1(n35322), .Q(n9255) );
  or2s1 U27823 ( .DIN1(n33924), .DIN2(n15491), .Q(n35322) );
  hi1s1 U27824 ( .DIN1(n35323), .Q(n9254) );
  or2s1 U27825 ( .DIN1(n33924), .DIN2(n15490), .Q(n35323) );
  hi1s1 U27826 ( .DIN1(n35324), .Q(n9253) );
  or2s1 U27827 ( .DIN1(n33924), .DIN2(n15489), .Q(n35324) );
  hi1s1 U27828 ( .DIN1(n15511), .Q(n33924) );
  or2s1 U27829 ( .DIN1(n35325), .DIN2(n35326), .Q(n9252) );
  and2s1 U27830 ( .DIN1(n34315), .DIN2(n35054), .Q(n35326) );
  and2s1 U27831 ( .DIN1(n33035), .DIN2(n35327), .Q(n35325) );
  and2s1 U27832 ( .DIN1(wb_stb_i), .DIN2(wb_we_i), .Q(n33035) );
  or2s1 U27833 ( .DIN1(n35328), .DIN2(n35329), .Q(n9251) );
  and2s1 U27834 ( .DIN1(n35330), .DIN2(n35331), .Q(n35329) );
  and2s1 U27835 ( .DIN1(n35332), .DIN2(wb_addr_i[2]), .Q(n35328) );
  or2s1 U27836 ( .DIN1(n35333), .DIN2(n35334), .Q(n9250) );
  and2s1 U27837 ( .DIN1(n35330), .DIN2(n35335), .Q(n35334) );
  and2s1 U27838 ( .DIN1(n35332), .DIN2(wb_addr_i[3]), .Q(n35333) );
  or2s1 U27839 ( .DIN1(n35336), .DIN2(n35337), .Q(n9249) );
  and2s1 U27840 ( .DIN1(n35330), .DIN2(n35338), .Q(n35337) );
  and2s1 U27841 ( .DIN1(n35332), .DIN2(wb_addr_i[4]), .Q(n35336) );
  or2s1 U27842 ( .DIN1(n35339), .DIN2(n35340), .Q(n9248) );
  and2s1 U27843 ( .DIN1(n35330), .DIN2(n35341), .Q(n35340) );
  and2s1 U27844 ( .DIN1(n35332), .DIN2(wb_addr_i[5]), .Q(n35339) );
  or2s1 U27845 ( .DIN1(n35342), .DIN2(n35343), .Q(n9247) );
  and2s1 U27846 ( .DIN1(n35330), .DIN2(n35344), .Q(n35343) );
  and2s1 U27847 ( .DIN1(n35332), .DIN2(wb_addr_i[6]), .Q(n35342) );
  or2s1 U27848 ( .DIN1(n35345), .DIN2(n35346), .Q(n9246) );
  and2s1 U27849 ( .DIN1(n35330), .DIN2(n35347), .Q(n35346) );
  and2s1 U27850 ( .DIN1(n35332), .DIN2(wb_addr_i[7]), .Q(n35345) );
  or2s1 U27851 ( .DIN1(n35348), .DIN2(n35349), .Q(n9245) );
  and2s1 U27852 ( .DIN1(n35330), .DIN2(n35350), .Q(n35349) );
  and2s1 U27853 ( .DIN1(n35332), .DIN2(wb_addr_i[8]), .Q(n35348) );
  or2s1 U27854 ( .DIN1(n35351), .DIN2(n35352), .Q(n9244) );
  and2s1 U27855 ( .DIN1(n35330), .DIN2(n35353), .Q(n35352) );
  and2s1 U27856 ( .DIN1(n35332), .DIN2(wb_addr_i[9]), .Q(n35351) );
  or2s1 U27857 ( .DIN1(n35354), .DIN2(n35355), .Q(n9243) );
  and2s1 U27858 ( .DIN1(n35330), .DIN2(n35356), .Q(n35355) );
  and2s1 U27859 ( .DIN1(n35357), .DIN2(n35332), .Q(n35354) );
  and2s1 U27860 ( .DIN1(wb_addr_i[10]), .DIN2(n35358), .Q(n35357) );
  or2s1 U27861 ( .DIN1(n35359), .DIN2(n34100), .Q(n35358) );
  and2s1 U27862 ( .DIN1(n35360), .DIN2(n34957), .Q(n35359) );
  or2s1 U27863 ( .DIN1(n35361), .DIN2(n35362), .Q(n9242) );
  and2s1 U27864 ( .DIN1(n35330), .DIN2(n35363), .Q(n35362) );
  and2s1 U27865 ( .DIN1(n35364), .DIN2(n5504), .Q(n35361) );
  and2s1 U27866 ( .DIN1(n35332), .DIN2(wb_addr_i[11]), .Q(n35364) );
  hi1s1 U27867 ( .DIN1(n35330), .Q(n35332) );
  or2s1 U27868 ( .DIN1(n35365), .DIN2(n35366), .Q(n35330) );
  or2s1 U27869 ( .DIN1(n35367), .DIN2(n35368), .Q(n35366) );
  and2s1 U27870 ( .DIN1(n15502), .DIN2(n32540), .Q(n35368) );
  hi1s1 U27871 ( .DIN1(wb_stb_i), .Q(n32540) );
  hi1s1 U27872 ( .DIN1(n35369), .Q(n35367) );
  or2s1 U27873 ( .DIN1(n15482), .DIN2(n15502), .Q(n35369) );
  or2s1 U27874 ( .DIN1(n35370), .DIN2(n35371), .Q(n35365) );
  and2s1 U27875 ( .DIN1(n35141), .DIN2(n35372), .Q(n35370) );
  or2s1 U27876 ( .DIN1(n35373), .DIN2(n35374), .Q(n9241) );
  or2s1 U27877 ( .DIN1(n35375), .DIN2(n35376), .Q(n35374) );
  and2s1 U27878 ( .DIN1(n33859), .DIN2(n35377), .Q(n35376) );
  and2s1 U27879 ( .DIN1(n33862), .DIN2(n35378), .Q(n35375) );
  or2s1 U27880 ( .DIN1(n35379), .DIN2(n35380), .Q(n35378) );
  hi1s1 U27881 ( .DIN1(n33863), .Q(n35380) );
  and2s1 U27882 ( .DIN1(u5_timer2[7]), .DIN2(n35381), .Q(n35379) );
  and2s1 U27883 ( .DIN1(n35382), .DIN2(n33865), .Q(n35373) );
  or2s1 U27884 ( .DIN1(n35383), .DIN2(n35384), .Q(n9240) );
  or2s1 U27885 ( .DIN1(n33865), .DIN2(n35385), .Q(n35384) );
  or2s1 U27886 ( .DIN1(n35386), .DIN2(n35387), .Q(n35385) );
  and2s1 U27887 ( .DIN1(n35388), .DIN2(n35389), .Q(n35387) );
  and2s1 U27888 ( .DIN1(n33859), .DIN2(n35390), .Q(n35386) );
  or2s1 U27889 ( .DIN1(n35391), .DIN2(n35392), .Q(n35383) );
  or2s1 U27890 ( .DIN1(n35393), .DIN2(n35394), .Q(n35392) );
  hi1s1 U27891 ( .DIN1(n35395), .Q(n35394) );
  or2s1 U27892 ( .DIN1(n35396), .DIN2(u5_timer2[0]), .Q(n35395) );
  and2s1 U27893 ( .DIN1(n35397), .DIN2(n35398), .Q(n35391) );
  or2s1 U27894 ( .DIN1(n35399), .DIN2(n35400), .Q(n9239) );
  or2s1 U27895 ( .DIN1(n35401), .DIN2(n35402), .Q(n35400) );
  or2s1 U27896 ( .DIN1(n35403), .DIN2(n35404), .Q(n35402) );
  and2s1 U27897 ( .DIN1(n35388), .DIN2(n32886), .Q(n35404) );
  and2s1 U27898 ( .DIN1(n35393), .DIN2(n35405), .Q(n35403) );
  and2s1 U27899 ( .DIN1(n35406), .DIN2(n33865), .Q(n35401) );
  or2s1 U27900 ( .DIN1(n35407), .DIN2(n35408), .Q(n35399) );
  or2s1 U27901 ( .DIN1(n35409), .DIN2(n35410), .Q(n35408) );
  and2s1 U27902 ( .DIN1(n33859), .DIN2(n35411), .Q(n35410) );
  and2s1 U27903 ( .DIN1(n35412), .DIN2(n35390), .Q(n35409) );
  or2s1 U27904 ( .DIN1(n35413), .DIN2(n35414), .Q(n35407) );
  and2s1 U27905 ( .DIN1(n35398), .DIN2(n32897), .Q(n35414) );
  or2s1 U27906 ( .DIN1(n35415), .DIN2(n35416), .Q(n32897) );
  or2s1 U27907 ( .DIN1(n35417), .DIN2(n35418), .Q(n35416) );
  and2s1 U27908 ( .DIN1(u0_sp_tms[13]), .DIN2(n35282), .Q(n35418) );
  and2s1 U27909 ( .DIN1(u0_tms[13]), .DIN2(n35283), .Q(n35417) );
  and2s1 U27910 ( .DIN1(n33862), .DIN2(n35419), .Q(n35413) );
  or2s1 U27911 ( .DIN1(n35420), .DIN2(n35421), .Q(n35419) );
  hi1s1 U27912 ( .DIN1(n35422), .Q(n35421) );
  and2s1 U27913 ( .DIN1(u5_timer2[1]), .DIN2(u5_timer2[0]), .Q(n35420) );
  or2s1 U27914 ( .DIN1(n35423), .DIN2(n35424), .Q(n9238) );
  or2s1 U27915 ( .DIN1(n35425), .DIN2(n35426), .Q(n35424) );
  or2s1 U27916 ( .DIN1(n35427), .DIN2(n35428), .Q(n35426) );
  and2s1 U27917 ( .DIN1(n32879), .DIN2(n33865), .Q(n35427) );
  or2s1 U27918 ( .DIN1(n35429), .DIN2(n35430), .Q(n35425) );
  and2s1 U27919 ( .DIN1(n35388), .DIN2(n35431), .Q(n35430) );
  and2s1 U27920 ( .DIN1(n33859), .DIN2(n32889), .Q(n35429) );
  or2s1 U27921 ( .DIN1(n35432), .DIN2(n35433), .Q(n35423) );
  or2s1 U27922 ( .DIN1(n35434), .DIN2(n35435), .Q(n35433) );
  and2s1 U27923 ( .DIN1(n35436), .DIN2(n35398), .Q(n35435) );
  and2s1 U27924 ( .DIN1(n35412), .DIN2(n35411), .Q(n35434) );
  or2s1 U27925 ( .DIN1(n35437), .DIN2(n35438), .Q(n35432) );
  and2s1 U27926 ( .DIN1(n35393), .DIN2(n32898), .Q(n35438) );
  or2s1 U27927 ( .DIN1(n35439), .DIN2(n35415), .Q(n32898) );
  and2s1 U27928 ( .DIN1(n33862), .DIN2(n35440), .Q(n35437) );
  or2s1 U27929 ( .DIN1(n35441), .DIN2(n35442), .Q(n35440) );
  hi1s1 U27930 ( .DIN1(n35443), .Q(n35442) );
  and2s1 U27931 ( .DIN1(u5_timer2[2]), .DIN2(n35422), .Q(n35441) );
  or2s1 U27932 ( .DIN1(n35444), .DIN2(n35445), .Q(n9237) );
  or2s1 U27933 ( .DIN1(n35446), .DIN2(n35447), .Q(n35445) );
  or2s1 U27934 ( .DIN1(n35448), .DIN2(n35449), .Q(n35447) );
  and2s1 U27935 ( .DIN1(n35388), .DIN2(n35377), .Q(n35449) );
  and2s1 U27936 ( .DIN1(n35393), .DIN2(n35450), .Q(n35448) );
  and2s1 U27937 ( .DIN1(n35451), .DIN2(n33865), .Q(n35446) );
  or2s1 U27938 ( .DIN1(n35452), .DIN2(n35453), .Q(n35444) );
  or2s1 U27939 ( .DIN1(n35454), .DIN2(n35455), .Q(n35453) );
  and2s1 U27940 ( .DIN1(n33859), .DIN2(n35456), .Q(n35455) );
  and2s1 U27941 ( .DIN1(n35398), .DIN2(n35457), .Q(n35454) );
  or2s1 U27942 ( .DIN1(n35458), .DIN2(n35459), .Q(n35452) );
  and2s1 U27943 ( .DIN1(n35412), .DIN2(n32889), .Q(n35459) );
  and2s1 U27944 ( .DIN1(n33862), .DIN2(n35460), .Q(n35458) );
  or2s1 U27945 ( .DIN1(n35461), .DIN2(n35462), .Q(n35460) );
  hi1s1 U27946 ( .DIN1(n35463), .Q(n35462) );
  and2s1 U27947 ( .DIN1(u5_timer2[3]), .DIN2(n35443), .Q(n35461) );
  or2s1 U27948 ( .DIN1(n35464), .DIN2(n35465), .Q(n9236) );
  or2s1 U27949 ( .DIN1(n35466), .DIN2(n35467), .Q(n35465) );
  or2s1 U27950 ( .DIN1(n35468), .DIN2(n35469), .Q(n35467) );
  and2s1 U27951 ( .DIN1(n35393), .DIN2(n35470), .Q(n35469) );
  and2s1 U27952 ( .DIN1(n35388), .DIN2(n33860), .Q(n35468) );
  and2s1 U27953 ( .DIN1(n35471), .DIN2(n33865), .Q(n35466) );
  or2s1 U27954 ( .DIN1(n35472), .DIN2(n35473), .Q(n35464) );
  or2s1 U27955 ( .DIN1(n35474), .DIN2(n35475), .Q(n35473) );
  and2s1 U27956 ( .DIN1(n35412), .DIN2(n35456), .Q(n35475) );
  and2s1 U27957 ( .DIN1(n35476), .DIN2(n34251), .Q(n35412) );
  hi1s1 U27958 ( .DIN1(n35398), .Q(n35476) );
  and2s1 U27959 ( .DIN1(n33862), .DIN2(n35477), .Q(n35474) );
  or2s1 U27960 ( .DIN1(n35478), .DIN2(n35479), .Q(n35477) );
  hi1s1 U27961 ( .DIN1(n35480), .Q(n35479) );
  and2s1 U27962 ( .DIN1(u5_timer2[4]), .DIN2(n35463), .Q(n35478) );
  and2s1 U27963 ( .DIN1(n33859), .DIN2(n35389), .Q(n35472) );
  or2s1 U27964 ( .DIN1(n35481), .DIN2(n35482), .Q(n9235) );
  or2s1 U27965 ( .DIN1(n35483), .DIN2(n35484), .Q(n35482) );
  and2s1 U27966 ( .DIN1(n35485), .DIN2(n33865), .Q(n35484) );
  and2s1 U27967 ( .DIN1(n33859), .DIN2(n32886), .Q(n35483) );
  or2s1 U27968 ( .DIN1(n35486), .DIN2(n35487), .Q(n35481) );
  and2s1 U27969 ( .DIN1(n35388), .DIN2(n32900), .Q(n35487) );
  or2s1 U27970 ( .DIN1(n35415), .DIN2(n35488), .Q(n32900) );
  or2s1 U27971 ( .DIN1(n35489), .DIN2(n35490), .Q(n35488) );
  and2s1 U27972 ( .DIN1(u0_sp_tms[25]), .DIN2(n35282), .Q(n35490) );
  and2s1 U27973 ( .DIN1(u0_tms[25]), .DIN2(n35283), .Q(n35489) );
  and2s1 U27974 ( .DIN1(n33862), .DIN2(n35491), .Q(n35486) );
  or2s1 U27975 ( .DIN1(n35492), .DIN2(n35493), .Q(n35491) );
  hi1s1 U27976 ( .DIN1(n35494), .Q(n35493) );
  and2s1 U27977 ( .DIN1(u5_timer2[5]), .DIN2(n35480), .Q(n35492) );
  or2s1 U27978 ( .DIN1(n35495), .DIN2(n35496), .Q(n9234) );
  or2s1 U27979 ( .DIN1(n35497), .DIN2(n35498), .Q(n35496) );
  and2s1 U27980 ( .DIN1(n33859), .DIN2(n35431), .Q(n35498) );
  and2s1 U27981 ( .DIN1(n33862), .DIN2(n35499), .Q(n35497) );
  or2s1 U27982 ( .DIN1(n35500), .DIN2(n35501), .Q(n35499) );
  hi1s1 U27983 ( .DIN1(n35381), .Q(n35501) );
  and2s1 U27984 ( .DIN1(u5_timer2[6]), .DIN2(n35494), .Q(n35500) );
  hi1s1 U27985 ( .DIN1(n35396), .Q(n33862) );
  or2s1 U27986 ( .DIN1(n35428), .DIN2(n35502), .Q(n35396) );
  or2s1 U27987 ( .DIN1(n33866), .DIN2(n33868), .Q(n35502) );
  or2s1 U27988 ( .DIN1(n35503), .DIN2(n35504), .Q(n33868) );
  or2s1 U27989 ( .DIN1(n35398), .DIN2(n35505), .Q(n35504) );
  or2s1 U27990 ( .DIN1(n35393), .DIN2(n33865), .Q(n35505) );
  or2s1 U27991 ( .DIN1(n35506), .DIN2(n34249), .Q(n35398) );
  and2s1 U27992 ( .DIN1(n34351), .DIN2(n15512), .Q(n35506) );
  or2s1 U27993 ( .DIN1(n34251), .DIN2(n35507), .Q(n35503) );
  or2s1 U27994 ( .DIN1(n35388), .DIN2(n33859), .Q(n35507) );
  and2s1 U27995 ( .DIN1(n32870), .DIN2(n35508), .Q(n33859) );
  and2s1 U27996 ( .DIN1(n35509), .DIN2(n35510), .Q(n35508) );
  or2s1 U27997 ( .DIN1(n35282), .DIN2(n35511), .Q(n35510) );
  and2s1 U27998 ( .DIN1(u0_csc[1]), .DIN2(n35512), .Q(n35511) );
  and2s1 U27999 ( .DIN1(n35513), .DIN2(u0_csc[2]), .Q(n35512) );
  hi1s1 U28000 ( .DIN1(u0_csc[3]), .Q(n35513) );
  or2s1 U28001 ( .DIN1(n35283), .DIN2(n35514), .Q(n35509) );
  and2s1 U28002 ( .DIN1(u0_sp_csc[2]), .DIN2(n35515), .Q(n35514) );
  and2s1 U28003 ( .DIN1(n35516), .DIN2(u0_sp_csc[1]), .Q(n35515) );
  hi1s1 U28004 ( .DIN1(u0_sp_csc[3]), .Q(n35516) );
  and2s1 U28005 ( .DIN1(u5_tmr2_done), .DIN2(n34351), .Q(n34251) );
  hi1s1 U28006 ( .DIN1(n35517), .Q(n33866) );
  or2s1 U28007 ( .DIN1(u5_timer2[8]), .DIN2(n33863), .Q(n35517) );
  or2s1 U28008 ( .DIN1(u5_timer2[7]), .DIN2(n35381), .Q(n33863) );
  or2s1 U28009 ( .DIN1(u5_timer2[6]), .DIN2(n35494), .Q(n35381) );
  or2s1 U28010 ( .DIN1(u5_timer2[5]), .DIN2(n35480), .Q(n35494) );
  or2s1 U28011 ( .DIN1(u5_timer2[4]), .DIN2(n35463), .Q(n35480) );
  or2s1 U28012 ( .DIN1(u5_timer2[3]), .DIN2(n35443), .Q(n35463) );
  or2s1 U28013 ( .DIN1(u5_timer2[2]), .DIN2(n35422), .Q(n35443) );
  or2s1 U28014 ( .DIN1(u5_timer2[0]), .DIN2(u5_timer2[1]), .Q(n35422) );
  or2s1 U28015 ( .DIN1(n35518), .DIN2(n34111), .Q(n35428) );
  and2s1 U28016 ( .DIN1(n35519), .DIN2(n32870), .Q(n35518) );
  and2s1 U28017 ( .DIN1(n35520), .DIN2(n35521), .Q(n35519) );
  or2s1 U28018 ( .DIN1(n35522), .DIN2(n35283), .Q(n35521) );
  and2s1 U28019 ( .DIN1(n35523), .DIN2(u0_sp_csc[1]), .Q(n35522) );
  hi1s1 U28020 ( .DIN1(n35524), .Q(n35523) );
  or2s1 U28021 ( .DIN1(u0_sp_csc[2]), .DIN2(u0_sp_csc[3]), .Q(n35524) );
  or2s1 U28022 ( .DIN1(n35525), .DIN2(n35282), .Q(n35520) );
  and2s1 U28023 ( .DIN1(u0_csc[1]), .DIN2(n34681), .Q(n35525) );
  hi1s1 U28024 ( .DIN1(n34685), .Q(n34681) );
  and2s1 U28025 ( .DIN1(n32885), .DIN2(n33865), .Q(n35495) );
  and2s1 U28026 ( .DIN1(n35526), .DIN2(n9141), .Q(n9233) );
  or2s1 U28027 ( .DIN1(n35527), .DIN2(n9142), .Q(n9232) );
  and2s1 U28028 ( .DIN1(n35526), .DIN2(n9143), .Q(n9231) );
  or2s1 U28029 ( .DIN1(n35527), .DIN2(n9144), .Q(n9230) );
  or2s1 U28030 ( .DIN1(n35528), .DIN2(n35529), .Q(n9229) );
  and2s1 U28031 ( .DIN1(wb_data_i[31]), .DIN2(n35527), .Q(n35529) );
  and2s1 U28032 ( .DIN1(n35526), .DIN2(n9176), .Q(n35528) );
  or2s1 U28033 ( .DIN1(n35530), .DIN2(n35531), .Q(n9228) );
  and2s1 U28034 ( .DIN1(wb_data_i[30]), .DIN2(n35527), .Q(n35531) );
  and2s1 U28035 ( .DIN1(n35526), .DIN2(n9175), .Q(n35530) );
  or2s1 U28036 ( .DIN1(n35532), .DIN2(n35533), .Q(n9227) );
  and2s1 U28037 ( .DIN1(wb_data_i[29]), .DIN2(n35527), .Q(n35533) );
  and2s1 U28038 ( .DIN1(n35526), .DIN2(n9174), .Q(n35532) );
  or2s1 U28039 ( .DIN1(n35534), .DIN2(n35535), .Q(n9226) );
  and2s1 U28040 ( .DIN1(wb_data_i[28]), .DIN2(n35527), .Q(n35535) );
  and2s1 U28041 ( .DIN1(n35526), .DIN2(n9173), .Q(n35534) );
  or2s1 U28042 ( .DIN1(n35536), .DIN2(n35537), .Q(n9225) );
  and2s1 U28043 ( .DIN1(wb_data_i[27]), .DIN2(n35527), .Q(n35537) );
  and2s1 U28044 ( .DIN1(n35526), .DIN2(n9172), .Q(n35536) );
  or2s1 U28045 ( .DIN1(n35538), .DIN2(n35539), .Q(n9224) );
  and2s1 U28046 ( .DIN1(wb_data_i[26]), .DIN2(n35527), .Q(n35539) );
  and2s1 U28047 ( .DIN1(n35526), .DIN2(n9171), .Q(n35538) );
  or2s1 U28048 ( .DIN1(n35540), .DIN2(n35541), .Q(n9223) );
  and2s1 U28049 ( .DIN1(wb_data_i[25]), .DIN2(n35527), .Q(n35541) );
  and2s1 U28050 ( .DIN1(n35526), .DIN2(n9170), .Q(n35540) );
  or2s1 U28051 ( .DIN1(n35542), .DIN2(n35543), .Q(n9222) );
  and2s1 U28052 ( .DIN1(wb_data_i[24]), .DIN2(n35527), .Q(n35543) );
  and2s1 U28053 ( .DIN1(n35526), .DIN2(n9169), .Q(n35542) );
  or2s1 U28054 ( .DIN1(n35544), .DIN2(n35545), .Q(n9221) );
  and2s1 U28055 ( .DIN1(wb_data_i[23]), .DIN2(n35527), .Q(n35545) );
  and2s1 U28056 ( .DIN1(n35526), .DIN2(n9168), .Q(n35544) );
  or2s1 U28057 ( .DIN1(n35546), .DIN2(n35547), .Q(n9220) );
  and2s1 U28058 ( .DIN1(wb_data_i[22]), .DIN2(n35527), .Q(n35547) );
  and2s1 U28059 ( .DIN1(n35526), .DIN2(n9167), .Q(n35546) );
  or2s1 U28060 ( .DIN1(n35548), .DIN2(n35549), .Q(n9219) );
  and2s1 U28061 ( .DIN1(wb_data_i[21]), .DIN2(n35527), .Q(n35549) );
  and2s1 U28062 ( .DIN1(n35526), .DIN2(n9166), .Q(n35548) );
  or2s1 U28063 ( .DIN1(n35550), .DIN2(n35551), .Q(n9218) );
  and2s1 U28064 ( .DIN1(wb_data_i[20]), .DIN2(n35527), .Q(n35551) );
  and2s1 U28065 ( .DIN1(n35526), .DIN2(n9165), .Q(n35550) );
  or2s1 U28066 ( .DIN1(n35552), .DIN2(n35553), .Q(n9217) );
  and2s1 U28067 ( .DIN1(wb_data_i[19]), .DIN2(n35527), .Q(n35553) );
  and2s1 U28068 ( .DIN1(n35526), .DIN2(n9164), .Q(n35552) );
  or2s1 U28069 ( .DIN1(n35554), .DIN2(n35555), .Q(n9216) );
  and2s1 U28070 ( .DIN1(wb_data_i[18]), .DIN2(n35527), .Q(n35555) );
  and2s1 U28071 ( .DIN1(n35526), .DIN2(n9163), .Q(n35554) );
  or2s1 U28072 ( .DIN1(n35556), .DIN2(n35557), .Q(n9215) );
  and2s1 U28073 ( .DIN1(wb_data_i[17]), .DIN2(n35527), .Q(n35557) );
  and2s1 U28074 ( .DIN1(n35526), .DIN2(n9162), .Q(n35556) );
  or2s1 U28075 ( .DIN1(n35558), .DIN2(n35559), .Q(n9214) );
  and2s1 U28076 ( .DIN1(wb_data_i[16]), .DIN2(n35527), .Q(n35559) );
  and2s1 U28077 ( .DIN1(n35526), .DIN2(n9161), .Q(n35558) );
  or2s1 U28078 ( .DIN1(n35560), .DIN2(n35561), .Q(n9213) );
  and2s1 U28079 ( .DIN1(wb_data_i[15]), .DIN2(n35527), .Q(n35561) );
  and2s1 U28080 ( .DIN1(n35526), .DIN2(n9160), .Q(n35560) );
  or2s1 U28081 ( .DIN1(n35562), .DIN2(n35563), .Q(n9212) );
  and2s1 U28082 ( .DIN1(wb_data_i[14]), .DIN2(n35527), .Q(n35563) );
  and2s1 U28083 ( .DIN1(n35526), .DIN2(n9159), .Q(n35562) );
  or2s1 U28084 ( .DIN1(n35564), .DIN2(n35565), .Q(n9211) );
  and2s1 U28085 ( .DIN1(wb_data_i[13]), .DIN2(n35527), .Q(n35565) );
  and2s1 U28086 ( .DIN1(n35526), .DIN2(n9158), .Q(n35564) );
  or2s1 U28087 ( .DIN1(n35566), .DIN2(n35567), .Q(n9210) );
  and2s1 U28088 ( .DIN1(wb_data_i[12]), .DIN2(n35527), .Q(n35567) );
  and2s1 U28089 ( .DIN1(n35526), .DIN2(n9157), .Q(n35566) );
  or2s1 U28090 ( .DIN1(n35568), .DIN2(n35569), .Q(n9209) );
  and2s1 U28091 ( .DIN1(wb_data_i[11]), .DIN2(n35527), .Q(n35569) );
  and2s1 U28092 ( .DIN1(n35526), .DIN2(n9156), .Q(n35568) );
  or2s1 U28093 ( .DIN1(n35570), .DIN2(n35571), .Q(n9208) );
  and2s1 U28094 ( .DIN1(wb_data_i[10]), .DIN2(n35527), .Q(n35571) );
  and2s1 U28095 ( .DIN1(n35526), .DIN2(n9155), .Q(n35570) );
  or2s1 U28096 ( .DIN1(n35572), .DIN2(n35573), .Q(n9207) );
  and2s1 U28097 ( .DIN1(wb_data_i[9]), .DIN2(n35527), .Q(n35573) );
  and2s1 U28098 ( .DIN1(n35526), .DIN2(n9154), .Q(n35572) );
  or2s1 U28099 ( .DIN1(n35574), .DIN2(n35575), .Q(n9206) );
  and2s1 U28100 ( .DIN1(wb_data_i[8]), .DIN2(n35527), .Q(n35575) );
  and2s1 U28101 ( .DIN1(n35526), .DIN2(n9153), .Q(n35574) );
  or2s1 U28102 ( .DIN1(n35576), .DIN2(n35577), .Q(n9205) );
  and2s1 U28103 ( .DIN1(wb_data_i[7]), .DIN2(n35527), .Q(n35577) );
  and2s1 U28104 ( .DIN1(n35526), .DIN2(n9152), .Q(n35576) );
  or2s1 U28105 ( .DIN1(n35578), .DIN2(n35579), .Q(n9204) );
  and2s1 U28106 ( .DIN1(wb_data_i[6]), .DIN2(n35527), .Q(n35579) );
  and2s1 U28107 ( .DIN1(n35526), .DIN2(n9151), .Q(n35578) );
  or2s1 U28108 ( .DIN1(n35580), .DIN2(n35581), .Q(n9203) );
  and2s1 U28109 ( .DIN1(wb_data_i[5]), .DIN2(n35527), .Q(n35581) );
  and2s1 U28110 ( .DIN1(n35526), .DIN2(n9150), .Q(n35580) );
  or2s1 U28111 ( .DIN1(n35582), .DIN2(n35583), .Q(n9202) );
  and2s1 U28112 ( .DIN1(wb_data_i[4]), .DIN2(n35527), .Q(n35583) );
  and2s1 U28113 ( .DIN1(n35526), .DIN2(n9149), .Q(n35582) );
  or2s1 U28114 ( .DIN1(n35584), .DIN2(n35585), .Q(n9201) );
  and2s1 U28115 ( .DIN1(wb_data_i[3]), .DIN2(n35527), .Q(n35585) );
  and2s1 U28116 ( .DIN1(n35526), .DIN2(n9148), .Q(n35584) );
  or2s1 U28117 ( .DIN1(n35586), .DIN2(n35587), .Q(n9200) );
  and2s1 U28118 ( .DIN1(wb_data_i[2]), .DIN2(n35527), .Q(n35587) );
  and2s1 U28119 ( .DIN1(n35526), .DIN2(n9147), .Q(n35586) );
  or2s1 U28120 ( .DIN1(n35588), .DIN2(n35589), .Q(n9199) );
  and2s1 U28121 ( .DIN1(wb_data_i[1]), .DIN2(n35527), .Q(n35589) );
  and2s1 U28122 ( .DIN1(n35526), .DIN2(n9146), .Q(n35588) );
  or2s1 U28123 ( .DIN1(n35590), .DIN2(n35591), .Q(n9198) );
  and2s1 U28124 ( .DIN1(wb_data_i[0]), .DIN2(n35527), .Q(n35591) );
  and2s1 U28125 ( .DIN1(n35526), .DIN2(n9145), .Q(n35590) );
  hi1s1 U28126 ( .DIN1(n35527), .Q(n35526) );
  or2s1 U28127 ( .DIN1(n34685), .DIN2(n35592), .Q(n35527) );
  or2s1 U28128 ( .DIN1(u0_csc[1]), .DIN2(n15482), .Q(n35592) );
  or2s1 U28129 ( .DIN1(u0_csc[2]), .DIN2(u0_csc[3]), .Q(n34685) );
  or2s1 U28130 ( .DIN1(n35593), .DIN2(n35594), .Q(n9195) );
  and2s1 U28131 ( .DIN1(n35054), .DIN2(n4536), .Q(n35594) );
  and2s1 U28132 ( .DIN1(n15502), .DIN2(n9197), .Q(n35593) );
  or2s1 U28133 ( .DIN1(n35595), .DIN2(n35596), .Q(n9197) );
  or2s1 U28134 ( .DIN1(n32907), .DIN2(n35597), .Q(n35596) );
  or2s1 U28135 ( .DIN1(n35598), .DIN2(n35599), .Q(n35595) );
  and2s1 U28136 ( .DIN1(n35600), .DIN2(n35052), .Q(n9194) );
  or2s1 U28137 ( .DIN1(n32869), .DIN2(n32907), .Q(n35600) );
  or2s1 U28138 ( .DIN1(n35601), .DIN2(n35602), .Q(n9193) );
  or2s1 U28139 ( .DIN1(n35603), .DIN2(n35604), .Q(n35602) );
  or2s1 U28140 ( .DIN1(n35605), .DIN2(n35606), .Q(n35604) );
  and2s1 U28141 ( .DIN1(u5_cke_r), .DIN2(n32907), .Q(n35606) );
  and2s1 U28142 ( .DIN1(n35607), .DIN2(n35052), .Q(n35605) );
  or2s1 U28143 ( .DIN1(n35608), .DIN2(n32943), .Q(n35607) );
  and2s1 U28144 ( .DIN1(n32940), .DIN2(n33017), .Q(n35608) );
  and2s1 U28145 ( .DIN1(u5_wb_cycle), .DIN2(n32934), .Q(n33017) );
  hi1s1 U28146 ( .DIN1(n32957), .Q(n32934) );
  or2s1 U28147 ( .DIN1(n34574), .DIN2(n35609), .Q(n35601) );
  or2s1 U28148 ( .DIN1(n35610), .DIN2(n35611), .Q(n9192) );
  and2s1 U28149 ( .DIN1(n32878), .DIN2(n33864), .Q(n35611) );
  or2s1 U28150 ( .DIN1(n35415), .DIN2(n35612), .Q(n33864) );
  or2s1 U28151 ( .DIN1(n35613), .DIN2(n35614), .Q(n35612) );
  and2s1 U28152 ( .DIN1(u0_sp_tms[7]), .DIN2(n35282), .Q(n35614) );
  and2s1 U28153 ( .DIN1(u0_tms[7]), .DIN2(n35283), .Q(n35613) );
  and2s1 U28154 ( .DIN1(u5_timer[7]), .DIN2(n35615), .Q(n35610) );
  or2s1 U28155 ( .DIN1(n35616), .DIN2(n35617), .Q(n35615) );
  and2s1 U28156 ( .DIN1(n32916), .DIN2(n35618), .Q(n35616) );
  or2s1 U28157 ( .DIN1(n35619), .DIN2(n35620), .Q(n9191) );
  or2s1 U28158 ( .DIN1(n35621), .DIN2(n35622), .Q(n35620) );
  or2s1 U28159 ( .DIN1(n35623), .DIN2(n32877), .Q(n35622) );
  and2s1 U28160 ( .DIN1(n32878), .DIN2(n35406), .Q(n35623) );
  or2s1 U28161 ( .DIN1(n35624), .DIN2(n35625), .Q(n35621) );
  or2s1 U28162 ( .DIN1(n35626), .DIN2(n35627), .Q(n35625) );
  and2s1 U28163 ( .DIN1(n32916), .DIN2(n35628), .Q(n35627) );
  hi1s1 U28164 ( .DIN1(u5_timer[0]), .Q(n35628) );
  and2s1 U28165 ( .DIN1(n35617), .DIN2(u5_timer[0]), .Q(n35626) );
  and2s1 U28166 ( .DIN1(n32888), .DIN2(n35411), .Q(n35624) );
  or2s1 U28167 ( .DIN1(n35629), .DIN2(n35630), .Q(n35619) );
  or2s1 U28168 ( .DIN1(n35631), .DIN2(n35632), .Q(n35630) );
  or2s1 U28169 ( .DIN1(n35633), .DIN2(n35634), .Q(n35632) );
  and2s1 U28170 ( .DIN1(n35389), .DIN2(n32887), .Q(n35634) );
  and2s1 U28171 ( .DIN1(n35405), .DIN2(n32899), .Q(n35633) );
  or2s1 U28172 ( .DIN1(n35415), .DIN2(n35635), .Q(n35405) );
  or2s1 U28173 ( .DIN1(n35636), .DIN2(n35637), .Q(n35635) );
  and2s1 U28174 ( .DIN1(u0_sp_tms[8]), .DIN2(n35282), .Q(n35637) );
  and2s1 U28175 ( .DIN1(u0_tms[8]), .DIN2(n35283), .Q(n35636) );
  and2s1 U28176 ( .DIN1(n32884), .DIN2(n35485), .Q(n35631) );
  or2s1 U28177 ( .DIN1(n35638), .DIN2(n35639), .Q(n35629) );
  or2s1 U28178 ( .DIN1(n35640), .DIN2(n35641), .Q(n35639) );
  and2s1 U28179 ( .DIN1(n33860), .DIN2(n32901), .Q(n35641) );
  or2s1 U28180 ( .DIN1(n35415), .DIN2(n35642), .Q(n33860) );
  or2s1 U28181 ( .DIN1(n35643), .DIN2(n35644), .Q(n35642) );
  and2s1 U28182 ( .DIN1(u0_sp_tms[24]), .DIN2(n35282), .Q(n35644) );
  and2s1 U28183 ( .DIN1(u0_tms[24]), .DIN2(n35283), .Q(n35643) );
  and2s1 U28184 ( .DIN1(n35645), .DIN2(n32907), .Q(n35640) );
  or2s1 U28185 ( .DIN1(n35646), .DIN2(n35647), .Q(n35645) );
  and2s1 U28186 ( .DIN1(n32913), .DIN2(n35457), .Q(n35647) );
  hi1s1 U28187 ( .DIN1(n35389), .Q(n32913) );
  and2s1 U28188 ( .DIN1(n32914), .DIN2(n35389), .Q(n35646) );
  hi1s1 U28189 ( .DIN1(n35457), .Q(n32914) );
  and2s1 U28190 ( .DIN1(n32896), .DIN2(n35397), .Q(n35638) );
  or2s1 U28191 ( .DIN1(n35415), .DIN2(n35648), .Q(n35397) );
  or2s1 U28192 ( .DIN1(n35649), .DIN2(n35650), .Q(n35648) );
  and2s1 U28193 ( .DIN1(u0_sp_tms[12]), .DIN2(n35282), .Q(n35650) );
  and2s1 U28194 ( .DIN1(u0_tms[12]), .DIN2(n35283), .Q(n35649) );
  or2s1 U28195 ( .DIN1(n35651), .DIN2(n35652), .Q(n9190) );
  or2s1 U28196 ( .DIN1(n35653), .DIN2(n35654), .Q(n35652) );
  or2s1 U28197 ( .DIN1(n35655), .DIN2(n35656), .Q(n35654) );
  and2s1 U28198 ( .DIN1(n32878), .DIN2(n35451), .Q(n35655) );
  or2s1 U28199 ( .DIN1(n35657), .DIN2(n35658), .Q(n35653) );
  or2s1 U28200 ( .DIN1(n35659), .DIN2(n35660), .Q(n35658) );
  and2s1 U28201 ( .DIN1(n32916), .DIN2(n35661), .Q(n35660) );
  and2s1 U28202 ( .DIN1(n32896), .DIN2(n35436), .Q(n35659) );
  or2s1 U28203 ( .DIN1(n35415), .DIN2(n35662), .Q(n35436) );
  or2s1 U28204 ( .DIN1(n35663), .DIN2(n35664), .Q(n35662) );
  and2s1 U28205 ( .DIN1(u0_sp_tms[14]), .DIN2(n35282), .Q(n35664) );
  and2s1 U28206 ( .DIN1(u0_tms[14]), .DIN2(n35283), .Q(n35663) );
  and2s1 U28207 ( .DIN1(n32888), .DIN2(n35456), .Q(n35657) );
  or2s1 U28208 ( .DIN1(n35665), .DIN2(n35666), .Q(n35651) );
  or2s1 U28209 ( .DIN1(n35667), .DIN2(n35668), .Q(n35666) );
  and2s1 U28210 ( .DIN1(n35450), .DIN2(n32899), .Q(n35668) );
  or2s1 U28211 ( .DIN1(n35415), .DIN2(n35669), .Q(n35450) );
  or2s1 U28212 ( .DIN1(n35670), .DIN2(n35671), .Q(n35669) );
  and2s1 U28213 ( .DIN1(u0_sp_tms[10]), .DIN2(n35282), .Q(n35671) );
  and2s1 U28214 ( .DIN1(u0_tms[10]), .DIN2(n35283), .Q(n35670) );
  and2s1 U28215 ( .DIN1(n35672), .DIN2(n35431), .Q(n35667) );
  or2s1 U28216 ( .DIN1(n35673), .DIN2(n35674), .Q(n35665) );
  or2s1 U28217 ( .DIN1(n35675), .DIN2(n35676), .Q(n35674) );
  and2s1 U28218 ( .DIN1(u5_timer[2]), .DIN2(n35677), .Q(n35676) );
  or2s1 U28219 ( .DIN1(n35678), .DIN2(n32918), .Q(n35677) );
  or2s1 U28220 ( .DIN1(n35679), .DIN2(n35617), .Q(n32918) );
  and2s1 U28221 ( .DIN1(u5_timer[0]), .DIN2(n32916), .Q(n35679) );
  and2s1 U28222 ( .DIN1(u5_timer[1]), .DIN2(n32916), .Q(n35678) );
  and2s1 U28223 ( .DIN1(n35680), .DIN2(n35681), .Q(n35675) );
  and2s1 U28224 ( .DIN1(n35682), .DIN2(n32907), .Q(n35680) );
  and2s1 U28225 ( .DIN1(n35683), .DIN2(n32901), .Q(n35673) );
  or2s1 U28226 ( .DIN1(n35415), .DIN2(n35684), .Q(n35683) );
  or2s1 U28227 ( .DIN1(n35685), .DIN2(n35686), .Q(n35684) );
  and2s1 U28228 ( .DIN1(u0_sp_tms[26]), .DIN2(n35282), .Q(n35686) );
  and2s1 U28229 ( .DIN1(u0_tms[26]), .DIN2(n35283), .Q(n35685) );
  or2s1 U28230 ( .DIN1(n35687), .DIN2(n35688), .Q(n9189) );
  or2s1 U28231 ( .DIN1(n35689), .DIN2(n35690), .Q(n35688) );
  or2s1 U28232 ( .DIN1(n35691), .DIN2(n35692), .Q(n35690) );
  and2s1 U28233 ( .DIN1(n32896), .DIN2(n35457), .Q(n35692) );
  and2s1 U28234 ( .DIN1(n32878), .DIN2(n35471), .Q(n35691) );
  or2s1 U28235 ( .DIN1(n35415), .DIN2(n35693), .Q(n35471) );
  or2s1 U28236 ( .DIN1(n35694), .DIN2(n35695), .Q(n35693) );
  and2s1 U28237 ( .DIN1(u0_sp_tms[3]), .DIN2(n35282), .Q(n35695) );
  and2s1 U28238 ( .DIN1(u0_tms[3]), .DIN2(n35283), .Q(n35694) );
  or2s1 U28239 ( .DIN1(n35696), .DIN2(n35697), .Q(n35689) );
  and2s1 U28240 ( .DIN1(n35470), .DIN2(n32899), .Q(n35697) );
  or2s1 U28241 ( .DIN1(n35415), .DIN2(n35698), .Q(n35470) );
  or2s1 U28242 ( .DIN1(n35699), .DIN2(n35700), .Q(n35698) );
  and2s1 U28243 ( .DIN1(u0_sp_tms[11]), .DIN2(n35282), .Q(n35700) );
  and2s1 U28244 ( .DIN1(u0_tms[11]), .DIN2(n35283), .Q(n35699) );
  and2s1 U28245 ( .DIN1(n35672), .DIN2(n35377), .Q(n35696) );
  or2s1 U28246 ( .DIN1(n35701), .DIN2(n32887), .Q(n35672) );
  and2s1 U28247 ( .DIN1(n35702), .DIN2(n32907), .Q(n35701) );
  hi1s1 U28248 ( .DIN1(n35682), .Q(n35702) );
  or2s1 U28249 ( .DIN1(n35703), .DIN2(n35704), .Q(n35687) );
  or2s1 U28250 ( .DIN1(n35705), .DIN2(n35706), .Q(n35704) );
  and2s1 U28251 ( .DIN1(n35707), .DIN2(n32901), .Q(n35706) );
  or2s1 U28252 ( .DIN1(n35415), .DIN2(n35708), .Q(n35707) );
  or2s1 U28253 ( .DIN1(n35709), .DIN2(n35710), .Q(n35708) );
  and2s1 U28254 ( .DIN1(u0_sp_tms[27]), .DIN2(n35282), .Q(n35710) );
  and2s1 U28255 ( .DIN1(u0_tms[27]), .DIN2(n35283), .Q(n35709) );
  and2s1 U28256 ( .DIN1(u5_timer[3]), .DIN2(n35711), .Q(n35705) );
  or2s1 U28257 ( .DIN1(n35712), .DIN2(n35713), .Q(n35703) );
  and2s1 U28258 ( .DIN1(n35714), .DIN2(n32907), .Q(n35713) );
  or2s1 U28259 ( .DIN1(n35715), .DIN2(n35716), .Q(n35714) );
  and2s1 U28260 ( .DIN1(n35681), .DIN2(n35377), .Q(n35716) );
  hi1s1 U28261 ( .DIN1(n35431), .Q(n35681) );
  and2s1 U28262 ( .DIN1(n35717), .DIN2(n35718), .Q(n35715) );
  hi1s1 U28263 ( .DIN1(n35377), .Q(n35718) );
  or2s1 U28264 ( .DIN1(n35415), .DIN2(n35719), .Q(n35377) );
  or2s1 U28265 ( .DIN1(n35720), .DIN2(n35721), .Q(n35719) );
  and2s1 U28266 ( .DIN1(u0_sp_tms[23]), .DIN2(n35282), .Q(n35721) );
  and2s1 U28267 ( .DIN1(u0_tms[23]), .DIN2(n35283), .Q(n35720) );
  and2s1 U28268 ( .DIN1(n35682), .DIN2(n35431), .Q(n35717) );
  or2s1 U28269 ( .DIN1(n35415), .DIN2(n35722), .Q(n35431) );
  or2s1 U28270 ( .DIN1(n35723), .DIN2(n35724), .Q(n35722) );
  and2s1 U28271 ( .DIN1(u0_sp_tms[22]), .DIN2(n35282), .Q(n35724) );
  and2s1 U28272 ( .DIN1(u0_tms[22]), .DIN2(n35283), .Q(n35723) );
  or2s1 U28273 ( .DIN1(n35725), .DIN2(n35726), .Q(n35682) );
  and2s1 U28274 ( .DIN1(n35390), .DIN2(n32886), .Q(n35726) );
  and2s1 U28275 ( .DIN1(n35727), .DIN2(n32910), .Q(n35725) );
  or2s1 U28276 ( .DIN1(n35728), .DIN2(n35729), .Q(n32910) );
  hi1s1 U28277 ( .DIN1(n35730), .Q(n35729) );
  or2s1 U28278 ( .DIN1(n35390), .DIN2(n35731), .Q(n35730) );
  and2s1 U28279 ( .DIN1(n35731), .DIN2(n35390), .Q(n35728) );
  hi1s1 U28280 ( .DIN1(n32886), .Q(n35731) );
  or2s1 U28281 ( .DIN1(n35415), .DIN2(n35732), .Q(n32886) );
  or2s1 U28282 ( .DIN1(n35733), .DIN2(n35734), .Q(n35732) );
  and2s1 U28283 ( .DIN1(u0_sp_tms[21]), .DIN2(n35282), .Q(n35734) );
  and2s1 U28284 ( .DIN1(u0_tms[21]), .DIN2(n35283), .Q(n35733) );
  and2s1 U28285 ( .DIN1(n35389), .DIN2(n35457), .Q(n35727) );
  or2s1 U28286 ( .DIN1(n35415), .DIN2(n35735), .Q(n35457) );
  or2s1 U28287 ( .DIN1(n35736), .DIN2(n35737), .Q(n35735) );
  and2s1 U28288 ( .DIN1(u0_sp_tms[15]), .DIN2(n35282), .Q(n35737) );
  and2s1 U28289 ( .DIN1(u0_tms[15]), .DIN2(n35283), .Q(n35736) );
  or2s1 U28290 ( .DIN1(n35415), .DIN2(n35738), .Q(n35389) );
  or2s1 U28291 ( .DIN1(n35739), .DIN2(n35740), .Q(n35738) );
  and2s1 U28292 ( .DIN1(u0_sp_tms[20]), .DIN2(n35282), .Q(n35740) );
  and2s1 U28293 ( .DIN1(u0_tms[20]), .DIN2(n35283), .Q(n35739) );
  and2s1 U28294 ( .DIN1(n35741), .DIN2(n32916), .Q(n35712) );
  and2s1 U28295 ( .DIN1(n35661), .DIN2(n35742), .Q(n35741) );
  hi1s1 U28296 ( .DIN1(u5_timer[3]), .Q(n35742) );
  hi1s1 U28297 ( .DIN1(n35743), .Q(n35661) );
  or2s1 U28298 ( .DIN1(n35744), .DIN2(n35745), .Q(n9188) );
  or2s1 U28299 ( .DIN1(n35746), .DIN2(n35747), .Q(n35745) );
  and2s1 U28300 ( .DIN1(n32878), .DIN2(n35485), .Q(n35747) );
  or2s1 U28301 ( .DIN1(n35415), .DIN2(n35748), .Q(n35485) );
  or2s1 U28302 ( .DIN1(n35749), .DIN2(n35750), .Q(n35748) );
  and2s1 U28303 ( .DIN1(u0_sp_tms[4]), .DIN2(n35282), .Q(n35750) );
  and2s1 U28304 ( .DIN1(u0_tms[4]), .DIN2(n35283), .Q(n35749) );
  and2s1 U28305 ( .DIN1(u5_timer[4]), .DIN2(n35751), .Q(n35746) );
  or2s1 U28306 ( .DIN1(n35752), .DIN2(n35711), .Q(n35751) );
  or2s1 U28307 ( .DIN1(n35753), .DIN2(n35617), .Q(n35711) );
  and2s1 U28308 ( .DIN1(n32916), .DIN2(n35743), .Q(n35753) );
  and2s1 U28309 ( .DIN1(u5_timer[3]), .DIN2(n32916), .Q(n35752) );
  and2s1 U28310 ( .DIN1(n32916), .DIN2(n35754), .Q(n35744) );
  or2s1 U28311 ( .DIN1(n35755), .DIN2(n35756), .Q(n9187) );
  or2s1 U28312 ( .DIN1(n35757), .DIN2(n35758), .Q(n35756) );
  and2s1 U28313 ( .DIN1(u5_timer[5]), .DIN2(n35759), .Q(n35758) );
  and2s1 U28314 ( .DIN1(n35760), .DIN2(n32916), .Q(n35757) );
  and2s1 U28315 ( .DIN1(n35754), .DIN2(n35761), .Q(n35760) );
  hi1s1 U28316 ( .DIN1(u5_timer[5]), .Q(n35761) );
  hi1s1 U28317 ( .DIN1(n35762), .Q(n35754) );
  and2s1 U28318 ( .DIN1(n32878), .DIN2(n32885), .Q(n35755) );
  or2s1 U28319 ( .DIN1(n35415), .DIN2(n35763), .Q(n32885) );
  or2s1 U28320 ( .DIN1(n35764), .DIN2(n35765), .Q(n35763) );
  and2s1 U28321 ( .DIN1(u0_sp_tms[5]), .DIN2(n35282), .Q(n35765) );
  and2s1 U28322 ( .DIN1(u0_tms[5]), .DIN2(n35283), .Q(n35764) );
  or2s1 U28323 ( .DIN1(n35766), .DIN2(n35767), .Q(n9186) );
  or2s1 U28324 ( .DIN1(n35768), .DIN2(n35769), .Q(n35767) );
  and2s1 U28325 ( .DIN1(n32878), .DIN2(n35382), .Q(n35769) );
  or2s1 U28326 ( .DIN1(n35415), .DIN2(n35770), .Q(n35382) );
  or2s1 U28327 ( .DIN1(n35771), .DIN2(n35772), .Q(n35770) );
  and2s1 U28328 ( .DIN1(u0_sp_tms[6]), .DIN2(n35282), .Q(n35772) );
  and2s1 U28329 ( .DIN1(u0_tms[6]), .DIN2(n35283), .Q(n35771) );
  and2s1 U28330 ( .DIN1(u5_timer[6]), .DIN2(n35773), .Q(n35768) );
  or2s1 U28331 ( .DIN1(n35774), .DIN2(n35759), .Q(n35773) );
  or2s1 U28332 ( .DIN1(n35775), .DIN2(n35617), .Q(n35759) );
  and2s1 U28333 ( .DIN1(n35776), .DIN2(n35777), .Q(n35617) );
  hi1s1 U28334 ( .DIN1(n35778), .Q(n35777) );
  and2s1 U28335 ( .DIN1(n32916), .DIN2(n35762), .Q(n35775) );
  and2s1 U28336 ( .DIN1(u5_timer[5]), .DIN2(n32916), .Q(n35774) );
  and2s1 U28337 ( .DIN1(n32916), .DIN2(n35779), .Q(n35766) );
  hi1s1 U28338 ( .DIN1(n35776), .Q(n32916) );
  or2s1 U28339 ( .DIN1(n32970), .DIN2(n35780), .Q(n35776) );
  or2s1 U28340 ( .DIN1(n19412), .DIN2(n35778), .Q(n35780) );
  or2s1 U28341 ( .DIN1(n35781), .DIN2(n35782), .Q(n35778) );
  or2s1 U28342 ( .DIN1(n32899), .DIN2(n33875), .Q(n35782) );
  or2s1 U28343 ( .DIN1(n32896), .DIN2(n32878), .Q(n33875) );
  or2s1 U28344 ( .DIN1(n34333), .DIN2(n33007), .Q(n32899) );
  and2s1 U28345 ( .DIN1(u5_tmr_done), .DIN2(n34368), .Q(n34333) );
  or2s1 U28346 ( .DIN1(n32877), .DIN2(n35783), .Q(n35781) );
  or2s1 U28347 ( .DIN1(n32907), .DIN2(n35784), .Q(n35783) );
  or2s1 U28348 ( .DIN1(n32865), .DIN2(n35656), .Q(n32877) );
  hi1s1 U28349 ( .DIN1(n9764), .Q(n32970) );
  or2s1 U28350 ( .DIN1(n35785), .DIN2(n35786), .Q(n9185) );
  or2s1 U28351 ( .DIN1(n35787), .DIN2(n35788), .Q(n9178) );
  or2s1 U28352 ( .DIN1(n34261), .DIN2(n34263), .Q(n35788) );
  and2s1 U28353 ( .DIN1(n35789), .DIN2(n35790), .Q(n35787) );
  and2s1 U28354 ( .DIN1(n34577), .DIN2(n33919), .Q(n35790) );
  hi1s1 U28355 ( .DIN1(n36662), .Q(n33919) );
  hi1s1 U28356 ( .DIN1(n35313), .Q(n34577) );
  or2s1 U28357 ( .DIN1(u4_rfr_req), .DIN2(u0_init_req), .Q(n35313) );
  and2s1 U28358 ( .DIN1(n15515), .DIN2(n32865), .Q(n35789) );
  and2s1 U28359 ( .DIN1(n35791), .DIN2(n9689), .Q(n9177) );
  and2s1 U28360 ( .DIN1(n35792), .DIN2(n34322), .Q(n35791) );
  or2s1 U28361 ( .DIN1(n35793), .DIN2(n35794), .Q(n9140) );
  or2s1 U28362 ( .DIN1(n35795), .DIN2(n35796), .Q(n35794) );
  and2s1 U28363 ( .DIN1(n35797), .DIN2(n32539), .Q(n35796) );
  hi1s1 U28364 ( .DIN1(n36663), .Q(n32539) );
  and2s1 U28365 ( .DIN1(n35798), .DIN2(wb_addr_i[25]), .Q(n35795) );
  and2s1 U28366 ( .DIN1(n35799), .DIN2(n34942), .Q(n35793) );
  hi1s1 U28367 ( .DIN1(n36664), .Q(n34942) );
  or2s1 U28368 ( .DIN1(n35800), .DIN2(n35801), .Q(n9139) );
  or2s1 U28369 ( .DIN1(n35802), .DIN2(n35803), .Q(n35801) );
  and2s1 U28370 ( .DIN1(n35797), .DIN2(n32543), .Q(n35803) );
  hi1s1 U28371 ( .DIN1(n36665), .Q(n32543) );
  and2s1 U28372 ( .DIN1(n35798), .DIN2(wb_addr_i[24]), .Q(n35802) );
  and2s1 U28373 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[22]), .Q(n35800) );
  or2s1 U28374 ( .DIN1(n35804), .DIN2(n35805), .Q(n9138) );
  or2s1 U28375 ( .DIN1(n35806), .DIN2(n35807), .Q(n35805) );
  and2s1 U28376 ( .DIN1(n35797), .DIN2(n32546), .Q(n35807) );
  hi1s1 U28377 ( .DIN1(n36666), .Q(n32546) );
  and2s1 U28378 ( .DIN1(n35798), .DIN2(wb_addr_i[23]), .Q(n35806) );
  and2s1 U28379 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[21]), .Q(n35804) );
  or2s1 U28380 ( .DIN1(n35808), .DIN2(n35809), .Q(n9137) );
  or2s1 U28381 ( .DIN1(n35810), .DIN2(n35811), .Q(n35809) );
  and2s1 U28382 ( .DIN1(n35797), .DIN2(n32549), .Q(n35811) );
  hi1s1 U28383 ( .DIN1(n36667), .Q(n32549) );
  and2s1 U28384 ( .DIN1(n35798), .DIN2(wb_addr_i[22]), .Q(n35810) );
  and2s1 U28385 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[20]), .Q(n35808) );
  or2s1 U28386 ( .DIN1(n35812), .DIN2(n35813), .Q(n9136) );
  or2s1 U28387 ( .DIN1(n35814), .DIN2(n35815), .Q(n35813) );
  and2s1 U28388 ( .DIN1(n35797), .DIN2(n32552), .Q(n35815) );
  hi1s1 U28389 ( .DIN1(n36668), .Q(n32552) );
  and2s1 U28390 ( .DIN1(n35798), .DIN2(wb_addr_i[21]), .Q(n35814) );
  and2s1 U28391 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[19]), .Q(n35812) );
  or2s1 U28392 ( .DIN1(n35816), .DIN2(n35817), .Q(n9135) );
  or2s1 U28393 ( .DIN1(n35818), .DIN2(n35819), .Q(n35817) );
  and2s1 U28394 ( .DIN1(n35797), .DIN2(n32555), .Q(n35819) );
  hi1s1 U28395 ( .DIN1(n36669), .Q(n32555) );
  and2s1 U28396 ( .DIN1(n35798), .DIN2(wb_addr_i[20]), .Q(n35818) );
  and2s1 U28397 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[18]), .Q(n35816) );
  or2s1 U28398 ( .DIN1(n35820), .DIN2(n35821), .Q(n9134) );
  or2s1 U28399 ( .DIN1(n35822), .DIN2(n35823), .Q(n35821) );
  and2s1 U28400 ( .DIN1(n35797), .DIN2(n32558), .Q(n35823) );
  hi1s1 U28401 ( .DIN1(n36670), .Q(n32558) );
  and2s1 U28402 ( .DIN1(n35798), .DIN2(wb_addr_i[19]), .Q(n35822) );
  and2s1 U28403 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[17]), .Q(n35820) );
  or2s1 U28404 ( .DIN1(n35824), .DIN2(n35825), .Q(n9133) );
  or2s1 U28405 ( .DIN1(n35826), .DIN2(n35827), .Q(n35825) );
  and2s1 U28406 ( .DIN1(n35797), .DIN2(n32561), .Q(n35827) );
  hi1s1 U28407 ( .DIN1(n36671), .Q(n32561) );
  and2s1 U28408 ( .DIN1(n35798), .DIN2(wb_addr_i[18]), .Q(n35826) );
  and2s1 U28409 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[16]), .Q(n35824) );
  or2s1 U28410 ( .DIN1(n35828), .DIN2(n35829), .Q(n9132) );
  or2s1 U28411 ( .DIN1(n35830), .DIN2(n35831), .Q(n35829) );
  and2s1 U28412 ( .DIN1(n35797), .DIN2(n32564), .Q(n35831) );
  hi1s1 U28413 ( .DIN1(n36672), .Q(n32564) );
  and2s1 U28414 ( .DIN1(n35798), .DIN2(wb_addr_i[17]), .Q(n35830) );
  and2s1 U28415 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[15]), .Q(n35828) );
  or2s1 U28416 ( .DIN1(n35832), .DIN2(n35833), .Q(n9131) );
  or2s1 U28417 ( .DIN1(n35834), .DIN2(n35835), .Q(n35833) );
  and2s1 U28418 ( .DIN1(n35836), .DIN2(n35096), .Q(n35835) );
  hi1s1 U28419 ( .DIN1(n36673), .Q(n35096) );
  and2s1 U28420 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[14]), .Q(n35834) );
  or2s1 U28421 ( .DIN1(n35837), .DIN2(n35838), .Q(n35832) );
  and2s1 U28422 ( .DIN1(n35797), .DIN2(n32567), .Q(n35838) );
  hi1s1 U28423 ( .DIN1(n36674), .Q(n32567) );
  and2s1 U28424 ( .DIN1(n35798), .DIN2(wb_addr_i[16]), .Q(n35837) );
  or2s1 U28425 ( .DIN1(n35839), .DIN2(n35840), .Q(n9130) );
  or2s1 U28426 ( .DIN1(n35841), .DIN2(n35842), .Q(n35840) );
  and2s1 U28427 ( .DIN1(n35836), .DIN2(n35084), .Q(n35842) );
  hi1s1 U28428 ( .DIN1(n36675), .Q(n35084) );
  and2s1 U28429 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[13]), .Q(n35841) );
  or2s1 U28430 ( .DIN1(n35843), .DIN2(n35844), .Q(n35839) );
  and2s1 U28431 ( .DIN1(n35797), .DIN2(n32570), .Q(n35844) );
  hi1s1 U28432 ( .DIN1(n36676), .Q(n32570) );
  and2s1 U28433 ( .DIN1(n35798), .DIN2(wb_addr_i[15]), .Q(n35843) );
  or2s1 U28434 ( .DIN1(n35845), .DIN2(n35846), .Q(n9129) );
  or2s1 U28435 ( .DIN1(n35847), .DIN2(n35848), .Q(n35846) );
  and2s1 U28436 ( .DIN1(n35849), .DIN2(u0_sp_tms[12]), .Q(n35848) );
  and2s1 U28437 ( .DIN1(n35850), .DIN2(n35099), .Q(n35847) );
  hi1s1 U28438 ( .DIN1(n36678), .Q(n35099) );
  or2s1 U28439 ( .DIN1(n35851), .DIN2(n35852), .Q(n35845) );
  or2s1 U28440 ( .DIN1(n35853), .DIN2(n35854), .Q(n35852) );
  and2s1 U28441 ( .DIN1(n35797), .DIN2(n32573), .Q(n35854) );
  hi1s1 U28442 ( .DIN1(n36677), .Q(n32573) );
  and2s1 U28443 ( .DIN1(n35798), .DIN2(wb_addr_i[14]), .Q(n35853) );
  and2s1 U28444 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[12]), .Q(n35851) );
  or2s1 U28445 ( .DIN1(n35855), .DIN2(n35856), .Q(n9128) );
  or2s1 U28446 ( .DIN1(n35857), .DIN2(n35858), .Q(n35856) );
  and2s1 U28447 ( .DIN1(n35849), .DIN2(u0_sp_tms[11]), .Q(n35858) );
  and2s1 U28448 ( .DIN1(n35850), .DIN2(n35128), .Q(n35857) );
  hi1s1 U28449 ( .DIN1(n36680), .Q(n35128) );
  or2s1 U28450 ( .DIN1(n35859), .DIN2(n35860), .Q(n35855) );
  or2s1 U28451 ( .DIN1(n35861), .DIN2(n35862), .Q(n35860) );
  and2s1 U28452 ( .DIN1(n35797), .DIN2(n32576), .Q(n35862) );
  hi1s1 U28453 ( .DIN1(n36679), .Q(n32576) );
  and2s1 U28454 ( .DIN1(n35798), .DIN2(wb_addr_i[13]), .Q(n35861) );
  and2s1 U28455 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[11]), .Q(n35859) );
  or2s1 U28456 ( .DIN1(n35863), .DIN2(n35864), .Q(n9127) );
  or2s1 U28457 ( .DIN1(n35865), .DIN2(n35866), .Q(n35864) );
  or2s1 U28458 ( .DIN1(n35867), .DIN2(n35868), .Q(n35866) );
  and2s1 U28459 ( .DIN1(n35850), .DIN2(n35142), .Q(n35868) );
  hi1s1 U28460 ( .DIN1(n36682), .Q(n35142) );
  and2s1 U28461 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[10]), .Q(n35867) );
  and2s1 U28462 ( .DIN1(n35849), .DIN2(u0_sp_tms[10]), .Q(n35865) );
  or2s1 U28463 ( .DIN1(n35869), .DIN2(n35870), .Q(n35863) );
  or2s1 U28464 ( .DIN1(n35871), .DIN2(n35872), .Q(n35870) );
  and2s1 U28465 ( .DIN1(n35797), .DIN2(n32579), .Q(n35872) );
  hi1s1 U28466 ( .DIN1(n36681), .Q(n32579) );
  and2s1 U28467 ( .DIN1(n35798), .DIN2(wb_addr_i[12]), .Q(n35871) );
  or2s1 U28468 ( .DIN1(rfr_ack), .DIN2(n35873), .Q(n35869) );
  and2s1 U28469 ( .DIN1(n35874), .DIN2(n35786), .Q(n35873) );
  or2s1 U28470 ( .DIN1(n35875), .DIN2(n35876), .Q(n35786) );
  or2s1 U28471 ( .DIN1(n35877), .DIN2(n35878), .Q(n35876) );
  and2s1 U28472 ( .DIN1(u5_ap_en), .DIN2(n35879), .Q(n35877) );
  or2s1 U28473 ( .DIN1(n32861), .DIN2(n35880), .Q(n35879) );
  or2s1 U28474 ( .DIN1(n35881), .DIN2(n32901), .Q(n35880) );
  or2s1 U28475 ( .DIN1(n35656), .DIN2(n33012), .Q(n32861) );
  or2s1 U28476 ( .DIN1(n35882), .DIN2(n35883), .Q(n33012) );
  or2s1 U28477 ( .DIN1(n32907), .DIN2(n35884), .Q(n35883) );
  or2s1 U28478 ( .DIN1(n35885), .DIN2(n34347), .Q(n35884) );
  or2s1 U28479 ( .DIN1(n35886), .DIN2(n35887), .Q(n35882) );
  or2s1 U28480 ( .DIN1(n33492), .DIN2(n34574), .Q(n35887) );
  or2s1 U28481 ( .DIN1(n35888), .DIN2(n35889), .Q(n35875) );
  or2s1 U28482 ( .DIN1(n34136), .DIN2(n35890), .Q(n35889) );
  and2s1 U28483 ( .DIN1(n35891), .DIN2(n32962), .Q(n35890) );
  and2s1 U28484 ( .DIN1(n34570), .DIN2(n32907), .Q(n35891) );
  and2s1 U28485 ( .DIN1(n35892), .DIN2(n4535), .Q(n35888) );
  or2s1 U28486 ( .DIN1(n34545), .DIN2(n35893), .Q(n35892) );
  or2s1 U28487 ( .DIN1(n35894), .DIN2(n35895), .Q(n9126) );
  or2s1 U28488 ( .DIN1(n35896), .DIN2(n35897), .Q(n35895) );
  or2s1 U28489 ( .DIN1(n35898), .DIN2(n35899), .Q(n35897) );
  and2s1 U28490 ( .DIN1(n35874), .DIN2(n35363), .Q(n35899) );
  hi1s1 U28491 ( .DIN1(n36685), .Q(n35363) );
  and2s1 U28492 ( .DIN1(n35850), .DIN2(n35155), .Q(n35898) );
  hi1s1 U28493 ( .DIN1(n36684), .Q(n35155) );
  and2s1 U28494 ( .DIN1(n35849), .DIN2(n35439), .Q(n35896) );
  or2s1 U28495 ( .DIN1(n35900), .DIN2(n35901), .Q(n35894) );
  or2s1 U28496 ( .DIN1(n35902), .DIN2(n35903), .Q(n35901) );
  and2s1 U28497 ( .DIN1(n35797), .DIN2(n32582), .Q(n35903) );
  hi1s1 U28498 ( .DIN1(n36683), .Q(n32582) );
  and2s1 U28499 ( .DIN1(n35798), .DIN2(wb_addr_i[11]), .Q(n35902) );
  and2s1 U28500 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[9]), .Q(n35900) );
  or2s1 U28501 ( .DIN1(n35904), .DIN2(n35905), .Q(n9125) );
  or2s1 U28502 ( .DIN1(n35906), .DIN2(n35907), .Q(n35905) );
  or2s1 U28503 ( .DIN1(n35908), .DIN2(n35909), .Q(n35907) );
  and2s1 U28504 ( .DIN1(n35874), .DIN2(n35356), .Q(n35909) );
  hi1s1 U28505 ( .DIN1(n36688), .Q(n35356) );
  and2s1 U28506 ( .DIN1(n35850), .DIN2(n35168), .Q(n35908) );
  hi1s1 U28507 ( .DIN1(n36687), .Q(n35168) );
  and2s1 U28508 ( .DIN1(n35849), .DIN2(u0_sp_tms[8]), .Q(n35906) );
  or2s1 U28509 ( .DIN1(n35910), .DIN2(n35911), .Q(n35904) );
  or2s1 U28510 ( .DIN1(n35912), .DIN2(n35913), .Q(n35911) );
  and2s1 U28511 ( .DIN1(n35797), .DIN2(n32585), .Q(n35913) );
  hi1s1 U28512 ( .DIN1(n36686), .Q(n32585) );
  and2s1 U28513 ( .DIN1(n35798), .DIN2(wb_addr_i[10]), .Q(n35912) );
  and2s1 U28514 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[8]), .Q(n35910) );
  or2s1 U28515 ( .DIN1(n35914), .DIN2(n35915), .Q(n9124) );
  or2s1 U28516 ( .DIN1(n35916), .DIN2(n35917), .Q(n35915) );
  or2s1 U28517 ( .DIN1(n35918), .DIN2(n35919), .Q(n35917) );
  and2s1 U28518 ( .DIN1(n35874), .DIN2(n35353), .Q(n35919) );
  hi1s1 U28519 ( .DIN1(n36691), .Q(n35353) );
  and2s1 U28520 ( .DIN1(n35850), .DIN2(n35180), .Q(n35918) );
  hi1s1 U28521 ( .DIN1(n36690), .Q(n35180) );
  and2s1 U28522 ( .DIN1(n35849), .DIN2(u0_sp_tms[7]), .Q(n35916) );
  or2s1 U28523 ( .DIN1(n35920), .DIN2(n35921), .Q(n35914) );
  or2s1 U28524 ( .DIN1(n35922), .DIN2(n35923), .Q(n35921) );
  and2s1 U28525 ( .DIN1(n35797), .DIN2(n32588), .Q(n35923) );
  hi1s1 U28526 ( .DIN1(n36689), .Q(n32588) );
  and2s1 U28527 ( .DIN1(n35798), .DIN2(wb_addr_i[9]), .Q(n35922) );
  and2s1 U28528 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[7]), .Q(n35920) );
  or2s1 U28529 ( .DIN1(n35924), .DIN2(n35925), .Q(n9123) );
  or2s1 U28530 ( .DIN1(n35926), .DIN2(n35927), .Q(n35925) );
  or2s1 U28531 ( .DIN1(n35928), .DIN2(n35929), .Q(n35927) );
  and2s1 U28532 ( .DIN1(n35874), .DIN2(n35350), .Q(n35929) );
  hi1s1 U28533 ( .DIN1(n36694), .Q(n35350) );
  and2s1 U28534 ( .DIN1(n35850), .DIN2(n35190), .Q(n35928) );
  hi1s1 U28535 ( .DIN1(n36693), .Q(n35190) );
  and2s1 U28536 ( .DIN1(n35849), .DIN2(u0_sp_tms[6]), .Q(n35926) );
  or2s1 U28537 ( .DIN1(n35930), .DIN2(n35931), .Q(n35924) );
  or2s1 U28538 ( .DIN1(n35932), .DIN2(n35933), .Q(n35931) );
  and2s1 U28539 ( .DIN1(n35797), .DIN2(n32591), .Q(n35933) );
  hi1s1 U28540 ( .DIN1(n36692), .Q(n32591) );
  and2s1 U28541 ( .DIN1(n35798), .DIN2(wb_addr_i[8]), .Q(n35932) );
  and2s1 U28542 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[6]), .Q(n35930) );
  or2s1 U28543 ( .DIN1(n35934), .DIN2(n35935), .Q(n9122) );
  or2s1 U28544 ( .DIN1(n35936), .DIN2(n35937), .Q(n35935) );
  or2s1 U28545 ( .DIN1(n35938), .DIN2(n35939), .Q(n35937) );
  and2s1 U28546 ( .DIN1(n35874), .DIN2(n35347), .Q(n35939) );
  hi1s1 U28547 ( .DIN1(n36697), .Q(n35347) );
  and2s1 U28548 ( .DIN1(n35850), .DIN2(n35200), .Q(n35938) );
  hi1s1 U28549 ( .DIN1(n36696), .Q(n35200) );
  and2s1 U28550 ( .DIN1(n35849), .DIN2(u0_sp_tms[5]), .Q(n35936) );
  or2s1 U28551 ( .DIN1(n35940), .DIN2(n35941), .Q(n35934) );
  or2s1 U28552 ( .DIN1(n35942), .DIN2(n35943), .Q(n35941) );
  and2s1 U28553 ( .DIN1(n35797), .DIN2(n32594), .Q(n35943) );
  hi1s1 U28554 ( .DIN1(n36695), .Q(n32594) );
  and2s1 U28555 ( .DIN1(n35798), .DIN2(wb_addr_i[7]), .Q(n35942) );
  and2s1 U28556 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[5]), .Q(n35940) );
  or2s1 U28557 ( .DIN1(n35944), .DIN2(n35945), .Q(n9121) );
  or2s1 U28558 ( .DIN1(n35946), .DIN2(n35947), .Q(n35945) );
  or2s1 U28559 ( .DIN1(n35948), .DIN2(n35949), .Q(n35947) );
  and2s1 U28560 ( .DIN1(n35874), .DIN2(n35344), .Q(n35949) );
  hi1s1 U28561 ( .DIN1(n36700), .Q(n35344) );
  and2s1 U28562 ( .DIN1(n35850), .DIN2(n35210), .Q(n35948) );
  hi1s1 U28563 ( .DIN1(n36699), .Q(n35210) );
  and2s1 U28564 ( .DIN1(n35849), .DIN2(u0_sp_tms[4]), .Q(n35946) );
  or2s1 U28565 ( .DIN1(n35950), .DIN2(n35951), .Q(n35944) );
  or2s1 U28566 ( .DIN1(n35952), .DIN2(n35953), .Q(n35951) );
  and2s1 U28567 ( .DIN1(n35797), .DIN2(n32597), .Q(n35953) );
  hi1s1 U28568 ( .DIN1(n36698), .Q(n32597) );
  and2s1 U28569 ( .DIN1(n35798), .DIN2(wb_addr_i[6]), .Q(n35952) );
  and2s1 U28570 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[4]), .Q(n35950) );
  or2s1 U28571 ( .DIN1(n35954), .DIN2(n35955), .Q(n9120) );
  or2s1 U28572 ( .DIN1(n35956), .DIN2(n35957), .Q(n35955) );
  or2s1 U28573 ( .DIN1(n35958), .DIN2(n35959), .Q(n35957) );
  and2s1 U28574 ( .DIN1(n35874), .DIN2(n35341), .Q(n35959) );
  hi1s1 U28575 ( .DIN1(n36703), .Q(n35341) );
  and2s1 U28576 ( .DIN1(n35850), .DIN2(n35220), .Q(n35958) );
  hi1s1 U28577 ( .DIN1(n36702), .Q(n35220) );
  and2s1 U28578 ( .DIN1(n35849), .DIN2(u0_sp_tms[3]), .Q(n35956) );
  or2s1 U28579 ( .DIN1(n35960), .DIN2(n35961), .Q(n35954) );
  or2s1 U28580 ( .DIN1(n35962), .DIN2(n35963), .Q(n35961) );
  and2s1 U28581 ( .DIN1(n35797), .DIN2(n32600), .Q(n35963) );
  hi1s1 U28582 ( .DIN1(n36701), .Q(n32600) );
  and2s1 U28583 ( .DIN1(n35798), .DIN2(wb_addr_i[5]), .Q(n35962) );
  and2s1 U28584 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[3]), .Q(n35960) );
  or2s1 U28585 ( .DIN1(n35964), .DIN2(n35965), .Q(n9119) );
  or2s1 U28586 ( .DIN1(n35966), .DIN2(n35967), .Q(n35965) );
  or2s1 U28587 ( .DIN1(n35968), .DIN2(n35969), .Q(n35967) );
  and2s1 U28588 ( .DIN1(n35874), .DIN2(n35338), .Q(n35969) );
  hi1s1 U28589 ( .DIN1(n36706), .Q(n35338) );
  and2s1 U28590 ( .DIN1(n35850), .DIN2(n35230), .Q(n35968) );
  hi1s1 U28591 ( .DIN1(n36705), .Q(n35230) );
  and2s1 U28592 ( .DIN1(n35849), .DIN2(n35970), .Q(n35966) );
  or2s1 U28593 ( .DIN1(n35971), .DIN2(n35972), .Q(n35964) );
  or2s1 U28594 ( .DIN1(n35973), .DIN2(n35974), .Q(n35972) );
  and2s1 U28595 ( .DIN1(n35797), .DIN2(n32603), .Q(n35974) );
  hi1s1 U28596 ( .DIN1(n36704), .Q(n32603) );
  and2s1 U28597 ( .DIN1(n35798), .DIN2(wb_addr_i[4]), .Q(n35973) );
  and2s1 U28598 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[2]), .Q(n35971) );
  or2s1 U28599 ( .DIN1(n35975), .DIN2(n35976), .Q(n9118) );
  or2s1 U28600 ( .DIN1(n35977), .DIN2(n35978), .Q(n35976) );
  or2s1 U28601 ( .DIN1(n35979), .DIN2(n35980), .Q(n35978) );
  and2s1 U28602 ( .DIN1(n35874), .DIN2(n35335), .Q(n35980) );
  hi1s1 U28603 ( .DIN1(n36709), .Q(n35335) );
  and2s1 U28604 ( .DIN1(n35850), .DIN2(n35246), .Q(n35979) );
  hi1s1 U28605 ( .DIN1(n36708), .Q(n35246) );
  and2s1 U28606 ( .DIN1(n35849), .DIN2(n35981), .Q(n35977) );
  or2s1 U28607 ( .DIN1(n35982), .DIN2(n35983), .Q(n35975) );
  or2s1 U28608 ( .DIN1(n35984), .DIN2(n35985), .Q(n35983) );
  and2s1 U28609 ( .DIN1(n35797), .DIN2(n32606), .Q(n35985) );
  hi1s1 U28610 ( .DIN1(n36707), .Q(n32606) );
  and2s1 U28611 ( .DIN1(n35798), .DIN2(wb_addr_i[3]), .Q(n35984) );
  and2s1 U28612 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[1]), .Q(n35982) );
  or2s1 U28613 ( .DIN1(n35986), .DIN2(n35987), .Q(n9117) );
  or2s1 U28614 ( .DIN1(n35988), .DIN2(n35989), .Q(n35987) );
  or2s1 U28615 ( .DIN1(n35990), .DIN2(n35991), .Q(n35989) );
  and2s1 U28616 ( .DIN1(n35874), .DIN2(n35331), .Q(n35991) );
  hi1s1 U28617 ( .DIN1(n36712), .Q(n35331) );
  hi1s1 U28618 ( .DIN1(n35992), .Q(n35874) );
  or2s1 U28619 ( .DIN1(n35993), .DIN2(n35994), .Q(n35992) );
  or2s1 U28620 ( .DIN1(n35995), .DIN2(n35996), .Q(n35994) );
  and2s1 U28621 ( .DIN1(n35850), .DIN2(n35284), .Q(n35990) );
  hi1s1 U28622 ( .DIN1(n36711), .Q(n35284) );
  and2s1 U28623 ( .DIN1(n35836), .DIN2(n35997), .Q(n35850) );
  and2s1 U28624 ( .DIN1(n35998), .DIN2(n35993), .Q(n35997) );
  or2s1 U28625 ( .DIN1(n33911), .DIN2(n32888), .Q(n35993) );
  and2s1 U28626 ( .DIN1(n35849), .DIN2(n35999), .Q(n35988) );
  and2s1 U28627 ( .DIN1(n35836), .DIN2(n35995), .Q(n35849) );
  hi1s1 U28628 ( .DIN1(n35998), .Q(n35995) );
  or2s1 U28629 ( .DIN1(\u5_temp_cs[1] ), .DIN2(n35283), .Q(n35998) );
  or2s1 U28630 ( .DIN1(n36000), .DIN2(n36001), .Q(\u5_temp_cs[1] ) );
  and2s1 U28631 ( .DIN1(n35054), .DIN2(n4531), .Q(n36001) );
  and2s1 U28632 ( .DIN1(n15502), .DIN2(n9180), .Q(n36000) );
  or2s1 U28633 ( .DIN1(n36002), .DIN2(n36003), .Q(n9180) );
  or2s1 U28634 ( .DIN1(n36004), .DIN2(n36005), .Q(n36003) );
  or2s1 U28635 ( .DIN1(n36006), .DIN2(n36007), .Q(n36005) );
  and2s1 U28636 ( .DIN1(n32943), .DIN2(n36008), .Q(n36006) );
  or2s1 U28637 ( .DIN1(n34136), .DIN2(n36009), .Q(n36002) );
  or2s1 U28638 ( .DIN1(n33901), .DIN2(n34536), .Q(n36009) );
  or2s1 U28639 ( .DIN1(n36010), .DIN2(n36011), .Q(n35986) );
  or2s1 U28640 ( .DIN1(n36012), .DIN2(n36013), .Q(n36011) );
  and2s1 U28641 ( .DIN1(n35797), .DIN2(n32609), .Q(n36013) );
  hi1s1 U28642 ( .DIN1(n36710), .Q(n32609) );
  and2s1 U28643 ( .DIN1(n35798), .DIN2(wb_addr_i[2]), .Q(n36012) );
  hi1s1 U28644 ( .DIN1(n36014), .Q(n35798) );
  or2s1 U28645 ( .DIN1(n35836), .DIN2(n36015), .Q(n36014) );
  or2s1 U28646 ( .DIN1(n35799), .DIN2(n35797), .Q(n36015) );
  hi1s1 U28647 ( .DIN1(n36016), .Q(n35797) );
  or2s1 U28648 ( .DIN1(n36017), .DIN2(n36018), .Q(n36016) );
  or2s1 U28649 ( .DIN1(n36019), .DIN2(n36020), .Q(n36018) );
  or2s1 U28650 ( .DIN1(n15514), .DIN2(n36021), .Q(n36017) );
  hi1s1 U28651 ( .DIN1(n35996), .Q(n35836) );
  or2s1 U28652 ( .DIN1(n36020), .DIN2(n36022), .Q(n35996) );
  or2s1 U28653 ( .DIN1(n36019), .DIN2(n36023), .Q(n36022) );
  and2s1 U28654 ( .DIN1(n35799), .DIN2(u1_u0_inc_in[0]), .Q(n36010) );
  and2s1 U28655 ( .DIN1(n36021), .DIN2(n36024), .Q(n35799) );
  and2s1 U28656 ( .DIN1(n36020), .DIN2(n36025), .Q(n36024) );
  hi1s1 U28657 ( .DIN1(n36019), .Q(n36025) );
  or2s1 U28658 ( .DIN1(n36026), .DIN2(n36027), .Q(n36019) );
  and2s1 U28659 ( .DIN1(u0_sp_csc[3]), .DIN2(n35282), .Q(n36027) );
  and2s1 U28660 ( .DIN1(u0_csc[3]), .DIN2(n35283), .Q(n36026) );
  or2s1 U28661 ( .DIN1(n36028), .DIN2(n36029), .Q(n36020) );
  and2s1 U28662 ( .DIN1(u0_sp_csc[2]), .DIN2(n35282), .Q(n36029) );
  and2s1 U28663 ( .DIN1(u0_csc[2]), .DIN2(n35283), .Q(n36028) );
  hi1s1 U28664 ( .DIN1(n36023), .Q(n36021) );
  or2s1 U28665 ( .DIN1(n36030), .DIN2(n36031), .Q(n36023) );
  and2s1 U28666 ( .DIN1(u0_sp_csc[1]), .DIN2(n35282), .Q(n36031) );
  and2s1 U28667 ( .DIN1(u0_csc[1]), .DIN2(n35283), .Q(n36030) );
  or2s1 U28668 ( .DIN1(n36032), .DIN2(n36033), .Q(n9116) );
  and2s1 U28669 ( .DIN1(wb_sel_i[3]), .DIN2(n32625), .Q(n36033) );
  and2s1 U28670 ( .DIN1(n32621), .DIN2(n9112), .Q(n36032) );
  or2s1 U28671 ( .DIN1(n36034), .DIN2(n36035), .Q(n9115) );
  and2s1 U28672 ( .DIN1(wb_sel_i[2]), .DIN2(n32625), .Q(n36035) );
  and2s1 U28673 ( .DIN1(n32621), .DIN2(n9111), .Q(n36034) );
  or2s1 U28674 ( .DIN1(n36036), .DIN2(n36037), .Q(n9114) );
  and2s1 U28675 ( .DIN1(wb_sel_i[1]), .DIN2(n32625), .Q(n36037) );
  and2s1 U28676 ( .DIN1(n32621), .DIN2(n9110), .Q(n36036) );
  or2s1 U28677 ( .DIN1(n36038), .DIN2(n36039), .Q(n9113) );
  and2s1 U28678 ( .DIN1(wb_sel_i[0]), .DIN2(n32625), .Q(n36039) );
  and2s1 U28679 ( .DIN1(n32621), .DIN2(n9109), .Q(n36038) );
  hi1s1 U28680 ( .DIN1(n32625), .Q(n32621) );
  and2s1 U28681 ( .DIN1(wb_cyc_i), .DIN2(wb_stb_i), .Q(n32625) );
  or2s1 U28682 ( .DIN1(n36040), .DIN2(n36041), .Q(n9108) );
  and2s1 U28683 ( .DIN1(n35792), .DIN2(n4993), .Q(n36040) );
  or2s1 U28684 ( .DIN1(n36042), .DIN2(n36041), .Q(n9107) );
  and2s1 U28685 ( .DIN1(n35792), .DIN2(n4994), .Q(n36042) );
  or2s1 U28686 ( .DIN1(n36043), .DIN2(n36041), .Q(n9106) );
  and2s1 U28687 ( .DIN1(n35792), .DIN2(n4995), .Q(n36043) );
  or2s1 U28688 ( .DIN1(n36044), .DIN2(n36041), .Q(n9105) );
  or2s1 U28689 ( .DIN1(n36045), .DIN2(u5_susp_sel_r), .Q(n36041) );
  and2s1 U28690 ( .DIN1(n15501), .DIN2(n36046), .Q(n36045) );
  or2s1 U28691 ( .DIN1(n32938), .DIN2(n35054), .Q(n36046) );
  hi1s1 U28692 ( .DIN1(u5_wb_cycle), .Q(n32938) );
  and2s1 U28693 ( .DIN1(n35792), .DIN2(n4996), .Q(n36044) );
  hi1s1 U28694 ( .DIN1(n15501), .Q(n35792) );
  or2s1 U28695 ( .DIN1(u5_susp_sel_r), .DIN2(n4533), .Q(n9104) );
  or2s1 U28696 ( .DIN1(n36047), .DIN2(n36048), .Q(n9103) );
  and2s1 U28697 ( .DIN1(n35054), .DIN2(n4532), .Q(n36048) );
  and2s1 U28698 ( .DIN1(n15502), .DIN2(n9182), .Q(n36047) );
  or2s1 U28699 ( .DIN1(n36049), .DIN2(n36050), .Q(n9182) );
  or2s1 U28700 ( .DIN1(n36051), .DIN2(n36052), .Q(n36050) );
  or2s1 U28701 ( .DIN1(n36053), .DIN2(n34347), .Q(n36052) );
  and2s1 U28702 ( .DIN1(n36054), .DIN2(n32943), .Q(n36053) );
  and2s1 U28703 ( .DIN1(n36055), .DIN2(n36008), .Q(n36054) );
  hi1s1 U28704 ( .DIN1(n36056), .Q(n36008) );
  or2s1 U28705 ( .DIN1(n36057), .DIN2(n36058), .Q(n36049) );
  or2s1 U28706 ( .DIN1(n34152), .DIN2(n34324), .Q(n36058) );
  or2s1 U28707 ( .DIN1(n35893), .DIN2(n33006), .Q(n36057) );
  and2s1 U28708 ( .DIN1(u5_tmr_done), .DIN2(n35598), .Q(n33006) );
  or2s1 U28709 ( .DIN1(n36059), .DIN2(n36060), .Q(n9102) );
  and2s1 U28710 ( .DIN1(n35054), .DIN2(n4530), .Q(n36060) );
  and2s1 U28711 ( .DIN1(n15502), .DIN2(n9184), .Q(n36059) );
  or2s1 U28712 ( .DIN1(n36061), .DIN2(n36062), .Q(n9184) );
  or2s1 U28713 ( .DIN1(n32907), .DIN2(n36004), .Q(n36062) );
  or2s1 U28714 ( .DIN1(n36063), .DIN2(n36064), .Q(n36004) );
  or2s1 U28715 ( .DIN1(n35599), .DIN2(n36051), .Q(n36064) );
  or2s1 U28716 ( .DIN1(n36065), .DIN2(n36066), .Q(n36051) );
  or2s1 U28717 ( .DIN1(n36067), .DIN2(n36068), .Q(n36066) );
  or2s1 U28718 ( .DIN1(n35881), .DIN2(n36069), .Q(n36068) );
  or2s1 U28719 ( .DIN1(n36070), .DIN2(n36071), .Q(n35881) );
  or2s1 U28720 ( .DIN1(n32869), .DIN2(n36072), .Q(n36071) );
  or2s1 U28721 ( .DIN1(n34273), .DIN2(n34274), .Q(n36070) );
  or2s1 U28722 ( .DIN1(n34117), .DIN2(n35885), .Q(n36067) );
  or2s1 U28723 ( .DIN1(n36073), .DIN2(n36074), .Q(n36065) );
  or2s1 U28724 ( .DIN1(n33896), .DIN2(n34574), .Q(n36074) );
  hi1s1 U28725 ( .DIN1(n36075), .Q(n34574) );
  or2s1 U28726 ( .DIN1(n32907), .DIN2(n36076), .Q(n36075) );
  or2s1 U28727 ( .DIN1(n35603), .DIN2(n34347), .Q(n36076) );
  or2s1 U28728 ( .DIN1(n34161), .DIN2(n35609), .Q(n34347) );
  or2s1 U28729 ( .DIN1(n34536), .DIN2(n32884), .Q(n35609) );
  or2s1 U28730 ( .DIN1(n36077), .DIN2(n36078), .Q(n35603) );
  or2s1 U28731 ( .DIN1(n33011), .DIN2(n35885), .Q(n36078) );
  or2s1 U28732 ( .DIN1(n36079), .DIN2(n36080), .Q(n35885) );
  or2s1 U28733 ( .DIN1(n36081), .DIN2(n36082), .Q(n36080) );
  or2s1 U28734 ( .DIN1(n33889), .DIN2(n36083), .Q(n36082) );
  or2s1 U28735 ( .DIN1(n35327), .DIN2(n34366), .Q(n36083) );
  or2s1 U28736 ( .DIN1(n36084), .DIN2(n34158), .Q(n34366) );
  and2s1 U28737 ( .DIN1(n36085), .DIN2(n36086), .Q(n34158) );
  hi1s1 U28738 ( .DIN1(n36087), .Q(n36085) );
  and2s1 U28739 ( .DIN1(n36088), .DIN2(n32928), .Q(n36084) );
  hi1s1 U28740 ( .DIN1(n36089), .Q(n32928) );
  and2s1 U28741 ( .DIN1(n32929), .DIN2(n36090), .Q(n36088) );
  hi1s1 U28742 ( .DIN1(n36091), .Q(n32929) );
  or2s1 U28743 ( .DIN1(n33910), .DIN2(n33911), .Q(n35327) );
  and2s1 U28744 ( .DIN1(u5_state[7]), .DIN2(n36092), .Q(n33911) );
  hi1s1 U28745 ( .DIN1(n36093), .Q(n36092) );
  or2s1 U28746 ( .DIN1(u5_state[9]), .DIN2(n36094), .Q(n36093) );
  and2s1 U28747 ( .DIN1(u5_state[8]), .DIN2(n36095), .Q(n33910) );
  hi1s1 U28748 ( .DIN1(n36096), .Q(n36095) );
  or2s1 U28749 ( .DIN1(u5_state[1]), .DIN2(n36097), .Q(n36096) );
  or2s1 U28750 ( .DIN1(n35393), .DIN2(n36098), .Q(n33889) );
  or2s1 U28751 ( .DIN1(n35388), .DIN2(n33879), .Q(n36098) );
  and2s1 U28752 ( .DIN1(u5_state[65]), .DIN2(n36099), .Q(n33879) );
  hi1s1 U28753 ( .DIN1(n36100), .Q(n36099) );
  or2s1 U28754 ( .DIN1(u5_state[63]), .DIN2(n36101), .Q(n36100) );
  hi1s1 U28755 ( .DIN1(n36102), .Q(n35388) );
  or2s1 U28756 ( .DIN1(n36103), .DIN2(n36104), .Q(n36102) );
  or2s1 U28757 ( .DIN1(n36105), .DIN2(n36106), .Q(n36104) );
  or2s1 U28758 ( .DIN1(n36107), .DIN2(n36108), .Q(n36106) );
  hi1s1 U28759 ( .DIN1(u5_state[51]), .Q(n36105) );
  or2s1 U28760 ( .DIN1(u5_state[57]), .DIN2(n36109), .Q(n36103) );
  and2s1 U28761 ( .DIN1(u5_state[40]), .DIN2(n36110), .Q(n35393) );
  and2s1 U28762 ( .DIN1(n36111), .DIN2(n36112), .Q(n36110) );
  or2s1 U28763 ( .DIN1(n33007), .DIN2(n36113), .Q(n36081) );
  or2s1 U28764 ( .DIN1(n34560), .DIN2(n34243), .Q(n36113) );
  hi1s1 U28765 ( .DIN1(n36114), .Q(n34243) );
  or2s1 U28766 ( .DIN1(n36115), .DIN2(n36116), .Q(n36114) );
  or2s1 U28767 ( .DIN1(n36117), .DIN2(n36118), .Q(n36116) );
  hi1s1 U28768 ( .DIN1(u5_state[21]), .Q(n36118) );
  or2s1 U28769 ( .DIN1(u5_state[22]), .DIN2(u5_state[18]), .Q(n36115) );
  hi1s1 U28770 ( .DIN1(n36119), .Q(n34560) );
  or2s1 U28771 ( .DIN1(n36120), .DIN2(n36121), .Q(n36119) );
  or2s1 U28772 ( .DIN1(n36122), .DIN2(n36123), .Q(n36121) );
  hi1s1 U28773 ( .DIN1(u5_state[3]), .Q(n36123) );
  or2s1 U28774 ( .DIN1(u5_state[37]), .DIN2(n36124), .Q(n36120) );
  hi1s1 U28775 ( .DIN1(n36125), .Q(n33007) );
  or2s1 U28776 ( .DIN1(n36126), .DIN2(n36127), .Q(n36125) );
  or2s1 U28777 ( .DIN1(n36128), .DIN2(n36129), .Q(n36127) );
  hi1s1 U28778 ( .DIN1(u5_state[62]), .Q(n36129) );
  or2s1 U28779 ( .DIN1(u5_state[5]), .DIN2(u5_state[57]), .Q(n36126) );
  or2s1 U28780 ( .DIN1(n36130), .DIN2(n36131), .Q(n36079) );
  or2s1 U28781 ( .DIN1(n32960), .DIN2(n36132), .Q(n36131) );
  or2s1 U28782 ( .DIN1(n34125), .DIN2(n33487), .Q(n36132) );
  hi1s1 U28783 ( .DIN1(n36133), .Q(n32960) );
  or2s1 U28784 ( .DIN1(n36134), .DIN2(n36135), .Q(n36133) );
  or2s1 U28785 ( .DIN1(n36136), .DIN2(n36137), .Q(n36135) );
  hi1s1 U28786 ( .DIN1(u5_state[12]), .Q(n36137) );
  or2s1 U28787 ( .DIN1(u5_state[13]), .DIN2(n36138), .Q(n36134) );
  or2s1 U28788 ( .DIN1(n33871), .DIN2(n36139), .Q(n36130) );
  or2s1 U28789 ( .DIN1(n34544), .DIN2(n32858), .Q(n36139) );
  hi1s1 U28790 ( .DIN1(n36140), .Q(n34544) );
  or2s1 U28791 ( .DIN1(n36141), .DIN2(n36142), .Q(n36140) );
  or2s1 U28792 ( .DIN1(n36143), .DIN2(n36144), .Q(n36142) );
  hi1s1 U28793 ( .DIN1(u5_state[0]), .Q(n36144) );
  or2s1 U28794 ( .DIN1(n32864), .DIN2(n36072), .Q(n33011) );
  or2s1 U28795 ( .DIN1(n36145), .DIN2(n36146), .Q(n36072) );
  or2s1 U28796 ( .DIN1(n32865), .DIN2(n32868), .Q(n36146) );
  hi1s1 U28797 ( .DIN1(n36147), .Q(n32868) );
  or2s1 U28798 ( .DIN1(n36148), .DIN2(n36149), .Q(n36147) );
  or2s1 U28799 ( .DIN1(n36150), .DIN2(n36151), .Q(n36149) );
  hi1s1 U28800 ( .DIN1(u5_state[19]), .Q(n36151) );
  or2s1 U28801 ( .DIN1(u5_state[17]), .DIN2(u5_state[16]), .Q(n36148) );
  hi1s1 U28802 ( .DIN1(n36152), .Q(n32865) );
  or2s1 U28803 ( .DIN1(n36153), .DIN2(n36154), .Q(n36152) );
  or2s1 U28804 ( .DIN1(n36155), .DIN2(n36156), .Q(n36154) );
  or2s1 U28805 ( .DIN1(u5_state[34]), .DIN2(u5_state[27]), .Q(n36153) );
  or2s1 U28806 ( .DIN1(n34263), .DIN2(n36157), .Q(n36145) );
  or2s1 U28807 ( .DIN1(n34261), .DIN2(n32870), .Q(n36157) );
  and2s1 U28808 ( .DIN1(u5_state[33]), .DIN2(n36158), .Q(n34261) );
  hi1s1 U28809 ( .DIN1(n36159), .Q(n36158) );
  or2s1 U28810 ( .DIN1(u5_state[39]), .DIN2(n36160), .Q(n36159) );
  hi1s1 U28811 ( .DIN1(n36161), .Q(n34263) );
  or2s1 U28812 ( .DIN1(n36162), .DIN2(n36163), .Q(n36161) );
  or2s1 U28813 ( .DIN1(n36164), .DIN2(n36155), .Q(n36163) );
  or2s1 U28814 ( .DIN1(n36165), .DIN2(n36166), .Q(n32864) );
  or2s1 U28815 ( .DIN1(n36007), .DIN2(n36167), .Q(n36166) );
  or2s1 U28816 ( .DIN1(n34324), .DIN2(n34290), .Q(n36167) );
  or2s1 U28817 ( .DIN1(n34545), .DIN2(n36168), .Q(n36165) );
  or2s1 U28818 ( .DIN1(u5_init_ack), .DIN2(n33901), .Q(n36168) );
  or2s1 U28819 ( .DIN1(n35886), .DIN2(n36169), .Q(n36077) );
  or2s1 U28820 ( .DIN1(u5_suspended_d), .DIN2(n32869), .Q(n36169) );
  hi1s1 U28821 ( .DIN1(n36170), .Q(n32869) );
  or2s1 U28822 ( .DIN1(n36171), .DIN2(n36172), .Q(n36170) );
  or2s1 U28823 ( .DIN1(n36089), .DIN2(n36090), .Q(n36172) );
  hi1s1 U28824 ( .DIN1(u5_state[11]), .Q(n36090) );
  or2s1 U28825 ( .DIN1(u5_state[10]), .DIN2(n36091), .Q(n36171) );
  or2s1 U28826 ( .DIN1(n36173), .DIN2(n36174), .Q(n35886) );
  or2s1 U28827 ( .DIN1(n36175), .DIN2(n36176), .Q(n36174) );
  or2s1 U28828 ( .DIN1(n34584), .DIN2(n36177), .Q(n36173) );
  hi1s1 U28829 ( .DIN1(n9092), .Q(n34584) );
  or2s1 U28830 ( .DIN1(n34116), .DIN2(n36178), .Q(n36073) );
  or2s1 U28831 ( .DIN1(u5_suspended_d), .DIN2(n34545), .Q(n36178) );
  hi1s1 U28832 ( .DIN1(n36179), .Q(n34545) );
  or2s1 U28833 ( .DIN1(n36180), .DIN2(n36181), .Q(n36179) );
  or2s1 U28834 ( .DIN1(n36182), .DIN2(n36183), .Q(n36181) );
  hi1s1 U28835 ( .DIN1(u5_state[2]), .Q(n36183) );
  or2s1 U28836 ( .DIN1(n33492), .DIN2(n35656), .Q(u5_suspended_d) );
  or2s1 U28837 ( .DIN1(n34257), .DIN2(n33013), .Q(n35656) );
  hi1s1 U28838 ( .DIN1(n36184), .Q(n33013) );
  or2s1 U28839 ( .DIN1(n36185), .DIN2(n36186), .Q(n36184) );
  or2s1 U28840 ( .DIN1(n36182), .DIN2(n36187), .Q(n36186) );
  hi1s1 U28841 ( .DIN1(u5_state[31]), .Q(n36187) );
  or2s1 U28842 ( .DIN1(u5_state[30]), .DIN2(u5_state[2]), .Q(n36185) );
  hi1s1 U28843 ( .DIN1(n34343), .Q(n34257) );
  or2s1 U28844 ( .DIN1(n36188), .DIN2(n36189), .Q(n34343) );
  or2s1 U28845 ( .DIN1(n36182), .DIN2(n36190), .Q(n36189) );
  hi1s1 U28846 ( .DIN1(u5_state[30]), .Q(n36190) );
  or2s1 U28847 ( .DIN1(n36191), .DIN2(n36192), .Q(n36182) );
  or2s1 U28848 ( .DIN1(n36193), .DIN2(n36194), .Q(n36192) );
  or2s1 U28849 ( .DIN1(u5_state[29]), .DIN2(n36195), .Q(n36191) );
  or2s1 U28850 ( .DIN1(u5_state[31]), .DIN2(u5_state[2]), .Q(n36188) );
  hi1s1 U28851 ( .DIN1(n36196), .Q(n33492) );
  or2s1 U28852 ( .DIN1(n36197), .DIN2(n36198), .Q(n36196) );
  or2s1 U28853 ( .DIN1(n36194), .DIN2(n36199), .Q(n36198) );
  hi1s1 U28854 ( .DIN1(u5_state[32]), .Q(n36199) );
  or2s1 U28855 ( .DIN1(n36200), .DIN2(n36201), .Q(n36197) );
  or2s1 U28856 ( .DIN1(n36202), .DIN2(n36203), .Q(n36201) );
  and2s1 U28857 ( .DIN1(u5_state[54]), .DIN2(n36204), .Q(n34116) );
  and2s1 U28858 ( .DIN1(n36205), .DIN2(n36206), .Q(n36204) );
  or2s1 U28859 ( .DIN1(n34121), .DIN2(n36177), .Q(n36063) );
  or2s1 U28860 ( .DIN1(n35598), .DIN2(n32967), .Q(n36177) );
  or2s1 U28861 ( .DIN1(n32943), .DIN2(n32940), .Q(n32907) );
  or2s1 U28862 ( .DIN1(n36207), .DIN2(n36208), .Q(n36061) );
  or2s1 U28863 ( .DIN1(n32884), .DIN2(n35893), .Q(n36208) );
  and2s1 U28864 ( .DIN1(n36209), .DIN2(n33901), .Q(n35893) );
  or2s1 U28865 ( .DIN1(n34363), .DIN2(n33902), .Q(n36209) );
  and2s1 U28866 ( .DIN1(n34536), .DIN2(u5_wb_wait_r), .Q(n36207) );
  or2s1 U28867 ( .DIN1(n36210), .DIN2(n36211), .Q(n9101) );
  or2s1 U28868 ( .DIN1(n36212), .DIN2(n36213), .Q(n36211) );
  and2s1 U28869 ( .DIN1(n36214), .DIN2(n33954), .Q(n36213) );
  or2s1 U28870 ( .DIN1(n33754), .DIN2(n34310), .Q(n33954) );
  or2s1 U28871 ( .DIN1(n32750), .DIN2(n36215), .Q(n34310) );
  or2s1 U28872 ( .DIN1(u0_csc0[3]), .DIN2(u0_csc0[2]), .Q(n36215) );
  hi1s1 U28873 ( .DIN1(u0_csc0[0]), .Q(n33754) );
  and2s1 U28874 ( .DIN1(n36216), .DIN2(n36217), .Q(n36212) );
  or2s1 U28875 ( .DIN1(n36218), .DIN2(n36219), .Q(n36217) );
  and2s1 U28876 ( .DIN1(n35282), .DIN2(n33952), .Q(n36219) );
  hi1s1 U28877 ( .DIN1(u0_spec_req_cs[0]), .Q(n33952) );
  hi1s1 U28878 ( .DIN1(n36220), .Q(n36218) );
  or2s1 U28879 ( .DIN1(n35282), .DIN2(u0_cs[0]), .Q(n36220) );
  or2s1 U28880 ( .DIN1(n36210), .DIN2(n36221), .Q(n9100) );
  or2s1 U28881 ( .DIN1(n36222), .DIN2(n36223), .Q(n36221) );
  and2s1 U28882 ( .DIN1(n36214), .DIN2(n33939), .Q(n36223) );
  or2s1 U28883 ( .DIN1(n33812), .DIN2(n34303), .Q(n33939) );
  or2s1 U28884 ( .DIN1(n32426), .DIN2(n36224), .Q(n34303) );
  or2s1 U28885 ( .DIN1(u0_csc1[3]), .DIN2(u0_csc1[2]), .Q(n36224) );
  hi1s1 U28886 ( .DIN1(u0_csc1[0]), .Q(n33812) );
  and2s1 U28887 ( .DIN1(n36216), .DIN2(n36225), .Q(n36222) );
  or2s1 U28888 ( .DIN1(n36226), .DIN2(n36227), .Q(n36225) );
  and2s1 U28889 ( .DIN1(n35282), .DIN2(n33937), .Q(n36227) );
  hi1s1 U28890 ( .DIN1(u0_spec_req_cs[1]), .Q(n33937) );
  hi1s1 U28891 ( .DIN1(n36228), .Q(n36226) );
  or2s1 U28892 ( .DIN1(n35282), .DIN2(u0_cs[1]), .Q(n36228) );
  or2s1 U28893 ( .DIN1(n36229), .DIN2(n36230), .Q(n9099) );
  or2s1 U28894 ( .DIN1(n36231), .DIN2(n36232), .Q(n36230) );
  and2s1 U28895 ( .DIN1(n15494), .DIN2(n35282), .Q(n36232) );
  and2s1 U28896 ( .DIN1(n15500), .DIN2(n35283), .Q(n36231) );
  or2s1 U28897 ( .DIN1(n36229), .DIN2(n36233), .Q(n9098) );
  or2s1 U28898 ( .DIN1(n36234), .DIN2(n36235), .Q(n36233) );
  and2s1 U28899 ( .DIN1(n15493), .DIN2(n35282), .Q(n36235) );
  and2s1 U28900 ( .DIN1(n15499), .DIN2(n35283), .Q(n36234) );
  or2s1 U28901 ( .DIN1(n36229), .DIN2(n36236), .Q(n9097) );
  or2s1 U28902 ( .DIN1(n36237), .DIN2(n36238), .Q(n36236) );
  and2s1 U28903 ( .DIN1(n15492), .DIN2(n35282), .Q(n36238) );
  and2s1 U28904 ( .DIN1(n15498), .DIN2(n35283), .Q(n36237) );
  or2s1 U28905 ( .DIN1(n36229), .DIN2(n36239), .Q(n9096) );
  or2s1 U28906 ( .DIN1(n36240), .DIN2(n36241), .Q(n36239) );
  and2s1 U28907 ( .DIN1(n15491), .DIN2(n35282), .Q(n36241) );
  and2s1 U28908 ( .DIN1(n15497), .DIN2(n35283), .Q(n36240) );
  or2s1 U28909 ( .DIN1(n36229), .DIN2(n36242), .Q(n9095) );
  or2s1 U28910 ( .DIN1(n36243), .DIN2(n36244), .Q(n36242) );
  and2s1 U28911 ( .DIN1(n15490), .DIN2(n35282), .Q(n36244) );
  and2s1 U28912 ( .DIN1(n15496), .DIN2(n35283), .Q(n36243) );
  or2s1 U28913 ( .DIN1(n36229), .DIN2(n36245), .Q(n9094) );
  or2s1 U28914 ( .DIN1(n36246), .DIN2(n36247), .Q(n36245) );
  and2s1 U28915 ( .DIN1(n15489), .DIN2(n35282), .Q(n36247) );
  and2s1 U28916 ( .DIN1(n15495), .DIN2(n35283), .Q(n36246) );
  or2s1 U28917 ( .DIN1(n36214), .DIN2(n36210), .Q(n36229) );
  or2s1 U28918 ( .DIN1(n36248), .DIN2(n36249), .Q(n36210) );
  and2s1 U28919 ( .DIN1(n35054), .DIN2(n4997), .Q(n36249) );
  hi1s1 U28920 ( .DIN1(n36250), .Q(n36248) );
  or2s1 U28921 ( .DIN1(n35054), .DIN2(n9682), .Q(n36250) );
  or2s1 U28922 ( .DIN1(n36251), .DIN2(n36252), .Q(n9682) );
  or2s1 U28923 ( .DIN1(n36253), .DIN2(n36254), .Q(n36252) );
  or2s1 U28924 ( .DIN1(n35784), .DIN2(n35597), .Q(n36254) );
  or2s1 U28925 ( .DIN1(n36255), .DIN2(n34121), .Q(n35597) );
  and2s1 U28926 ( .DIN1(n33487), .DIN2(n36256), .Q(n36255) );
  or2s1 U28927 ( .DIN1(n36257), .DIN2(n36258), .Q(n36256) );
  or2s1 U28928 ( .DIN1(n35411), .DIN2(n32889), .Q(n36258) );
  or2s1 U28929 ( .DIN1(n35415), .DIN2(n36259), .Q(n32889) );
  or2s1 U28930 ( .DIN1(n36260), .DIN2(n36261), .Q(n36259) );
  and2s1 U28931 ( .DIN1(u0_sp_tms[18]), .DIN2(n35282), .Q(n36261) );
  and2s1 U28932 ( .DIN1(u0_tms[18]), .DIN2(n35283), .Q(n36260) );
  or2s1 U28933 ( .DIN1(n35415), .DIN2(n36262), .Q(n35411) );
  or2s1 U28934 ( .DIN1(n36263), .DIN2(n36264), .Q(n36262) );
  and2s1 U28935 ( .DIN1(u0_sp_tms[17]), .DIN2(n35282), .Q(n36264) );
  and2s1 U28936 ( .DIN1(u0_tms[17]), .DIN2(n35283), .Q(n36263) );
  or2s1 U28937 ( .DIN1(n35390), .DIN2(n35456), .Q(n36257) );
  or2s1 U28938 ( .DIN1(n35415), .DIN2(n36265), .Q(n35456) );
  or2s1 U28939 ( .DIN1(n36266), .DIN2(n36267), .Q(n36265) );
  and2s1 U28940 ( .DIN1(u0_sp_tms[19]), .DIN2(n35282), .Q(n36267) );
  and2s1 U28941 ( .DIN1(u0_tms[19]), .DIN2(n35283), .Q(n36266) );
  or2s1 U28942 ( .DIN1(n35415), .DIN2(n36268), .Q(n35390) );
  or2s1 U28943 ( .DIN1(n36269), .DIN2(n36270), .Q(n36268) );
  and2s1 U28944 ( .DIN1(u0_sp_tms[16]), .DIN2(n35282), .Q(n36270) );
  and2s1 U28945 ( .DIN1(u0_tms[16]), .DIN2(n35283), .Q(n36269) );
  hi1s1 U28946 ( .DIN1(n36271), .Q(n33487) );
  or2s1 U28947 ( .DIN1(n36272), .DIN2(n36273), .Q(n36271) );
  or2s1 U28948 ( .DIN1(n36274), .DIN2(n36275), .Q(n36273) );
  hi1s1 U28949 ( .DIN1(u5_state[49]), .Q(n36275) );
  or2s1 U28950 ( .DIN1(u5_state[48]), .DIN2(u5_state[14]), .Q(n36272) );
  or2s1 U28951 ( .DIN1(n34352), .DIN2(n36276), .Q(n35784) );
  or2s1 U28952 ( .DIN1(n32888), .DIN2(n32884), .Q(n36276) );
  and2s1 U28953 ( .DIN1(u5_state[9]), .DIN2(n36277), .Q(n32884) );
  hi1s1 U28954 ( .DIN1(n36278), .Q(n36277) );
  or2s1 U28955 ( .DIN1(u5_state[7]), .DIN2(n36094), .Q(n36278) );
  or2s1 U28956 ( .DIN1(n36279), .DIN2(n36280), .Q(n36094) );
  and2s1 U28957 ( .DIN1(n33908), .DIN2(n34536), .Q(n32888) );
  and2s1 U28958 ( .DIN1(u5_state[6]), .DIN2(n36281), .Q(n34536) );
  hi1s1 U28959 ( .DIN1(n36282), .Q(n36281) );
  or2s1 U28960 ( .DIN1(u5_state[64]), .DIN2(n36283), .Q(n36282) );
  hi1s1 U28961 ( .DIN1(u5_wb_wait_r), .Q(n33908) );
  or2s1 U28962 ( .DIN1(n32887), .DIN2(n32901), .Q(n34352) );
  or2s1 U28963 ( .DIN1(n34152), .DIN2(n32990), .Q(n32901) );
  or2s1 U28964 ( .DIN1(n34290), .DIN2(n36284), .Q(n32990) );
  or2s1 U28965 ( .DIN1(n36285), .DIN2(n34324), .Q(n36284) );
  hi1s1 U28966 ( .DIN1(n36286), .Q(n34290) );
  or2s1 U28967 ( .DIN1(n36287), .DIN2(n36288), .Q(n36286) );
  or2s1 U28968 ( .DIN1(n36289), .DIN2(n36290), .Q(n36288) );
  hi1s1 U28969 ( .DIN1(u5_state[20]), .Q(n36290) );
  or2s1 U28970 ( .DIN1(n36291), .DIN2(n36292), .Q(n36287) );
  or2s1 U28971 ( .DIN1(u5_state[17]), .DIN2(n36091), .Q(n36292) );
  or2s1 U28972 ( .DIN1(n32967), .DIN2(n32966), .Q(n32887) );
  or2s1 U28973 ( .DIN1(n36007), .DIN2(n36293), .Q(n32966) );
  or2s1 U28974 ( .DIN1(n32992), .DIN2(n34136), .Q(n36293) );
  and2s1 U28975 ( .DIN1(u5_tmr_done), .DIN2(n36294), .Q(n32992) );
  and2s1 U28976 ( .DIN1(n32962), .DIN2(n33901), .Q(n36294) );
  hi1s1 U28977 ( .DIN1(n36295), .Q(n33901) );
  or2s1 U28978 ( .DIN1(n36296), .DIN2(n36297), .Q(n36295) );
  or2s1 U28979 ( .DIN1(n36150), .DIN2(n36298), .Q(n36297) );
  hi1s1 U28980 ( .DIN1(u5_state[16]), .Q(n36298) );
  or2s1 U28981 ( .DIN1(u5_state[19]), .DIN2(u5_state[17]), .Q(n36296) );
  hi1s1 U28982 ( .DIN1(n33902), .Q(n32962) );
  or2s1 U28983 ( .DIN1(n36299), .DIN2(n36300), .Q(n33902) );
  and2s1 U28984 ( .DIN1(u0_sp_csc_10), .DIN2(n35282), .Q(n36300) );
  and2s1 U28985 ( .DIN1(u0_csc_10), .DIN2(n35283), .Q(n36299) );
  or2s1 U28986 ( .DIN1(n34254), .DIN2(n35878), .Q(n36007) );
  or2s1 U28987 ( .DIN1(n36301), .DIN2(n34283), .Q(n35878) );
  and2s1 U28988 ( .DIN1(u5_state[18]), .DIN2(n36302), .Q(n34283) );
  hi1s1 U28989 ( .DIN1(n36303), .Q(n36302) );
  or2s1 U28990 ( .DIN1(n36304), .DIN2(n36117), .Q(n36303) );
  and2s1 U28991 ( .DIN1(n34266), .DIN2(n34268), .Q(n36301) );
  and2s1 U28992 ( .DIN1(n36162), .DIN2(n36156), .Q(n34268) );
  hi1s1 U28993 ( .DIN1(u5_state[35]), .Q(n36156) );
  hi1s1 U28994 ( .DIN1(u5_state[34]), .Q(n36162) );
  and2s1 U28995 ( .DIN1(u5_state[27]), .DIN2(n36305), .Q(n34266) );
  hi1s1 U28996 ( .DIN1(n36155), .Q(n36305) );
  or2s1 U28997 ( .DIN1(n36306), .DIN2(n36307), .Q(n36155) );
  or2s1 U28998 ( .DIN1(u5_state[60]), .DIN2(n36308), .Q(n36306) );
  hi1s1 U28999 ( .DIN1(n36309), .Q(n32967) );
  or2s1 U29000 ( .DIN1(n36310), .DIN2(n36311), .Q(n36309) );
  or2s1 U29001 ( .DIN1(n36312), .DIN2(n36313), .Q(n36311) );
  hi1s1 U29002 ( .DIN1(u5_state[15]), .Q(n36312) );
  or2s1 U29003 ( .DIN1(u5_state[18]), .DIN2(n36314), .Q(n36310) );
  or2s1 U29004 ( .DIN1(n36175), .DIN2(n36315), .Q(n36253) );
  or2s1 U29005 ( .DIN1(n36316), .DIN2(n34355), .Q(n36315) );
  and2s1 U29006 ( .DIN1(n35598), .DIN2(n34363), .Q(n34355) );
  hi1s1 U29007 ( .DIN1(u5_tmr_done), .Q(n34363) );
  and2s1 U29008 ( .DIN1(u5_state[64]), .DIN2(n36317), .Q(n35598) );
  hi1s1 U29009 ( .DIN1(n36318), .Q(n36317) );
  or2s1 U29010 ( .DIN1(u5_state[6]), .DIN2(n36283), .Q(n36318) );
  or2s1 U29011 ( .DIN1(n36319), .DIN2(n36320), .Q(n36283) );
  or2s1 U29012 ( .DIN1(u5_state[65]), .DIN2(u5_state[63]), .Q(n36320) );
  and2s1 U29013 ( .DIN1(n32943), .DIN2(n36321), .Q(n36316) );
  or2s1 U29014 ( .DIN1(n36056), .DIN2(n32942), .Q(n36321) );
  hi1s1 U29015 ( .DIN1(n36055), .Q(n32942) );
  or2s1 U29016 ( .DIN1(n34567), .DIN2(n34569), .Q(n36055) );
  or2s1 U29017 ( .DIN1(n34570), .DIN2(n36322), .Q(n34569) );
  or2s1 U29018 ( .DIN1(u5_wb_write_go_r), .DIN2(n32957), .Q(n36322) );
  or2s1 U29019 ( .DIN1(n34331), .DIN2(n33480), .Q(n32957) );
  hi1s1 U29020 ( .DIN1(n9537), .Q(n33480) );
  or2s1 U29021 ( .DIN1(n34966), .DIN2(n36323), .Q(n9537) );
  or2s1 U29022 ( .DIN1(u5_burst_cnt[9]), .DIN2(u5_burst_cnt[10]), .Q(n36323) );
  or2s1 U29023 ( .DIN1(n35021), .DIN2(n36324), .Q(n34966) );
  or2s1 U29024 ( .DIN1(u5_burst_cnt[8]), .DIN2(u5_burst_cnt[7]), .Q(n36324) );
  or2s1 U29025 ( .DIN1(n35005), .DIN2(n36325), .Q(n35021) );
  or2s1 U29026 ( .DIN1(u5_burst_cnt[6]), .DIN2(u5_burst_cnt[5]), .Q(n36325) );
  or2s1 U29027 ( .DIN1(n34990), .DIN2(n36326), .Q(n35005) );
  or2s1 U29028 ( .DIN1(u5_burst_cnt[4]), .DIN2(u5_burst_cnt[3]), .Q(n36326) );
  or2s1 U29029 ( .DIN1(u5_burst_cnt[2]), .DIN2(n34979), .Q(n34990) );
  or2s1 U29030 ( .DIN1(u5_burst_cnt[0]), .DIN2(u5_burst_cnt[1]), .Q(n34979) );
  hi1s1 U29031 ( .DIN1(n32956), .Q(n34567) );
  or2s1 U29032 ( .DIN1(n36327), .DIN2(u5_cke_r), .Q(n32956) );
  and2s1 U29033 ( .DIN1(n32941), .DIN2(n35052), .Q(n36327) );
  hi1s1 U29034 ( .DIN1(u5_cnt), .Q(n35052) );
  and2s1 U29035 ( .DIN1(n34570), .DIN2(u5_wb_cycle), .Q(n36056) );
  hi1s1 U29036 ( .DIN1(n32941), .Q(n34570) );
  and2s1 U29037 ( .DIN1(n36328), .DIN2(n36329), .Q(n32941) );
  hi1s1 U29038 ( .DIN1(n35439), .Q(n36329) );
  or2s1 U29039 ( .DIN1(n36330), .DIN2(n36331), .Q(n35439) );
  and2s1 U29040 ( .DIN1(u0_sp_tms[9]), .DIN2(n35282), .Q(n36331) );
  and2s1 U29041 ( .DIN1(u0_tms[9]), .DIN2(n35283), .Q(n36330) );
  or2s1 U29042 ( .DIN1(n36332), .DIN2(n35970), .Q(n36328) );
  or2s1 U29043 ( .DIN1(n35999), .DIN2(n35981), .Q(n36332) );
  hi1s1 U29044 ( .DIN1(n36333), .Q(n32943) );
  or2s1 U29045 ( .DIN1(n36334), .DIN2(n36335), .Q(n36333) );
  or2s1 U29046 ( .DIN1(n36274), .DIN2(n36336), .Q(n36335) );
  hi1s1 U29047 ( .DIN1(u5_state[14]), .Q(n36336) );
  or2s1 U29048 ( .DIN1(n35599), .DIN2(n36337), .Q(n36175) );
  or2s1 U29049 ( .DIN1(n34955), .DIN2(n36338), .Q(n36337) );
  or2s1 U29050 ( .DIN1(n34351), .DIN2(n36339), .Q(n35599) );
  or2s1 U29051 ( .DIN1(n34249), .DIN2(n32896), .Q(n36339) );
  and2s1 U29052 ( .DIN1(u5_state[63]), .DIN2(n36340), .Q(n32896) );
  hi1s1 U29053 ( .DIN1(n36341), .Q(n36340) );
  or2s1 U29054 ( .DIN1(u5_state[65]), .DIN2(n36101), .Q(n36341) );
  or2s1 U29055 ( .DIN1(n36319), .DIN2(n36342), .Q(n36101) );
  or2s1 U29056 ( .DIN1(u5_state[6]), .DIN2(u5_state[64]), .Q(n36342) );
  or2s1 U29057 ( .DIN1(n36343), .DIN2(n36344), .Q(n36319) );
  or2s1 U29058 ( .DIN1(n36345), .DIN2(n36346), .Q(n36344) );
  and2s1 U29059 ( .DIN1(n36347), .DIN2(n36348), .Q(n34249) );
  and2s1 U29060 ( .DIN1(n36349), .DIN2(u5_state[47]), .Q(n36348) );
  hi1s1 U29061 ( .DIN1(n36350), .Q(n36347) );
  or2s1 U29062 ( .DIN1(u5_state[46]), .DIN2(n36351), .Q(n36350) );
  hi1s1 U29063 ( .DIN1(n36352), .Q(n34351) );
  or2s1 U29064 ( .DIN1(n36353), .DIN2(n36354), .Q(n36352) );
  or2s1 U29065 ( .DIN1(n36274), .DIN2(n36355), .Q(n36354) );
  hi1s1 U29066 ( .DIN1(u5_state[48]), .Q(n36355) );
  or2s1 U29067 ( .DIN1(n36356), .DIN2(n36136), .Q(n36274) );
  or2s1 U29068 ( .DIN1(u5_state[49]), .DIN2(u5_state[14]), .Q(n36353) );
  or2s1 U29069 ( .DIN1(n36357), .DIN2(n36358), .Q(n36251) );
  or2s1 U29070 ( .DIN1(n32940), .DIN2(n34161), .Q(n36358) );
  hi1s1 U29071 ( .DIN1(n32984), .Q(n32940) );
  or2s1 U29072 ( .DIN1(n36359), .DIN2(n36360), .Q(n32984) );
  or2s1 U29073 ( .DIN1(n36136), .DIN2(n36361), .Q(n36360) );
  hi1s1 U29074 ( .DIN1(u5_state[13]), .Q(n36361) );
  or2s1 U29075 ( .DIN1(n36362), .DIN2(n36363), .Q(n36136) );
  or2s1 U29076 ( .DIN1(u5_state[12]), .DIN2(n36138), .Q(n36359) );
  or2s1 U29077 ( .DIN1(n34111), .DIN2(n36364), .Q(n36357) );
  or2s1 U29078 ( .DIN1(n34341), .DIN2(n32858), .Q(n36364) );
  and2s1 U29079 ( .DIN1(u5_state[39]), .DIN2(n36365), .Q(n32858) );
  hi1s1 U29080 ( .DIN1(n36366), .Q(n36365) );
  or2s1 U29081 ( .DIN1(u5_state[33]), .DIN2(n36160), .Q(n36366) );
  or2s1 U29082 ( .DIN1(n36367), .DIN2(n36368), .Q(n36160) );
  or2s1 U29083 ( .DIN1(n36107), .DIN2(n36369), .Q(n36368) );
  or2s1 U29084 ( .DIN1(u5_state[29]), .DIN2(n36370), .Q(n36367) );
  and2s1 U29085 ( .DIN1(n34350), .DIN2(n33871), .Q(n34341) );
  and2s1 U29086 ( .DIN1(u5_state[50]), .DIN2(n36371), .Q(n33871) );
  hi1s1 U29087 ( .DIN1(n36372), .Q(n36371) );
  or2s1 U29088 ( .DIN1(u5_state[4]), .DIN2(n36373), .Q(n36372) );
  hi1s1 U29089 ( .DIN1(u5_tmr2_done), .Q(n34350) );
  hi1s1 U29090 ( .DIN1(n15502), .Q(n35054) );
  or2s1 U29091 ( .DIN1(n36374), .DIN2(n36375), .Q(n9092) );
  and2s1 U29092 ( .DIN1(n36376), .DIN2(n36377), .Q(n36374) );
  or2s1 U29093 ( .DIN1(u5_state[53]), .DIN2(n36378), .Q(n36377) );
  or2s1 U29094 ( .DIN1(u5_state[54]), .DIN2(n36205), .Q(n36376) );
  hi1s1 U29095 ( .DIN1(u5_state[53]), .Q(n36205) );
  and2s1 U29096 ( .DIN1(n15474), .DIN2(n36379), .Q(n19413) );
  and2s1 U29097 ( .DIN1(n34143), .DIN2(n15508), .Q(n36379) );
  hi1s1 U29098 ( .DIN1(n34151), .Q(n34143) );
  or2s1 U29099 ( .DIN1(u5_ir_cnt[1]), .DIN2(u5_ir_cnt[0]), .Q(n34151) );
  and2s1 U29100 ( .DIN1(n36380), .DIN2(n35779), .Q(n19412) );
  hi1s1 U29101 ( .DIN1(n35618), .Q(n35779) );
  or2s1 U29102 ( .DIN1(n35762), .DIN2(n36381), .Q(n35618) );
  or2s1 U29103 ( .DIN1(u5_timer[6]), .DIN2(u5_timer[5]), .Q(n36381) );
  or2s1 U29104 ( .DIN1(n35743), .DIN2(n36382), .Q(n35762) );
  or2s1 U29105 ( .DIN1(u5_timer[4]), .DIN2(u5_timer[3]), .Q(n36382) );
  or2s1 U29106 ( .DIN1(u5_timer[0]), .DIN2(n36383), .Q(n35743) );
  or2s1 U29107 ( .DIN1(u5_timer[2]), .DIN2(u5_timer[1]), .Q(n36383) );
  hi1s1 U29108 ( .DIN1(u5_timer[7]), .Q(n36380) );
  hi1s1 U29109 ( .DIN1(n36176), .Q(n19410) );
  or2s1 U29110 ( .DIN1(n34348), .DIN2(n36384), .Q(n36176) );
  or2s1 U29111 ( .DIN1(n33896), .DIN2(n34117), .Q(n36384) );
  or2s1 U29112 ( .DIN1(n36385), .DIN2(n36386), .Q(n34117) );
  and2s1 U29113 ( .DIN1(n36387), .DIN2(n36388), .Q(n36386) );
  hi1s1 U29114 ( .DIN1(n36389), .Q(n36388) );
  and2s1 U29115 ( .DIN1(n36390), .DIN2(n36391), .Q(n36387) );
  or2s1 U29116 ( .DIN1(n36392), .DIN2(n36393), .Q(n36390) );
  and2s1 U29117 ( .DIN1(u5_state[59]), .DIN2(n36394), .Q(n36393) );
  hi1s1 U29118 ( .DIN1(n36395), .Q(n36394) );
  and2s1 U29119 ( .DIN1(n36396), .DIN2(n36397), .Q(n36392) );
  hi1s1 U29120 ( .DIN1(n36398), .Q(n36397) );
  or2s1 U29121 ( .DIN1(n36351), .DIN2(u5_state[59]), .Q(n36398) );
  and2s1 U29122 ( .DIN1(u5_state[55]), .DIN2(n36399), .Q(n36396) );
  and2s1 U29123 ( .DIN1(n36400), .DIN2(n36401), .Q(n36385) );
  and2s1 U29124 ( .DIN1(n36402), .DIN2(n36399), .Q(n36401) );
  hi1s1 U29125 ( .DIN1(n36403), .Q(n36399) );
  and2s1 U29126 ( .DIN1(n36404), .DIN2(n36405), .Q(n36402) );
  and2s1 U29127 ( .DIN1(u5_state[56]), .DIN2(n36349), .Q(n36400) );
  hi1s1 U29128 ( .DIN1(n36406), .Q(n33896) );
  or2s1 U29129 ( .DIN1(n36109), .DIN2(n36407), .Q(n36406) );
  or2s1 U29130 ( .DIN1(n36128), .DIN2(n36408), .Q(n36407) );
  hi1s1 U29131 ( .DIN1(u5_state[57]), .Q(n36408) );
  or2s1 U29132 ( .DIN1(n34121), .DIN2(n34111), .Q(n34348) );
  hi1s1 U29133 ( .DIN1(n36409), .Q(n34121) );
  or2s1 U29134 ( .DIN1(n36410), .DIN2(n36411), .Q(n36409) );
  or2s1 U29135 ( .DIN1(n36389), .DIN2(n36391), .Q(n36411) );
  hi1s1 U29136 ( .DIN1(u5_state[58]), .Q(n36391) );
  or2s1 U29137 ( .DIN1(u5_state[59]), .DIN2(n36395), .Q(n36410) );
  hi1s1 U29138 ( .DIN1(n36069), .Q(n19409) );
  or2s1 U29139 ( .DIN1(n36338), .DIN2(n36412), .Q(n36069) );
  or2s1 U29140 ( .DIN1(n34111), .DIN2(n34361), .Q(n36412) );
  or2s1 U29141 ( .DIN1(n34114), .DIN2(n34955), .Q(n34361) );
  or2s1 U29142 ( .DIN1(n36413), .DIN2(n34295), .Q(n34955) );
  hi1s1 U29143 ( .DIN1(n36414), .Q(n34295) );
  or2s1 U29144 ( .DIN1(n36415), .DIN2(n36416), .Q(n36414) );
  or2s1 U29145 ( .DIN1(n36417), .DIN2(n36404), .Q(n36416) );
  hi1s1 U29146 ( .DIN1(u5_state[44]), .Q(n36404) );
  or2s1 U29147 ( .DIN1(n36403), .DIN2(n36418), .Q(n36415) );
  and2s1 U29148 ( .DIN1(n34107), .DIN2(n34106), .Q(n36413) );
  and2s1 U29149 ( .DIN1(n36419), .DIN2(n36420), .Q(n34106) );
  hi1s1 U29150 ( .DIN1(n36421), .Q(n36420) );
  and2s1 U29151 ( .DIN1(n36422), .DIN2(n36111), .Q(n36419) );
  hi1s1 U29152 ( .DIN1(u5_state[41]), .Q(n36111) );
  and2s1 U29153 ( .DIN1(u5_state[42]), .DIN2(n36423), .Q(n34107) );
  and2s1 U29154 ( .DIN1(u5_state[53]), .DIN2(n36424), .Q(n34114) );
  and2s1 U29155 ( .DIN1(n36378), .DIN2(n36206), .Q(n36424) );
  hi1s1 U29156 ( .DIN1(n36375), .Q(n36206) );
  or2s1 U29157 ( .DIN1(n36425), .DIN2(n36426), .Q(n36375) );
  hi1s1 U29158 ( .DIN1(u5_state[54]), .Q(n36378) );
  hi1s1 U29159 ( .DIN1(n35041), .Q(n34111) );
  or2s1 U29160 ( .DIN1(n36427), .DIN2(n36428), .Q(n35041) );
  or2s1 U29161 ( .DIN1(n36417), .DIN2(n36405), .Q(n36428) );
  hi1s1 U29162 ( .DIN1(u5_state[52]), .Q(n36405) );
  or2s1 U29163 ( .DIN1(n36403), .DIN2(n36429), .Q(n36427) );
  or2s1 U29164 ( .DIN1(u5_state[56]), .DIN2(u5_state[44]), .Q(n36429) );
  or2s1 U29165 ( .DIN1(n36430), .DIN2(n36431), .Q(n36338) );
  or2s1 U29166 ( .DIN1(n33865), .DIN2(n36432), .Q(n36431) );
  or2s1 U29167 ( .DIN1(n32853), .DIN2(n34297), .Q(n36432) );
  hi1s1 U29168 ( .DIN1(n36433), .Q(n34297) );
  or2s1 U29169 ( .DIN1(n36434), .DIN2(n36435), .Q(n36433) );
  or2s1 U29170 ( .DIN1(n36122), .DIN2(n36436), .Q(n36435) );
  hi1s1 U29171 ( .DIN1(u5_state[37]), .Q(n36436) );
  or2s1 U29172 ( .DIN1(u5_state[3]), .DIN2(n36124), .Q(n36434) );
  hi1s1 U29173 ( .DIN1(n36437), .Q(n32853) );
  or2s1 U29174 ( .DIN1(n36438), .DIN2(n36439), .Q(n36437) );
  or2s1 U29175 ( .DIN1(n36143), .DIN2(n36440), .Q(n36439) );
  hi1s1 U29176 ( .DIN1(u5_state[38]), .Q(n36440) );
  or2s1 U29177 ( .DIN1(u5_state[36]), .DIN2(u5_state[0]), .Q(n36438) );
  or2s1 U29178 ( .DIN1(n36441), .DIN2(n36442), .Q(n33865) );
  or2s1 U29179 ( .DIN1(n32846), .DIN2(n34102), .Q(n36442) );
  and2s1 U29180 ( .DIN1(u5_state[41]), .DIN2(n36443), .Q(n34102) );
  and2s1 U29181 ( .DIN1(n36422), .DIN2(n36112), .Q(n36443) );
  and2s1 U29182 ( .DIN1(n36423), .DIN2(n36444), .Q(n36112) );
  hi1s1 U29183 ( .DIN1(n36445), .Q(n36444) );
  or2s1 U29184 ( .DIN1(u5_state[42]), .DIN2(n36421), .Q(n36445) );
  hi1s1 U29185 ( .DIN1(n36446), .Q(n36423) );
  hi1s1 U29186 ( .DIN1(u5_state[40]), .Q(n36422) );
  hi1s1 U29187 ( .DIN1(n36447), .Q(n32846) );
  or2s1 U29188 ( .DIN1(n36448), .DIN2(n36449), .Q(n36447) );
  or2s1 U29189 ( .DIN1(n36143), .DIN2(n36450), .Q(n36449) );
  hi1s1 U29190 ( .DIN1(u5_state[36]), .Q(n36450) );
  or2s1 U29191 ( .DIN1(n36122), .DIN2(n36451), .Q(n36143) );
  or2s1 U29192 ( .DIN1(n36452), .DIN2(n36446), .Q(n36122) );
  or2s1 U29193 ( .DIN1(n36453), .DIN2(n36454), .Q(n36446) );
  or2s1 U29194 ( .DIN1(n36455), .DIN2(n36395), .Q(n36453) );
  or2s1 U29195 ( .DIN1(u5_state[38]), .DIN2(u5_state[0]), .Q(n36448) );
  or2s1 U29196 ( .DIN1(n19411), .DIN2(n34247), .Q(n36441) );
  and2s1 U29197 ( .DIN1(u5_state[45]), .DIN2(n36456), .Q(n34247) );
  hi1s1 U29198 ( .DIN1(n36457), .Q(n36456) );
  or2s1 U29199 ( .DIN1(u5_state[43]), .DIN2(n36458), .Q(n36457) );
  and2s1 U29200 ( .DIN1(u5_state[43]), .DIN2(n36459), .Q(n19411) );
  hi1s1 U29201 ( .DIN1(n36460), .Q(n36459) );
  or2s1 U29202 ( .DIN1(u5_state[45]), .DIN2(n36458), .Q(n36460) );
  or2s1 U29203 ( .DIN1(n36461), .DIN2(n36426), .Q(n36458) );
  or2s1 U29204 ( .DIN1(n36370), .DIN2(n36108), .Q(n36426) );
  or2s1 U29205 ( .DIN1(n32856), .DIN2(n36462), .Q(n36430) );
  or2s1 U29206 ( .DIN1(n34368), .DIN2(n32878), .Q(n36462) );
  and2s1 U29207 ( .DIN1(u5_state[60]), .DIN2(n36463), .Q(n32878) );
  hi1s1 U29208 ( .DIN1(n36464), .Q(n36463) );
  or2s1 U29209 ( .DIN1(n36308), .DIN2(n36465), .Q(n36464) );
  hi1s1 U29210 ( .DIN1(n36466), .Q(n34368) );
  or2s1 U29211 ( .DIN1(n36467), .DIN2(n36468), .Q(n36466) );
  or2s1 U29212 ( .DIN1(n36469), .DIN2(n36470), .Q(n36468) );
  hi1s1 U29213 ( .DIN1(u5_state[61]), .Q(n36469) );
  or2s1 U29214 ( .DIN1(n36471), .DIN2(n36472), .Q(n36467) );
  or2s1 U29215 ( .DIN1(u5_state[8]), .DIN2(u5_state[1]), .Q(n36472) );
  and2s1 U29216 ( .DIN1(n36473), .DIN2(n36474), .Q(n32856) );
  and2s1 U29217 ( .DIN1(n36349), .DIN2(u5_state[46]), .Q(n36474) );
  hi1s1 U29218 ( .DIN1(n36417), .Q(n36349) );
  or2s1 U29219 ( .DIN1(n36389), .DIN2(n36475), .Q(n36417) );
  or2s1 U29220 ( .DIN1(u5_state[55]), .DIN2(n36455), .Q(n36475) );
  or2s1 U29221 ( .DIN1(n36476), .DIN2(n36454), .Q(n36389) );
  or2s1 U29222 ( .DIN1(n36477), .DIN2(n36478), .Q(n36454) );
  or2s1 U29223 ( .DIN1(n36452), .DIN2(n36421), .Q(n36476) );
  hi1s1 U29224 ( .DIN1(n36479), .Q(n36473) );
  or2s1 U29225 ( .DIN1(u5_state[47]), .DIN2(n36351), .Q(n36479) );
  and2s1 U29226 ( .DIN1(n36480), .DIN2(n15523), .Q(n19407) );
  and2s1 U29227 ( .DIN1(n15488), .DIN2(n15470), .Q(n36480) );
  hi1s1 U29228 ( .DIN1(n32217), .Q(n19406) );
  or2s1 U29229 ( .DIN1(n36481), .DIN2(n36482), .Q(n32217) );
  or2s1 U29230 ( .DIN1(n36483), .DIN2(n36484), .Q(n36482) );
  or2s1 U29231 ( .DIN1(n36485), .DIN2(n36486), .Q(n36484) );
  hi1s1 U29232 ( .DIN1(n36590), .Q(n36483) );
  or2s1 U29233 ( .DIN1(n36487), .DIN2(n36488), .Q(n36481) );
  or2s1 U29234 ( .DIN1(n32033), .DIN2(n36489), .Q(n36488) );
  hi1s1 U29235 ( .DIN1(n36490), .Q(n19405) );
  or2s1 U29236 ( .DIN1(n36491), .DIN2(n36492), .Q(n36490) );
  or2s1 U29237 ( .DIN1(n36486), .DIN2(n36493), .Q(n36492) );
  or2s1 U29238 ( .DIN1(n36487), .DIN2(n36485), .Q(n36493) );
  hi1s1 U29239 ( .DIN1(n36592), .Q(n36485) );
  hi1s1 U29240 ( .DIN1(n36593), .Q(n36487) );
  hi1s1 U29241 ( .DIN1(n36591), .Q(n36486) );
  or2s1 U29242 ( .DIN1(n36489), .DIN2(n36494), .Q(n36491) );
  or2s1 U29243 ( .DIN1(n36590), .DIN2(n32033), .Q(n36494) );
  hi1s1 U29244 ( .DIN1(n36609), .Q(n32033) );
  hi1s1 U29245 ( .DIN1(n36594), .Q(n36489) );
  and2s1 U29246 ( .DIN1(wb_cyc_i), .DIN2(n36495), .Q(n19404) );
  hi1s1 U29247 ( .DIN1(n36597), .Q(n36495) );
  and2s1 U29248 ( .DIN1(n36496), .DIN2(u1_u0_inc_in[11]), .Q(N884) );
  or2s1 U29249 ( .DIN1(n36497), .DIN2(n36498), .Q(N883) );
  hi1s1 U29250 ( .DIN1(n36499), .Q(n36498) );
  or2s1 U29251 ( .DIN1(n36500), .DIN2(u1_u0_inc_in[11]), .Q(n36499) );
  and2s1 U29252 ( .DIN1(u1_u0_inc_in[11]), .DIN2(n36500), .Q(n36497) );
  hi1s1 U29253 ( .DIN1(n36496), .Q(n36500) );
  and2s1 U29254 ( .DIN1(n36501), .DIN2(n36502), .Q(n36496) );
  and2s1 U29255 ( .DIN1(u1_u0_inc_in[9]), .DIN2(u1_u0_inc_in[10]), .Q(n36502) );
  or2s1 U29256 ( .DIN1(n36503), .DIN2(n36504), .Q(N882) );
  hi1s1 U29257 ( .DIN1(n36505), .Q(n36504) );
  or2s1 U29258 ( .DIN1(n36506), .DIN2(u1_u0_inc_in[10]), .Q(n36505) );
  and2s1 U29259 ( .DIN1(u1_u0_inc_in[10]), .DIN2(n36506), .Q(n36503) );
  or2s1 U29260 ( .DIN1(n36507), .DIN2(n36508), .Q(n36506) );
  or2s1 U29261 ( .DIN1(n36509), .DIN2(n36510), .Q(N881) );
  and2s1 U29262 ( .DIN1(n36501), .DIN2(n36507), .Q(n36510) );
  hi1s1 U29263 ( .DIN1(u1_u0_inc_in[9]), .Q(n36507) );
  and2s1 U29264 ( .DIN1(u1_u0_inc_in[9]), .DIN2(n36508), .Q(n36509) );
  hi1s1 U29265 ( .DIN1(n36501), .Q(n36508) );
  and2s1 U29266 ( .DIN1(u1_u0_inc_in[8]), .DIN2(n36511), .Q(n36501) );
  or2s1 U29267 ( .DIN1(n36512), .DIN2(n36513), .Q(N880) );
  hi1s1 U29268 ( .DIN1(n36514), .Q(n36513) );
  or2s1 U29269 ( .DIN1(n36515), .DIN2(u1_u0_inc_in[8]), .Q(n36514) );
  and2s1 U29270 ( .DIN1(u1_u0_inc_in[8]), .DIN2(n36515), .Q(n36512) );
  hi1s1 U29271 ( .DIN1(n36511), .Q(n36515) );
  and2s1 U29272 ( .DIN1(u1_u0_inc_in[7]), .DIN2(n36516), .Q(n36511) );
  or2s1 U29273 ( .DIN1(n36517), .DIN2(n36518), .Q(N879) );
  hi1s1 U29274 ( .DIN1(n36519), .Q(n36518) );
  or2s1 U29275 ( .DIN1(n36520), .DIN2(u1_u0_inc_in[7]), .Q(n36519) );
  and2s1 U29276 ( .DIN1(u1_u0_inc_in[7]), .DIN2(n36520), .Q(n36517) );
  hi1s1 U29277 ( .DIN1(n36516), .Q(n36520) );
  and2s1 U29278 ( .DIN1(u1_u0_inc_in[6]), .DIN2(n36521), .Q(n36516) );
  or2s1 U29279 ( .DIN1(n36522), .DIN2(n36523), .Q(N878) );
  and2s1 U29280 ( .DIN1(n36521), .DIN2(n36524), .Q(n36523) );
  hi1s1 U29281 ( .DIN1(u1_u0_inc_in[6]), .Q(n36524) );
  hi1s1 U29282 ( .DIN1(n36525), .Q(n36521) );
  and2s1 U29283 ( .DIN1(u1_u0_inc_in[6]), .DIN2(n36525), .Q(n36522) );
  or2s1 U29284 ( .DIN1(n36526), .DIN2(n36527), .Q(n36525) );
  or2s1 U29285 ( .DIN1(n36528), .DIN2(n36529), .Q(N877) );
  and2s1 U29286 ( .DIN1(n36530), .DIN2(n36526), .Q(n36529) );
  hi1s1 U29287 ( .DIN1(u1_u0_inc_in[5]), .Q(n36526) );
  hi1s1 U29288 ( .DIN1(n36527), .Q(n36530) );
  and2s1 U29289 ( .DIN1(u1_u0_inc_in[5]), .DIN2(n36527), .Q(n36528) );
  or2s1 U29290 ( .DIN1(n36531), .DIN2(n36532), .Q(n36527) );
  or2s1 U29291 ( .DIN1(n36533), .DIN2(n36534), .Q(N876) );
  and2s1 U29292 ( .DIN1(n36535), .DIN2(n36531), .Q(n36534) );
  hi1s1 U29293 ( .DIN1(u1_u0_inc_in[4]), .Q(n36531) );
  hi1s1 U29294 ( .DIN1(n36532), .Q(n36535) );
  and2s1 U29295 ( .DIN1(u1_u0_inc_in[4]), .DIN2(n36532), .Q(n36533) );
  or2s1 U29296 ( .DIN1(n36536), .DIN2(n36537), .Q(n36532) );
  or2s1 U29297 ( .DIN1(n36538), .DIN2(n36539), .Q(N875) );
  and2s1 U29298 ( .DIN1(n36540), .DIN2(n36536), .Q(n36539) );
  hi1s1 U29299 ( .DIN1(u1_u0_inc_in[3]), .Q(n36536) );
  hi1s1 U29300 ( .DIN1(n36537), .Q(n36540) );
  and2s1 U29301 ( .DIN1(u1_u0_inc_in[3]), .DIN2(n36537), .Q(n36538) );
  or2s1 U29302 ( .DIN1(n36541), .DIN2(n36542), .Q(n36537) );
  or2s1 U29303 ( .DIN1(n36543), .DIN2(n36544), .Q(N874) );
  and2s1 U29304 ( .DIN1(n36545), .DIN2(n36541), .Q(n36544) );
  hi1s1 U29305 ( .DIN1(u1_u0_inc_in[2]), .Q(n36541) );
  hi1s1 U29306 ( .DIN1(n36542), .Q(n36545) );
  and2s1 U29307 ( .DIN1(u1_u0_inc_in[2]), .DIN2(n36542), .Q(n36543) );
  or2s1 U29308 ( .DIN1(N872), .DIN2(n36546), .Q(n36542) );
  or2s1 U29309 ( .DIN1(n36547), .DIN2(n36548), .Q(N873) );
  and2s1 U29310 ( .DIN1(u1_u0_inc_in[0]), .DIN2(n36546), .Q(n36548) );
  hi1s1 U29311 ( .DIN1(u1_u0_inc_in[1]), .Q(n36546) );
  and2s1 U29312 ( .DIN1(u1_u0_inc_in[1]), .DIN2(N872), .Q(n36547) );
  hi1s1 U29313 ( .DIN1(u1_u0_inc_in[0]), .Q(N872) );
  hi1s1 U29314 ( .DIN1(n32812), .Q(N1549) );
  or2s1 U29315 ( .DIN1(n36549), .DIN2(n36550), .Q(n32812) );
  or2s1 U29316 ( .DIN1(n36551), .DIN2(n36552), .Q(n36550) );
  or2s1 U29317 ( .DIN1(n36553), .DIN2(n36554), .Q(n36552) );
  or2s1 U29318 ( .DIN1(n36555), .DIN2(n36556), .Q(n36554) );
  and2s1 U29319 ( .DIN1(u0_csr_r2[1]), .DIN2(n32770), .Q(n36556) );
  hi1s1 U29320 ( .DIN1(u4_ps_cnt[1]), .Q(n32770) );
  and2s1 U29321 ( .DIN1(u4_ps_cnt[1]), .DIN2(n32826), .Q(n36555) );
  hi1s1 U29322 ( .DIN1(u0_csr_r2[1]), .Q(n32826) );
  or2s1 U29323 ( .DIN1(n36557), .DIN2(n36558), .Q(n36553) );
  and2s1 U29324 ( .DIN1(u0_csr_r2[0]), .DIN2(n32775), .Q(n36558) );
  hi1s1 U29325 ( .DIN1(u4_ps_cnt[0]), .Q(n32775) );
  and2s1 U29326 ( .DIN1(u4_ps_cnt[0]), .DIN2(n32825), .Q(n36557) );
  hi1s1 U29327 ( .DIN1(u0_csr_r2[0]), .Q(n32825) );
  or2s1 U29328 ( .DIN1(n36559), .DIN2(n36560), .Q(n36551) );
  or2s1 U29329 ( .DIN1(n36561), .DIN2(n36562), .Q(n36560) );
  and2s1 U29330 ( .DIN1(u0_csr_r2[5]), .DIN2(n32799), .Q(n36562) );
  hi1s1 U29331 ( .DIN1(u4_ps_cnt[5]), .Q(n32799) );
  and2s1 U29332 ( .DIN1(u4_ps_cnt[5]), .DIN2(n32820), .Q(n36561) );
  hi1s1 U29333 ( .DIN1(u0_csr_r2[5]), .Q(n32820) );
  or2s1 U29334 ( .DIN1(n36563), .DIN2(n36564), .Q(n36559) );
  and2s1 U29335 ( .DIN1(u0_csr_r2[3]), .DIN2(n32784), .Q(n36564) );
  hi1s1 U29336 ( .DIN1(u4_ps_cnt[3]), .Q(n32784) );
  and2s1 U29337 ( .DIN1(u4_ps_cnt[3]), .DIN2(n32824), .Q(n36563) );
  hi1s1 U29338 ( .DIN1(u0_csr_r2[3]), .Q(n32824) );
  or2s1 U29339 ( .DIN1(n36565), .DIN2(n36566), .Q(n36549) );
  or2s1 U29340 ( .DIN1(n36567), .DIN2(n36568), .Q(n36566) );
  or2s1 U29341 ( .DIN1(n36569), .DIN2(n36570), .Q(n36568) );
  and2s1 U29342 ( .DIN1(u0_csr_r2[7]), .DIN2(n32762), .Q(n36570) );
  hi1s1 U29343 ( .DIN1(u4_ps_cnt[7]), .Q(n32762) );
  and2s1 U29344 ( .DIN1(u4_ps_cnt[7]), .DIN2(n32818), .Q(n36569) );
  hi1s1 U29345 ( .DIN1(u0_csr_r2[7]), .Q(n32818) );
  or2s1 U29346 ( .DIN1(n36571), .DIN2(n36572), .Q(n36567) );
  and2s1 U29347 ( .DIN1(u0_csr_r2[2]), .DIN2(n32778), .Q(n36572) );
  hi1s1 U29348 ( .DIN1(u4_ps_cnt[2]), .Q(n32778) );
  and2s1 U29349 ( .DIN1(u4_ps_cnt[2]), .DIN2(n32823), .Q(n36571) );
  hi1s1 U29350 ( .DIN1(u0_csr_r2[2]), .Q(n32823) );
  or2s1 U29351 ( .DIN1(n36573), .DIN2(n36574), .Q(n36565) );
  or2s1 U29352 ( .DIN1(n36575), .DIN2(n36576), .Q(n36574) );
  and2s1 U29353 ( .DIN1(u0_csr_r2[4]), .DIN2(n32793), .Q(n36576) );
  hi1s1 U29354 ( .DIN1(u4_ps_cnt[4]), .Q(n32793) );
  and2s1 U29355 ( .DIN1(u4_ps_cnt[4]), .DIN2(n32819), .Q(n36575) );
  hi1s1 U29356 ( .DIN1(u0_csr_r2[4]), .Q(n32819) );
  or2s1 U29357 ( .DIN1(n36577), .DIN2(n36578), .Q(n36573) );
  and2s1 U29358 ( .DIN1(u0_csr_r2[6]), .DIN2(n32759), .Q(n36578) );
  hi1s1 U29359 ( .DIN1(u4_ps_cnt[6]), .Q(n32759) );
  and2s1 U29360 ( .DIN1(u4_ps_cnt[6]), .DIN2(n32817), .Q(n36577) );
  hi1s1 U29361 ( .DIN1(u0_csr_r2[6]), .Q(n32817) );
endmodule

