module c1908 ( N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, N37, 
    N40, N43, N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79, N82, N85, 
    N88, N91, N94, N99, N104, N2753, N2754, N2755, N2756, N2762, N2767, N2768, 
    N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786, N2787, N2811, 
    N2886, N2887, N2888, N2889, N2890, N2891, N2892, N2899 );
input  N1, N4, N7, N10, N13, N16, N19, N22, N25, N28, N31, N34, N37, N40, N43, 
    N46, N49, N53, N56, N60, N63, N66, N69, N72, N76, N79, N82, N85, N88, N91, 
    N94, N99, N104;
output N2753, N2754, N2755, N2756, N2762, N2767, N2768, N2779, N2780, N2781, 
    N2782, N2783, N2784, N2785, N2786, N2787, N2811, N2886, N2887, N2888, 
    N2889, N2890, N2891, N2892, N2899;
    wire n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
        n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
        n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
        n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
        n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
        n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
        n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
        n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
        n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
        n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
        n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
        n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
        n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
        n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
        n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
        n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
        n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
        n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
        n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
        n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
        n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
        n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
        n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
        n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
        n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
        n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
        n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
        n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
        n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
        n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
        n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
        n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
        n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
        n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
        n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
        n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
        n811, n812, n813, n814, n815, n816, n817, n818, n819, n820;
    nor2s1 U1 ( .Q(N2899), .DIN1(n380), .DIN2(n381) );
    nor2s1 U2 ( .Q(N2887), .DIN1(n380), .DIN2(n382) );
    nor2s1 U3 ( .Q(N2886), .DIN1(n380), .DIN2(n383) );
    nnd2s1 U4 ( .Q(N2811), .DIN1(n384), .DIN2(n385) );
    nor2s1 U5 ( .Q(N2890), .DIN1(n380), .DIN2(n386) );
    nor2s1 U6 ( .Q(N2889), .DIN1(n380), .DIN2(n387) );
    nor2s1 U7 ( .Q(N2888), .DIN1(n380), .DIN2(n388) );
    nor2s1 U8 ( .Q(n389), .DIN1(n390), .DIN2(n391) );
    nor2s1 U9 ( .Q(n392), .DIN1(n393), .DIN2(n394) );
    nor2s1 U10 ( .Q(n395), .DIN1(n396), .DIN2(n397) );
    hi1s1 U11 ( .Q(n398), .DIN(N104) );
    hi1s1 U12 ( .Q(n399), .DIN(N72) );
    hi1s1 U13 ( .Q(n400), .DIN(N69) );
    hi1s1 U14 ( .Q(n401), .DIN(N94) );
    nor2s1 U15 ( .Q(n391), .DIN1(n390), .DIN2(n402) );
    nor2s1 U16 ( .Q(n403), .DIN1(n404), .DIN2(n405) );
    nnd2s1 U17 ( .Q(n406), .DIN1(n391), .DIN2(n407) );
    nnd2s1 U18 ( .Q(n408), .DIN1(n409), .DIN2(n410) );
    nor2s1 U19 ( .Q(n411), .DIN1(n406), .DIN2(n412) );
    nnd2s1 U20 ( .Q(n413), .DIN1(n414), .DIN2(n415) );
    nor2s1 U21 ( .Q(n416), .DIN1(n410), .DIN2(n409) );
    nnd2s1 U22 ( .Q(n417), .DIN1(n414), .DIN2(n418) );
    nor2s1 U23 ( .Q(n419), .DIN1(n420), .DIN2(n410) );
    nnd2s1 U24 ( .Q(n421), .DIN1(n415), .DIN2(n422) );
    nnd2s1 U25 ( .Q(n423), .DIN1(n404), .DIN2(n424) );
    nnd2s1 U26 ( .Q(n425), .DIN1(n410), .DIN2(n420) );
    nor2s1 U27 ( .Q(n426), .DIN1(n423), .DIN2(n406) );
    nor2s1 U28 ( .Q(n427), .DIN1(n398), .DIN2(N91) );
    nnd2s1 U29 ( .Q(n428), .DIN1(n390), .DIN2(n429) );
    nor2s1 U30 ( .Q(n430), .DIN1(n431), .DIN2(n428) );
    nor2s1 U31 ( .Q(n432), .DIN1(n433), .DIN2(n423) );
    nnd2s1 U32 ( .Q(n434), .DIN1(n435), .DIN2(n436) );
    nnd2s1 U33 ( .Q(n437), .DIN1(n438), .DIN2(n439) );
    nor2s1 U34 ( .Q(n440), .DIN1(n401), .DIN2(n441) );
    nnd2s1 U35 ( .Q(n393), .DIN1(n442), .DIN2(N99) );
    nor2s1 U36 ( .Q(n441), .DIN1(n437), .DIN2(n434) );
    nor2s1 U37 ( .Q(n443), .DIN1(n444), .DIN2(n445) );
    nnd2s1 U38 ( .Q(n446), .DIN1(n447), .DIN2(n448) );
    nor2s1 U39 ( .Q(n449), .DIN1(n450), .DIN2(n451) );
    nor2s1 U40 ( .Q(n452), .DIN1(n453), .DIN2(n454) );
    nor2s1 U41 ( .Q(n455), .DIN1(n456), .DIN2(n457) );
    nnd2s1 U42 ( .Q(n458), .DIN1(n459), .DIN2(n460) );
    nor2s1 U43 ( .Q(n461), .DIN1(n462), .DIN2(n463) );
    nnd2s1 U44 ( .Q(n464), .DIN1(n465), .DIN2(n466) );
    nnd2s1 U45 ( .Q(n467), .DIN1(n468), .DIN2(n469) );
    nnd2s1 U46 ( .Q(n422), .DIN1(n470), .DIN2(n471) );
    nnd2s1 U47 ( .Q(n472), .DIN1(n473), .DIN2(n474) );
    nor2s1 U48 ( .Q(n415), .DIN1(n475), .DIN2(n476) );
    nnd2s1 U49 ( .Q(n477), .DIN1(n478), .DIN2(n479) );
    nnd2s1 U50 ( .Q(n420), .DIN1(n480), .DIN2(n481) );
    nor2s1 U51 ( .Q(n410), .DIN1(n482), .DIN2(n483) );
    nor2s1 U52 ( .Q(n484), .DIN1(n485), .DIN2(n486) );
    nor2s1 U53 ( .Q(n487), .DIN1(n488), .DIN2(n489) );
    nnd2s1 U54 ( .Q(n404), .DIN1(n490), .DIN2(n491) );
    nnd2s1 U55 ( .Q(n492), .DIN1(n493), .DIN2(n494) );
    nor2s1 U56 ( .Q(n495), .DIN1(n496), .DIN2(n497) );
    nor2s1 U57 ( .Q(n390), .DIN1(n498), .DIN2(n499) );
    nnd2s1 U58 ( .Q(N2892), .DIN1(n500), .DIN2(n501) );
    nnd2s1 U59 ( .Q(N2891), .DIN1(n502), .DIN2(n503) );
    nnd2s1 U60 ( .Q(N2787), .DIN1(n504), .DIN2(n505) );
    nnd2s1 U61 ( .Q(N2786), .DIN1(n506), .DIN2(n507) );
    nnd2s1 U62 ( .Q(N2785), .DIN1(n508), .DIN2(n509) );
    nnd2s1 U63 ( .Q(N2784), .DIN1(n510), .DIN2(n511) );
    nnd2s1 U64 ( .Q(N2783), .DIN1(n512), .DIN2(n513) );
    nnd2s1 U65 ( .Q(N2782), .DIN1(n514), .DIN2(n515) );
    nnd2s1 U66 ( .Q(N2781), .DIN1(n516), .DIN2(n517) );
    nnd2s1 U67 ( .Q(N2780), .DIN1(n518), .DIN2(n519) );
    nnd2s1 U68 ( .Q(N2779), .DIN1(n520), .DIN2(n521) );
    nnd2s1 U69 ( .Q(N2768), .DIN1(n522), .DIN2(n523) );
    nnd2s1 U70 ( .Q(N2767), .DIN1(n524), .DIN2(n525) );
    nnd2s1 U71 ( .Q(N2762), .DIN1(n526), .DIN2(n527) );
    nnd2s1 U72 ( .Q(N2756), .DIN1(n528), .DIN2(n529) );
    nnd2s1 U73 ( .Q(N2755), .DIN1(n530), .DIN2(n531) );
    nnd2s1 U74 ( .Q(N2754), .DIN1(n532), .DIN2(n533) );
    nnd2s1 U75 ( .Q(N2753), .DIN1(n534), .DIN2(n535) );
    nnd2s1 U76 ( .Q(n382), .DIN1(n536), .DIN2(n537) );
    nnd2s1 U77 ( .Q(n383), .DIN1(n538), .DIN2(n539) );
    nor2s1 U78 ( .Q(n540), .DIN1(N104), .DIN2(N72) );
    nor2s1 U79 ( .Q(n541), .DIN1(n542), .DIN2(n543) );
    nnd2s1 U80 ( .Q(n544), .DIN1(n545), .DIN2(n546) );
    nor2s1 U81 ( .Q(n547), .DIN1(n548), .DIN2(n549) );
    nor2s1 U82 ( .Q(n550), .DIN1(n551), .DIN2(n552) );
    nnd2s1 U83 ( .Q(n553), .DIN1(n554), .DIN2(n555) );
    nor2s1 U84 ( .Q(n556), .DIN1(N104), .DIN2(n400) );
    nnd2s1 U85 ( .Q(n557), .DIN1(n558), .DIN2(n559) );
    nnd2s1 U86 ( .Q(n560), .DIN1(n561), .DIN2(n562) );
    nor2s1 U87 ( .Q(n563), .DIN1(n564), .DIN2(n565) );
    nor2s1 U88 ( .Q(n566), .DIN1(n567), .DIN2(n568) );
    nnd2s1 U89 ( .Q(n569), .DIN1(n570), .DIN2(n571) );
    nnd2s1 U90 ( .Q(n572), .DIN1(n573), .DIN2(n574) );
    nor2s1 U91 ( .Q(n575), .DIN1(n576), .DIN2(n577) );
    nor2s1 U92 ( .Q(n578), .DIN1(n579), .DIN2(n580) );
    nnd2s1 U93 ( .Q(n581), .DIN1(n582), .DIN2(n583) );
    nor2s1 U94 ( .Q(n584), .DIN1(n585), .DIN2(n586) );
    nnd2s1 U95 ( .Q(n587), .DIN1(n588), .DIN2(n589) );
    nor2s1 U96 ( .Q(n590), .DIN1(n591), .DIN2(n401) );
    nor2s1 U97 ( .Q(n442), .DIN1(N104), .DIN2(n591) );
    nnd2s1 U98 ( .Q(n592), .DIN1(n593), .DIN2(n594) );
    nnd2s1 U99 ( .Q(n595), .DIN1(n596), .DIN2(n597) );
    nor2s1 U100 ( .Q(n598), .DIN1(n599), .DIN2(n600) );
    nnd2s1 U101 ( .Q(n601), .DIN1(n602), .DIN2(n603) );
    nnd2s1 U102 ( .Q(n604), .DIN1(n605), .DIN2(n606) );
    nnd2s1 U103 ( .Q(n607), .DIN1(n608), .DIN2(n609) );
    nnd2s1 U104 ( .Q(n610), .DIN1(n611), .DIN2(n612) );
    nor2s1 U105 ( .Q(n613), .DIN1(n614), .DIN2(n615) );
    nnd2s1 U106 ( .Q(n431), .DIN1(n616), .DIN2(n617) );
    nor2s1 U107 ( .Q(n618), .DIN1(n421), .DIN2(n425) );
    nor2s1 U108 ( .Q(n619), .DIN1(n413), .DIN2(n620) );
    nor2s1 U109 ( .Q(n621), .DIN1(n417), .DIN2(n622) );
    nor2s1 U110 ( .Q(n623), .DIN1(n622), .DIN2(n421) );
    nnd2s1 U111 ( .Q(n433), .DIN1(n391), .DIN2(n616) );
    nor2s1 U112 ( .Q(n624), .DIN1(n412), .DIN2(n433) );
    nor2s1 U113 ( .Q(n625), .DIN1(n620), .DIN2(n421) );
    nnd2s1 U114 ( .Q(n626), .DIN1(n422), .DIN2(n418) );
    nnd2s1 U115 ( .Q(n627), .DIN1(n419), .DIN2(n432) );
    nor2s1 U116 ( .Q(n628), .DIN1(n620), .DIN2(n417) );
    nnd2s1 U117 ( .Q(n629), .DIN1(n630), .DIN2(n631) );
    nnd2s1 U118 ( .Q(n632), .DIN1(n633), .DIN2(n634) );
    nor2s1 U119 ( .Q(n436), .DIN1(n629), .DIN2(n632) );
    nnd2s1 U120 ( .Q(n635), .DIN1(n636), .DIN2(n637) );
    nnd2s1 U121 ( .Q(n638), .DIN1(n639), .DIN2(n640) );
    nor2s1 U122 ( .Q(n435), .DIN1(n635), .DIN2(n638) );
    nor2s1 U123 ( .Q(n641), .DIN1(N88), .DIN2(n591) );
    nor2s1 U124 ( .Q(n642), .DIN1(n398), .DIN2(n401) );
    nor2s1 U125 ( .Q(n643), .DIN1(n414), .DIN2(n415) );
    nor2s1 U126 ( .Q(n644), .DIN1(n408), .DIN2(n645) );
    nor2s1 U127 ( .Q(n646), .DIN1(n645), .DIN2(n413) );
    nor2s1 U128 ( .Q(n647), .DIN1(n645), .DIN2(n417) );
    nnd2s1 U129 ( .Q(n648), .DIN1(n411), .DIN2(n419) );
    nor2s1 U130 ( .Q(n649), .DIN1(n413), .DIN2(n425) );
    nor2s1 U131 ( .Q(n650), .DIN1(n408), .DIN2(n417) );
    nor2s1 U132 ( .Q(n651), .DIN1(n408), .DIN2(n421) );
    nor2s1 U133 ( .Q(n652), .DIN1(n413), .DIN2(n622) );
    nnd2s1 U134 ( .Q(n653), .DIN1(n654), .DIN2(n655) );
    nnd2s1 U135 ( .Q(n656), .DIN1(n657), .DIN2(n658) );
    nor2s1 U136 ( .Q(n439), .DIN1(n653), .DIN2(n656) );
    nnd2s1 U137 ( .Q(n659), .DIN1(n660), .DIN2(n661) );
    nnd2s1 U138 ( .Q(n662), .DIN1(n663), .DIN2(n664) );
    nor2s1 U139 ( .Q(n438), .DIN1(n659), .DIN2(n662) );
    nor2s1 U140 ( .Q(n665), .DIN1(n666), .DIN2(n667) );
    nnd2s1 U141 ( .Q(n668), .DIN1(n669), .DIN2(n670) );
    nnd2s1 U142 ( .Q(n671), .DIN1(n672), .DIN2(n673) );
    nor2s1 U143 ( .Q(n674), .DIN1(n389), .DIN2(n408) );
    nnd2s1 U144 ( .Q(n394), .DIN1(n403), .DIN2(n675) );
    nnd2s1 U145 ( .Q(n396), .DIN1(n676), .DIN2(n677) );
    nnd2s1 U146 ( .Q(n397), .DIN1(n678), .DIN2(n679) );
    nor2s1 U147 ( .Q(n385), .DIN1(N104), .DIN2(n392) );
    nor2s1 U148 ( .Q(n384), .DIN1(n395), .DIN2(n680) );
    hi1s1 U149 ( .Q(n681), .DIN(N37) );
    hi1s1 U150 ( .Q(n682), .DIN(N34) );
    hi1s1 U151 ( .Q(n683), .DIN(N43) );
    hi1s1 U152 ( .Q(n684), .DIN(N28) );
    hi1s1 U153 ( .Q(n685), .DIN(N46) );
    hi1s1 U154 ( .Q(n686), .DIN(N19) );
    hi1s1 U155 ( .Q(n687), .DIN(N16) );
    hi1s1 U156 ( .Q(n688), .DIN(N13) );
    nnd2s1 U157 ( .Q(n689), .DIN1(N63), .DIN2(n398) );
    hi1s1 U158 ( .Q(n690), .DIN(N22) );
    hi1s1 U159 ( .Q(n691), .DIN(N10) );
    hi1s1 U160 ( .Q(n692), .DIN(N7) );
    hi1s1 U161 ( .Q(n693), .DIN(N4) );
    hi1s1 U162 ( .Q(n694), .DIN(N1) );
    nor2s1 U163 ( .Q(n695), .DIN1(n495), .DIN2(N94) );
    nnd2s1 U164 ( .Q(n696), .DIN1(N49), .DIN2(n697) );
    hi1s1 U165 ( .Q(n698), .DIN(N40) );
    nnd2s1 U166 ( .Q(n699), .DIN1(N66), .DIN2(n398) );
    nnd2s1 U167 ( .Q(n700), .DIN1(n701), .DIN2(n401) );
    nnd2s1 U168 ( .Q(n702), .DIN1(n540), .DIN2(N53) );
    nnd2s1 U169 ( .Q(n703), .DIN1(n467), .DIN2(n401) );
    nnd2s1 U170 ( .Q(n704), .DIN1(n556), .DIN2(N56) );
    nnd2s1 U171 ( .Q(n705), .DIN1(n472), .DIN2(n401) );
    nnd2s1 U172 ( .Q(n706), .DIN1(n556), .DIN2(N60) );
    nnd2s1 U173 ( .Q(n707), .DIN1(N56), .DIN2(n708) );
    nnd2s1 U174 ( .Q(n709), .DIN1(n477), .DIN2(n401) );
    nnd2s1 U175 ( .Q(n710), .DIN1(n540), .DIN2(N49) );
    nnd2s1 U176 ( .Q(n711), .DIN1(n712), .DIN2(n401) );
    nnd2s1 U177 ( .Q(n713), .DIN1(n440), .DIN2(N79) );
    nnd2s1 U178 ( .Q(n714), .DIN1(n665), .DIN2(n458) );
    nor2s1 U179 ( .Q(n715), .DIN1(n458), .DIN2(n665) );
    nor2s1 U180 ( .Q(n381), .DIN1(n716), .DIN2(n715) );
    nor2s1 U181 ( .Q(n717), .DIN1(n718), .DIN2(n452) );
    nor2s1 U182 ( .Q(n719), .DIN1(n720), .DIN2(n461) );
    nor2s1 U183 ( .Q(n721), .DIN1(n717), .DIN2(n427) );
    nnd2s1 U184 ( .Q(n722), .DIN1(n434), .DIN2(n398) );
    nor2s1 U185 ( .Q(n723), .DIN1(n724), .DIN2(n719) );
    nnd2s1 U186 ( .Q(n725), .DIN1(N104), .DIN2(n726) );
    nnd2s1 U187 ( .Q(n727), .DIN1(n437), .DIN2(n398) );
    nor2s1 U188 ( .Q(n728), .DIN1(n492), .DIN2(n729) );
    nnd2s1 U189 ( .Q(n730), .DIN1(N104), .DIN2(n731) );
    nnd2s1 U190 ( .Q(n732), .DIN1(n440), .DIN2(N56) );
    nor2s1 U191 ( .Q(n733), .DIN1(n477), .DIN2(n732) );
    nnd2s1 U192 ( .Q(n734), .DIN1(n732), .DIN2(n477) );
    nor2s1 U193 ( .Q(n386), .DIN1(n733), .DIN2(n735) );
    nnd2s1 U194 ( .Q(n736), .DIN1(n440), .DIN2(N85) );
    nor2s1 U195 ( .Q(n737), .DIN1(n472), .DIN2(n736) );
    nnd2s1 U196 ( .Q(n738), .DIN1(n736), .DIN2(n472) );
    nor2s1 U197 ( .Q(n387), .DIN1(n737), .DIN2(n739) );
    nnd2s1 U198 ( .Q(n740), .DIN1(n440), .DIN2(N82) );
    nor2s1 U199 ( .Q(n741), .DIN1(n467), .DIN2(n740) );
    nnd2s1 U200 ( .Q(n742), .DIN1(n740), .DIN2(n467) );
    nor2s1 U201 ( .Q(n388), .DIN1(n741), .DIN2(n743) );
    nnd2s1 U202 ( .Q(n631), .DIN1(n618), .DIN2(n430) );
    nnd2s1 U203 ( .Q(n630), .DIN1(n619), .DIN2(n430) );
    nnd2s1 U204 ( .Q(n634), .DIN1(n621), .DIN2(n430) );
    nnd2s1 U205 ( .Q(n633), .DIN1(n623), .DIN2(n430) );
    nnd2s1 U206 ( .Q(n637), .DIN1(n618), .DIN2(n624) );
    nnd2s1 U207 ( .Q(n655), .DIN1(n644), .DIN2(n643) );
    nnd2s1 U208 ( .Q(n654), .DIN1(n646), .DIN2(n416) );
    nnd2s1 U209 ( .Q(n658), .DIN1(n647), .DIN2(n419) );
    nor2s1 U210 ( .Q(n744), .DIN1(n648), .DIN2(n421) );
    nnd2s1 U211 ( .Q(n636), .DIN1(n625), .DIN2(n432) );
    nor2s1 U212 ( .Q(n745), .DIN1(n627), .DIN2(n626) );
    nnd2s1 U213 ( .Q(n639), .DIN1(n628), .DIN2(n432) );
    nnd2s1 U214 ( .Q(n661), .DIN1(n649), .DIN2(n426) );
    nnd2s1 U215 ( .Q(n660), .DIN1(n650), .DIN2(n426) );
    nnd2s1 U216 ( .Q(n664), .DIN1(n651), .DIN2(n426) );
    nnd2s1 U217 ( .Q(n663), .DIN1(n652), .DIN2(n426) );
    hi1s1 U218 ( .Q(n746), .DIN(n393) );
    hi1s1 U219 ( .Q(n657), .DIN(n744) );
    hi1s1 U220 ( .Q(n640), .DIN(n745) );
    nor2s1 U221 ( .Q(n380), .DIN1(n398), .DIN2(N99) );
    hi1s1 U222 ( .Q(n676), .DIN(n408) );
    nnd2s1 U223 ( .Q(n708), .DIN1(N69), .DIN2(n401) );
    nnd2s1 U224 ( .Q(n424), .DIN1(N60), .DIN2(n708) );
    hi1s1 U225 ( .Q(n412), .DIN(n403) );
    nnd2s1 U226 ( .Q(n697), .DIN1(n399), .DIN2(n401) );
    nnd2s1 U227 ( .Q(n429), .DIN1(N53), .DIN2(n697) );
    nor2s1 U228 ( .Q(n591), .DIN1(n400), .DIN2(n399) );
    nnd2s1 U229 ( .Q(n747), .DIN1(n642), .DIN2(n641) );
    nnd2s1 U230 ( .Q(n407), .DIN1(n393), .DIN2(n747) );
    hi1s1 U231 ( .Q(n620), .DIN(n416) );
    hi1s1 U232 ( .Q(n679), .DIN(n413) );
    hi1s1 U233 ( .Q(n622), .DIN(n419) );
    nnd2s1 U234 ( .Q(n748), .DIN1(n590), .DIN2(n427) );
    nnd2s1 U235 ( .Q(n616), .DIN1(n393), .DIN2(n748) );
    nnd2s1 U236 ( .Q(n726), .DIN1(N91), .DIN2(N66) );
    nor2s1 U237 ( .Q(n729), .DIN1(n398), .DIN2(N88) );
    nnd2s1 U238 ( .Q(n731), .DIN1(N88), .DIN2(N63) );
    nnd2s1 U239 ( .Q(n749), .DIN1(n423), .DIN2(n404) );
    nnd2s1 U240 ( .Q(n750), .DIN1(n746), .DIN2(n749) );
    nnd2s1 U241 ( .Q(n677), .DIN1(n412), .DIN2(n750) );
    nnd2s1 U242 ( .Q(n751), .DIN1(n421), .DIN2(n417) );
    nnd2s1 U243 ( .Q(n752), .DIN1(n622), .DIN2(n425) );
    nnd2s1 U244 ( .Q(n753), .DIN1(n679), .DIN2(n752) );
    nnd2s1 U245 ( .Q(n754), .DIN1(n676), .DIN2(n751) );
    nnd2s1 U246 ( .Q(n755), .DIN1(n754), .DIN2(n753) );
    nnd2s1 U247 ( .Q(n756), .DIN1(n674), .DIN2(n679) );
    nnd2s1 U248 ( .Q(n757), .DIN1(n678), .DIN2(n755) );
    nnd2s1 U249 ( .Q(n675), .DIN1(n757), .DIN2(n756) );
    nnd2s1 U250 ( .Q(n758), .DIN1(n440), .DIN2(N76) );
    nnd2s1 U251 ( .Q(n759), .DIN1(n440), .DIN2(N49) );
    nnd2s1 U252 ( .Q(n583), .DIN1(N37), .DIN2(n682) );
    nnd2s1 U253 ( .Q(n582), .DIN1(N34), .DIN2(n681) );
    nnd2s1 U254 ( .Q(n448), .DIN1(N43), .DIN2(n684) );
    nnd2s1 U255 ( .Q(n447), .DIN1(N28), .DIN2(n683) );
    nor2s1 U256 ( .Q(n451), .DIN1(n685), .DIN2(n446) );
    nor2s1 U257 ( .Q(n450), .DIN1(n760), .DIN2(N46) );
    nor2s1 U258 ( .Q(n586), .DIN1(n761), .DIN2(n762) );
    nor2s1 U259 ( .Q(n585), .DIN1(n449), .DIN2(N31) );
    nnd2s1 U260 ( .Q(n763), .DIN1(n581), .DIN2(n584) );
    nor2s1 U261 ( .Q(n453), .DIN1(n584), .DIN2(n581) );
    hi1s1 U262 ( .Q(n720), .DIN(n452) );
    nnd2s1 U263 ( .Q(n589), .DIN1(N19), .DIN2(n687) );
    nnd2s1 U264 ( .Q(n588), .DIN1(N16), .DIN2(n686) );
    nor2s1 U265 ( .Q(n457), .DIN1(n688), .DIN2(n587) );
    nnd2s1 U266 ( .Q(n764), .DIN1(n587), .DIN2(n688) );
    hi1s1 U267 ( .Q(n765), .DIN(n455) );
    nnd2s1 U268 ( .Q(n460), .DIN1(n720), .DIN2(n455) );
    nnd2s1 U269 ( .Q(n459), .DIN1(n765), .DIN2(n452) );
    nnd2s1 U270 ( .Q(n612), .DIN1(N25), .DIN2(n689) );
    nnd2s1 U271 ( .Q(n611), .DIN1(n766), .DIN2(n767) );
    nnd2s1 U272 ( .Q(n606), .DIN1(N22), .DIN2(n691) );
    nnd2s1 U273 ( .Q(n605), .DIN1(N10), .DIN2(n690) );
    nnd2s1 U274 ( .Q(n594), .DIN1(N7), .DIN2(n693) );
    nnd2s1 U275 ( .Q(n593), .DIN1(N4), .DIN2(n692) );
    nor2s1 U276 ( .Q(n486), .DIN1(n694), .DIN2(n592) );
    nnd2s1 U277 ( .Q(n768), .DIN1(n592), .DIN2(n694) );
    hi1s1 U278 ( .Q(n769), .DIN(n484) );
    nnd2s1 U279 ( .Q(n609), .DIN1(n765), .DIN2(n484) );
    nnd2s1 U280 ( .Q(n608), .DIN1(n769), .DIN2(n455) );
    nor2s1 U281 ( .Q(n770), .DIN1(n771), .DIN2(n607) );
    nnd2s1 U282 ( .Q(n493), .DIN1(n607), .DIN2(n771) );
    nor2s1 U283 ( .Q(n615), .DIN1(n449), .DIN2(n492) );
    nor2s1 U284 ( .Q(n614), .DIN1(n772), .DIN2(n762) );
    nnd2s1 U285 ( .Q(n773), .DIN1(n610), .DIN2(n613) );
    nor2s1 U286 ( .Q(n496), .DIN1(n613), .DIN2(n610) );
    nnd2s1 U287 ( .Q(n774), .DIN1(n695), .DIN2(n696) );
    nor2s1 U288 ( .Q(n498), .DIN1(n696), .DIN2(n695) );
    nnd2s1 U289 ( .Q(n597), .DIN1(N40), .DIN2(n691) );
    nnd2s1 U290 ( .Q(n596), .DIN1(N10), .DIN2(n698) );
    nor2s1 U291 ( .Q(n600), .DIN1(n699), .DIN2(n595) );
    nnd2s1 U292 ( .Q(n775), .DIN1(n595), .DIN2(n699) );
    nnd2s1 U293 ( .Q(n603), .DIN1(n720), .DIN2(n484) );
    nnd2s1 U294 ( .Q(n602), .DIN1(n769), .DIN2(n452) );
    nor2s1 U295 ( .Q(n489), .DIN1(n598), .DIN2(n601) );
    nnd2s1 U296 ( .Q(n776), .DIN1(n601), .DIN2(n598) );
    hi1s1 U297 ( .Q(n701), .DIN(n487) );
    nnd2s1 U298 ( .Q(n491), .DIN1(N76), .DIN2(n700) );
    nor2s1 U299 ( .Q(n777), .DIN1(n700), .DIN2(N76) );
    nor2s1 U300 ( .Q(n543), .DIN1(n683), .DIN2(N31) );
    nor2s1 U301 ( .Q(n542), .DIN1(n761), .DIN2(N43) );
    nnd2s1 U302 ( .Q(n546), .DIN1(N22), .DIN2(n688) );
    nnd2s1 U303 ( .Q(n545), .DIN1(N13), .DIN2(n690) );
    nor2s1 U304 ( .Q(n549), .DIN1(n541), .DIN2(n544) );
    nnd2s1 U305 ( .Q(n778), .DIN1(n544), .DIN2(n541) );
    nor2s1 U306 ( .Q(n463), .DIN1(n698), .DIN2(N25) );
    nor2s1 U307 ( .Q(n462), .DIN1(n767), .DIN2(N40) );
    hi1s1 U308 ( .Q(n718), .DIN(n461) );
    nnd2s1 U309 ( .Q(n466), .DIN1(N46), .DIN2(n461) );
    nnd2s1 U310 ( .Q(n465), .DIN1(n718), .DIN2(n685) );
    nnd2s1 U311 ( .Q(n779), .DIN1(N4), .DIN2(n702) );
    nor2s1 U312 ( .Q(n551), .DIN1(n702), .DIN2(N4) );
    nnd2s1 U313 ( .Q(n555), .DIN1(n464), .DIN2(n550) );
    nor2s1 U314 ( .Q(n780), .DIN1(n550), .DIN2(n464) );
    nor2s1 U315 ( .Q(n781), .DIN1(n547), .DIN2(n553) );
    nnd2s1 U316 ( .Q(n468), .DIN1(n553), .DIN2(n547) );
    nnd2s1 U317 ( .Q(n471), .DIN1(N82), .DIN2(n703) );
    nor2s1 U318 ( .Q(n782), .DIN1(n703), .DIN2(N82) );
    hi1s1 U319 ( .Q(n414), .DIN(n422) );
    nnd2s1 U320 ( .Q(n559), .DIN1(N34), .DIN2(n690) );
    nnd2s1 U321 ( .Q(n558), .DIN1(N22), .DIN2(n682) );
    nor2s1 U322 ( .Q(n783), .DIN1(n687), .DIN2(n557) );
    nnd2s1 U323 ( .Q(n561), .DIN1(n557), .DIN2(n687) );
    nnd2s1 U324 ( .Q(n784), .DIN1(N7), .DIN2(n704) );
    nor2s1 U325 ( .Q(n564), .DIN1(n704), .DIN2(N7) );
    nnd2s1 U326 ( .Q(n785), .DIN1(n446), .DIN2(n563) );
    nor2s1 U327 ( .Q(n567), .DIN1(n563), .DIN2(n446) );
    nnd2s1 U328 ( .Q(n474), .DIN1(n560), .DIN2(n566) );
    nor2s1 U329 ( .Q(n786), .DIN1(n566), .DIN2(n560) );
    nnd2s1 U330 ( .Q(n787), .DIN1(N85), .DIN2(n705) );
    nor2s1 U331 ( .Q(n475), .DIN1(n705), .DIN2(N85) );
    nnd2s1 U332 ( .Q(n571), .DIN1(N37), .DIN2(n684) );
    nnd2s1 U333 ( .Q(n570), .DIN1(N28), .DIN2(n681) );
    nor2s1 U334 ( .Q(n788), .DIN1(n686), .DIN2(n569) );
    nnd2s1 U335 ( .Q(n573), .DIN1(n569), .DIN2(n686) );
    nnd2s1 U336 ( .Q(n789), .DIN1(N10), .DIN2(n706) );
    nor2s1 U337 ( .Q(n576), .DIN1(n706), .DIN2(N10) );
    nnd2s1 U338 ( .Q(n790), .DIN1(n464), .DIN2(n575) );
    nor2s1 U339 ( .Q(n579), .DIN1(n575), .DIN2(n464) );
    nnd2s1 U340 ( .Q(n479), .DIN1(n572), .DIN2(n578) );
    nor2s1 U341 ( .Q(n791), .DIN1(n578), .DIN2(n572) );
    nnd2s1 U342 ( .Q(n481), .DIN1(n792), .DIN2(n709) );
    nnd2s1 U343 ( .Q(n480), .DIN1(n793), .DIN2(n707) );
    hi1s1 U344 ( .Q(n409), .DIN(n420) );
    nor2s1 U345 ( .Q(n445), .DIN1(n710), .DIN2(N1) );
    nnd2s1 U346 ( .Q(n794), .DIN1(N1), .DIN2(n710) );
    nnd2s1 U347 ( .Q(n795), .DIN1(n796), .DIN2(n797) );
    nnd2s1 U348 ( .Q(n798), .DIN1(n458), .DIN2(n443) );
    nnd2s1 U349 ( .Q(n712), .DIN1(n798), .DIN2(n795) );
    nnd2s1 U350 ( .Q(n799), .DIN1(N79), .DIN2(n711) );
    nor2s1 U351 ( .Q(n482), .DIN1(n711), .DIN2(N79) );
    nor2s1 U352 ( .Q(n667), .DIN1(n713), .DIN2(n796) );
    nnd2s1 U353 ( .Q(n800), .DIN1(n796), .DIN2(n713) );
    nor2s1 U354 ( .Q(n801), .DIN1(n722), .DIN2(n723) );
    nnd2s1 U355 ( .Q(n669), .DIN1(n723), .DIN2(n722) );
    nor2s1 U356 ( .Q(n802), .DIN1(n725), .DIN2(n668) );
    nnd2s1 U357 ( .Q(n500), .DIN1(n668), .DIN2(n725) );
    nor2s1 U358 ( .Q(n803), .DIN1(n727), .DIN2(n728) );
    nnd2s1 U359 ( .Q(n672), .DIN1(n728), .DIN2(n727) );
    nor2s1 U360 ( .Q(n804), .DIN1(n730), .DIN2(n671) );
    nnd2s1 U361 ( .Q(n502), .DIN1(n671), .DIN2(n730) );
    nnd2s1 U362 ( .Q(n537), .DIN1(n487), .DIN2(n758) );
    nor2s1 U363 ( .Q(n805), .DIN1(n758), .DIN2(n487) );
    nnd2s1 U364 ( .Q(n539), .DIN1(n495), .DIN2(n759) );
    nor2s1 U365 ( .Q(n806), .DIN1(n759), .DIN2(n495) );
    nor2s1 U366 ( .Q(n807), .DIN1(n631), .DIN2(N40) );
    nnd2s1 U367 ( .Q(n504), .DIN1(N40), .DIN2(n631) );
    nor2s1 U368 ( .Q(n808), .DIN1(n630), .DIN2(N37) );
    nnd2s1 U369 ( .Q(n506), .DIN1(N37), .DIN2(n630) );
    nor2s1 U370 ( .Q(n809), .DIN1(n634), .DIN2(N34) );
    nnd2s1 U371 ( .Q(n508), .DIN1(N34), .DIN2(n634) );
    nnd2s1 U372 ( .Q(n511), .DIN1(n810), .DIN2(n761) );
    nnd2s1 U373 ( .Q(n510), .DIN1(N31), .DIN2(n633) );
    nnd2s1 U374 ( .Q(n513), .DIN1(n811), .DIN2(n767) );
    nnd2s1 U375 ( .Q(n512), .DIN1(N25), .DIN2(n637) );
    nor2s1 U376 ( .Q(n812), .DIN1(n655), .DIN2(N22) );
    nnd2s1 U377 ( .Q(n514), .DIN1(N22), .DIN2(n655) );
    nor2s1 U378 ( .Q(n813), .DIN1(n654), .DIN2(N19) );
    nnd2s1 U379 ( .Q(n516), .DIN1(N19), .DIN2(n654) );
    nor2s1 U380 ( .Q(n814), .DIN1(n658), .DIN2(N16) );
    nnd2s1 U381 ( .Q(n518), .DIN1(N16), .DIN2(n658) );
    nnd2s1 U382 ( .Q(n521), .DIN1(n744), .DIN2(n688) );
    nnd2s1 U383 ( .Q(n520), .DIN1(N13), .DIN2(n657) );
    nor2s1 U384 ( .Q(n815), .DIN1(n636), .DIN2(N46) );
    nnd2s1 U385 ( .Q(n522), .DIN1(N46), .DIN2(n636) );
    nnd2s1 U386 ( .Q(n525), .DIN1(n745), .DIN2(n683) );
    nnd2s1 U387 ( .Q(n524), .DIN1(N43), .DIN2(n640) );
    nor2s1 U388 ( .Q(n816), .DIN1(n639), .DIN2(N28) );
    nnd2s1 U389 ( .Q(n526), .DIN1(N28), .DIN2(n639) );
    nor2s1 U390 ( .Q(n817), .DIN1(n661), .DIN2(N10) );
    nnd2s1 U391 ( .Q(n528), .DIN1(N10), .DIN2(n661) );
    nor2s1 U392 ( .Q(n818), .DIN1(n660), .DIN2(N7) );
    nnd2s1 U393 ( .Q(n530), .DIN1(N7), .DIN2(n660) );
    nor2s1 U394 ( .Q(n819), .DIN1(n664), .DIN2(N4) );
    nnd2s1 U395 ( .Q(n532), .DIN1(N4), .DIN2(n664) );
    nor2s1 U396 ( .Q(n820), .DIN1(n663), .DIN2(N1) );
    nnd2s1 U397 ( .Q(n534), .DIN1(N1), .DIN2(n663) );
    hi1s1 U398 ( .Q(n599), .DIN(n775) );
    hi1s1 U399 ( .Q(n497), .DIN(n773) );
    hi1s1 U400 ( .Q(n680), .DIN(n441) );
    hi1s1 U401 ( .Q(n724), .DIN(n721) );
    hi1s1 U402 ( .Q(n538), .DIN(n806) );
    hi1s1 U403 ( .Q(n418), .DIN(n415) );
    hi1s1 U404 ( .Q(n645), .DIN(n411) );
    hi1s1 U405 ( .Q(n678), .DIN(n428) );
    hi1s1 U406 ( .Q(n554), .DIN(n780) );
    hi1s1 U407 ( .Q(n469), .DIN(n781) );
    hi1s1 U408 ( .Q(n473), .DIN(n786) );
    hi1s1 U409 ( .Q(n499), .DIN(n774) );
    hi1s1 U410 ( .Q(n402), .DIN(n429) );
    hi1s1 U411 ( .Q(n617), .DIN(n423) );
    hi1s1 U412 ( .Q(n501), .DIN(n802) );
    hi1s1 U413 ( .Q(n503), .DIN(n804) );
    hi1s1 U414 ( .Q(n739), .DIN(n738) );
    hi1s1 U415 ( .Q(n743), .DIN(n742) );
    hi1s1 U416 ( .Q(n548), .DIN(n778) );
    hi1s1 U417 ( .Q(n670), .DIN(n801) );
    hi1s1 U418 ( .Q(n673), .DIN(n803) );
    hi1s1 U419 ( .Q(n580), .DIN(n790) );
    hi1s1 U420 ( .Q(n483), .DIN(n799) );
    hi1s1 U421 ( .Q(n761), .DIN(N31) );
    hi1s1 U422 ( .Q(n760), .DIN(n446) );
    hi1s1 U423 ( .Q(n797), .DIN(n458) );
    hi1s1 U424 ( .Q(n796), .DIN(n443) );
    hi1s1 U425 ( .Q(n735), .DIN(n734) );
    hi1s1 U426 ( .Q(n444), .DIN(n794) );
    hi1s1 U427 ( .Q(n577), .DIN(n789) );
    hi1s1 U428 ( .Q(n767), .DIN(N25) );
    hi1s1 U429 ( .Q(n574), .DIN(n788) );
    hi1s1 U430 ( .Q(n478), .DIN(n791) );
    hi1s1 U431 ( .Q(n793), .DIN(n709) );
    hi1s1 U432 ( .Q(n792), .DIN(n707) );
    hi1s1 U433 ( .Q(n456), .DIN(n764) );
    hi1s1 U434 ( .Q(n762), .DIN(n449) );
    hi1s1 U435 ( .Q(n454), .DIN(n763) );
    hi1s1 U436 ( .Q(n552), .DIN(n779) );
    hi1s1 U437 ( .Q(n470), .DIN(n782) );
    hi1s1 U438 ( .Q(n565), .DIN(n784) );
    hi1s1 U439 ( .Q(n568), .DIN(n785) );
    hi1s1 U440 ( .Q(n562), .DIN(n783) );
    hi1s1 U441 ( .Q(n476), .DIN(n787) );
    hi1s1 U442 ( .Q(n485), .DIN(n768) );
    hi1s1 U443 ( .Q(n488), .DIN(n776) );
    hi1s1 U444 ( .Q(n490), .DIN(n777) );
    hi1s1 U445 ( .Q(n771), .DIN(n604) );
    hi1s1 U446 ( .Q(n494), .DIN(n770) );
    hi1s1 U447 ( .Q(n772), .DIN(n492) );
    hi1s1 U448 ( .Q(n766), .DIN(n689) );
    hi1s1 U449 ( .Q(n405), .DIN(n424) );
    hi1s1 U450 ( .Q(n666), .DIN(n800) );
    hi1s1 U451 ( .Q(n716), .DIN(n714) );
    hi1s1 U452 ( .Q(n536), .DIN(n805) );
    hi1s1 U453 ( .Q(n505), .DIN(n807) );
    hi1s1 U454 ( .Q(n507), .DIN(n808) );
    hi1s1 U455 ( .Q(n509), .DIN(n809) );
    hi1s1 U456 ( .Q(n810), .DIN(n633) );
    hi1s1 U457 ( .Q(n811), .DIN(n637) );
    hi1s1 U458 ( .Q(n515), .DIN(n812) );
    hi1s1 U459 ( .Q(n517), .DIN(n813) );
    hi1s1 U460 ( .Q(n519), .DIN(n814) );
    hi1s1 U461 ( .Q(n523), .DIN(n815) );
    hi1s1 U462 ( .Q(n527), .DIN(n816) );
    hi1s1 U463 ( .Q(n529), .DIN(n817) );
    hi1s1 U464 ( .Q(n531), .DIN(n818) );
    hi1s1 U465 ( .Q(n533), .DIN(n819) );
    hi1s1 U466 ( .Q(n535), .DIN(n820) );
endmodule

