
module s15850 ( CK, g100, g101, g102, g103, g10377, g10379, g104, 
        g10455, g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109, 
        g11163, g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185, 
        g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700, g18, 
        g1957, g1960, g1961, g23, g2355, g2601, g2602, g2603, g2604, g2605, 
        g2606, g2607, g2608, g2609, g2610, g2611, g2612, g2648, g27, g28, g29, 
        g2986, g30, g3007, g3069, g31, g3327, g41, g4171, g4172, g4173, g4174, 
        g4175, g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, 
        g4194, g4195, g4196, g4197, g4198, g4199, g42, g4200, g4201, g4202, 
        g4203, g4204, g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, 
        g4213, g4214, g4215, g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, 
        g5101, g5105, g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, 
        g6258, g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267, 
        g6268, g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276, g6277, 
        g6278, g6279, g6280, g6281, g6282, g6283, g6284, g6285, g6842, g6920, 
        g6926, g6932, g6942, g6949, g6955, g741, g742, g743, g744, g750, g7744, 
        g8061, g8062, g82, g8271, g83, g8313, g8316, g8318, g8323, g8328, 
        g8331, g8335, g8340, g8347, g8349, g8352, g84, g85, g8561, g8562, 
        g8563, g8564, g8565, g8566, g86, g87, g872, g873, g877, g88, g881, 
        g886, g889, g89, g892, g895, g8976, g8977, g8978, g8979, g898, g8980, 
        g8981, g8982, g8983, g8984, g8985, g8986, g90, g901, g904, g907, g91, 
        g910, g913, g916, g919, g92, g922, g925, g93, g94, g9451, g95, g96, 
        g99, g9961 );
  input  CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176,
         g1179, g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696,
         g1700, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41,
         g42, g43, g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82,
         g83, g84, g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89,
         g892, g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919,
         g92, g922, g925, g93, g94, g95, g96, g99;
  output g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
         g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601, g2602,
         g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612,
         g2648, g2986, g3007, g3069, g3327, g4171, g4172, g4173, g4174, g4175,
         g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194,
         g4195, g4196, g4197, g4198, g4199, g4200, g4201, g4202, g4203, g4204,
         g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214,
         g4215, g4216, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253,
         g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
         g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
         g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
         g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g7744,
         g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335,
         g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566,
         g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985,
         g8986, g9451, g9961;
  wire   g100, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, g1194,
         g1197, g1200, g1203, g18, g1960, g1961, g27, g30, g31, g41, g42, g43,
         g44, g45, g46, g47, g48, g82, g84, g85, g86, g87, g872, g873, g88,
         g886, g889, g89, g892, g895, g898, g90, g901, g904, g907, g91, g910,
         g913, g916, g919, g92, g922, g925, g93, g94, g95, g96, g99, g1289,
         g5660, g1882, g9349, g312, g5644, g452, g11257, g123, g8272, g207,
         g7315, g713, g9345, g1153, g6304, g1744, g5663, g1558, g7349, g695,
         g9343, g461, g11467, g940, g8572, g976, g11471, g709, g8432, g1092,
         g6810, g1574, g7354, g7816, g369, g11439, g1580, g7356, g1736, g6846,
         g39, g10774, g11182, g1424, g7330, g1737, g1672, g11037, g1077, g6805,
         g1231, g8279, g4, g8079, g774, g7785, g1104, g6815, g1304, g7290,
         g243, g7325, g1499, g8447, g1444, g8987, g757, g11179, g786, g8436,
         g1543, g7344, g315, g5645, g1534, g7341, g622, g9338, g1927, g9354,
         g1660, g11033, g278, g7765, g1436, g8989, g718, g8433, g7775, g554,
         g11047, g496, g11333, g981, g11472, g4896, g590, g5653, g829, g4182,
         g1095, g6811, g704, g9344, g1265, g7302, g1786, g7814, g682, g8429,
         g1296, g7292, g587, g6295, g7777, g646, g8065, g327, g5649, g1389,
         g6836, g7311, g1956, g1955, g1675, g11038, g354, g11508, g113, g7285,
         g639, g8063, g1684, g11041, g1639, g8448, g1791, g8080, g248, g7323,
         g1707, g4907, g1759, g5668, g351, g11507, g1604, g7364, g1098, g6812,
         g932, g8570, g1896, g8282, g736, g8435, g1019, g7807, g1362, g7305,
         g745, g2639, g1419, g7332, g7779, g11397, g1086, g6808, g1486, g8444,
         g1730, g10881, g1504, g7328, g1470, g8440, g8437, g583, g1678, g11039,
         g174, g8423, g1766, g7810, g1801, g8450, g186, g7317, g959, g11403,
         g1007, g7806, g1407, g8993, g1868, g7817, g758, g6797, g1718, g6337,
         g396, g11265, g1015, g7808, g38, g10872, g632, g5655, g1415, g7335,
         g1227, g8278, g1721, g10878, g16, g4906, g284, g7767, g426, g11256,
         g219, g7310, g1360, g7289, g1428, g8992, g579, g1564, g7351, g1741,
         g5662, g225, g7309, g281, g7766, g1308, g11627, g611, g9930, g5654,
         g1217, g9823, g1589, g7359, g1466, g8439, g1571, g7353, g1861, g7815,
         g1365, g7307, g1448, g11594, g1133, g6309, g1333, g11635, g153, g8426,
         g962, g11404, g766, g6799, g588, g6296, g486, g11331, g471, g11469,
         g1397, g7322, g580, g1950, g8288, g755, g5656, g1101, g6814, g549,
         g11044, g105, g11180, g1669, g11036, g7308, g1531, g7340, g1458,
         g7327, g572, g10877, g1011, g7805, g10867, g1411, g7331, g1074, g6813,
         g444, g11259, g1474, g8441, g1080, g6806, g6336, g333, g5651, g269,
         g7762, g401, g11266, g1857, g11409, g9, g7336, g664, g8782, g965,
         g11405, g7324, g309, g5652, g8077, g231, g7319, g557, g11048, g586,
         g6294, g869, g875, g7316, g158, g8425, g5657, g1023, g7799, g7755,
         g1327, g11633, g654, g8067, g293, g7770, g1346, g11656, g1633, g8873,
         g1753, g5666, g1508, g7329, g1240, g7297, g538, g11326, g416, g11269,
         g542, g11325, g1681, g11040, g374, g11440, g563, g11050, g1914, g8284,
         g530, g11328, g575, g11052, g1936, g9355, g7778, g1117, g6299, g1317,
         g1356, g357, g11509, g386, g11263, g1601, g7363, g166, g7747, g501,
         g11334, g7758, g1840, g8694, g7783, g318, g5646, g6818, g6800, g10870,
         g302, g7773, g342, g11513, g1250, g7299, g6301, g2044, g1032, g7800,
         g1432, g8990, g1453, g7326, g363, g11511, g330, g5650, g6303, g1357,
         g6330, g10869, g928, g8569, g7757, g516, g11337, g7759, g778, g8076,
         g861, g4190, g1627, g8871, g1292, g7293, g290, g7769, g1850, g5671,
         g770, g7288, g1583, g7357, g466, g11468, g1561, g7350, g1546, g7345,
         g287, g7768, g560, g11049, g617, g8780, g17, g4894, g336, g11653,
         g456, g11466, g305, g5643, g345, g11642, g8, g2613, g1771, g7811,
         g865, g8275, g7751, g1945, g9356, g1738, g5661, g1478, g8442, g4217,
         g1690, g6844, g1482, g8443, g1110, g6817, g296, g7771, g1663, g11034,
         g700, g8431, g1762, g5669, g360, g11510, g192, g6837, g1657, g10875,
         g722, g9346, g7780, g566, g11051, g7809, g1089, g6809, g4897, g1071,
         g6804, g986, g11473, g971, g11470, g6338, g143, g7746, g1814, g9825,
         g1212, g1918, g9353, g782, g8273, g1822, g9826, g237, g7306, g2638,
         g1462, g8438, g178, g7748, g366, g11512, g837, g4184, g599, g9819,
         g11408, g944, g11398, g1941, g8287, g170, g8422, g1520, g7334, g686,
         g9342, g953, g11401, g6339, g10775, g1765, g3329, g1733, g10882,
         g1270, g7303, g1610, g6845, g1796, g8280, g1324, g11632, g1540, g7343,
         g7312, g4898, g491, g11332, g5670, g213, g7313, g1781, g7813, g1900,
         g9351, g1245, g7298, g108, g11593, g7287, g148, g8427, g833, g4183,
         g1923, g8285, g936, g8571, g1314, g11629, g849, g4187, g1336, g11654,
         g272, g7763, g1806, g8573, g8568, g1887, g8281, g37, g10871, g968,
         g11406, g5673, g1137, g6310, g1891, g9350, g1255, g7300, g7753, g874,
         g9821, g591, g9818, g731, g9347, g8781, g1218, g8276, g605, g9820,
         g7776, g182, g7749, g950, g11400, g1129, g6308, g857, g4189, g448,
         g11258, g1828, g9827, g1727, g10880, g1592, g7360, g1703, g6843,
         g1932, g8286, g1624, g8870, g1068, g6803, g578, g440, g11260, g476,
         g11338, g119, g7745, g668, g9340, g139, g8418, g1149, g6305, g10868,
         g7366, g263, g7760, g8274, g1747, g5664, g6802, g275, g7764, g1524,
         g7338, g1577, g7355, g7786, g391, g11264, g658, g9339, g1386, g7318,
         g7750, g9822, g1125, g6307, g201, g7304, g1280, g7295, g1083, g6807,
         g8066, g1636, g8874, g853, g4188, g421, g11270, g762, g6798, g956,
         g11402, g378, g11441, g1756, g5667, g589, g6297, g841, g4185, g1027,
         g7798, g1003, g7803, g1403, g8991, g1145, g6312, g1107, g6816, g1223,
         g8277, g406, g11267, g1811, g11185, g11183, g1654, g10874, g6835,
         g1595, g7361, g1537, g7342, g727, g8434, g999, g7804, g6801, g481,
         g11324, g754, g4895, g1330, g11634, g845, g4186, g790, g8567, g1512,
         g8449, g1490, g8445, g6300, g348, g11506, g1260, g7301, g7756, g131,
         g8420, g7, g2731, g7754, g521, g11330, g1318, g11630, g1872, g9348,
         g677, g9341, g582, g7320, g1549, g7346, g947, g11399, g1834, g9895,
         g1598, g7362, g1121, g6306, g1321, g11631, g506, g11335, g546, g11043,
         g1909, g9352, g1552, g7347, g584, g6292, g1687, g11042, g1586, g7358,
         g324, g5648, g1141, g6311, g1341, g11655, g1710, g4901, g11184, g7321,
         g135, g8419, g525, g11329, g581, g1607, g7365, g321, g5647, g7782,
         g1275, g11443, g1311, g11628, g1615, g8868, g382, g11442, g6825, g266,
         g7761, g1284, g7294, g7314, g673, g8428, g5672, g162, g8424, g411,
         g11268, g431, g11262, g1905, g8283, g1515, g7333, g1630, g8872, g7774,
         g991, g7802, g1300, g7291, g339, g11505, g7752, g1750, g5665, g585,
         g6293, g1440, g8988, g1666, g11035, g1528, g7339, g1351, g11657,
         g11181, g127, g8421, g1618, g11611, g1235, g7296, g299, g7772, g435,
         g11261, g7781, g1555, g7348, g995, g7801, g1621, g8869, g6313, g643,
         g8064, g1494, g8446, g1567, g7352, g691, g8430, g534, g11327, g1776,
         g7812, g569, g10876, g6302, g9824, g1, g8078, g511, g11336, g1724,
         g10879, g12, g7337, g1878, g8695, g7784, g3435, g10408, g10336, g3399,
         g8226, g8814, g10417, g9931, g8241, g10405, g8214, g8187, g3431,
         g10712, g2791, g10411, g8203, g10414, g3418, g8816, g10515, g8815,
         g10583, g3425, g6919, g10779, g3438, g3414, g8812, g10402, g8221,
         g8200, g8811, g8818, g8236, g10339, g8206, g8817, g8810, g8230, g5287,
         g8819, g3407, g8806, g8813, g8210, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, \DFF_489/net776 , \DFF_452/net739 ,
         \DFF_441/net728 , \DFF_436/net723 , \DFF_385/net672 ,
         \DFF_384/net671 , \DFF_336/net623 , \DFF_330/net617 ,
         \DFF_319/net606 , \DFF_275/net562 , \DFF_270/net557 ,
         \DFF_242/net529 , \DFF_228/net515 , \DFF_194/net481 ,
         \DFF_168/net455 , \DFF_157/net444 , \DFF_136/net423 ,
         \DFF_126/net413 , \DFF_121/net408 , \DFF_93/net380 ;
  assign g6280 = g100;
  assign g4205 = g1170;
  assign g4209 = g1173;
  assign g4210 = g1176;
  assign g4211 = g1179;
  assign g4212 = g1182;
  assign g4213 = g1185;
  assign g4214 = g1188;
  assign g4215 = g1191;
  assign g4216 = g1194;
  assign g4206 = g1197;
  assign g4207 = g1200;
  assign g4208 = g1203;
  assign g2355 = g18;
  assign g4888 = g1960;
  assign g4887 = g1961;
  assign g7744 = g27;
  assign g6254 = g30;
  assign g6255 = g31;
  assign g6256 = g41;
  assign g6257 = g42;
  assign g6258 = g43;
  assign g6259 = g44;
  assign g6260 = g45;
  assign g6261 = g46;
  assign g6262 = g47;
  assign g6263 = g48;
  assign g6264 = g82;
  assign g6266 = g84;
  assign g6267 = g85;
  assign g6268 = g86;
  assign g6269 = g87;
  assign g8061 = g872;
  assign g5101 = g872;
  assign g8062 = g873;
  assign g5105 = g873;
  assign g6270 = g88;
  assign g4191 = g886;
  assign g4192 = g889;
  assign g6271 = g89;
  assign g4193 = g892;
  assign g4194 = g895;
  assign g4195 = g898;
  assign g6272 = g90;
  assign g4197 = g901;
  assign g4198 = g904;
  assign g4199 = g907;
  assign g6273 = g91;
  assign g4200 = g910;
  assign g4201 = g913;
  assign g4202 = g916;
  assign g4203 = g919;
  assign g6274 = g92;
  assign g4204 = g922;
  assign g4196 = g925;
  assign g6275 = g93;
  assign g6276 = g94;
  assign g6277 = g95;
  assign g6278 = g96;
  assign g6279 = g99;
  assign g4177 = g774;
  assign g4180 = g786;
  assign g2602 = g587;
  assign g6284 = g6295;
  assign g6295 = g104;
  assign g2609 = g583;
  assign g4173 = g758;
  assign g2605 = g579;
  assign g4175 = g766;
  assign g2603 = g588;
  assign g6285 = g6296;
  assign g6296 = g28;
  assign g2606 = g580;
  assign g2612 = g586;
  assign g6283 = g6294;
  assign g6294 = g103;
  assign g4178 = g778;
  assign g4176 = g770;
  assign g2648 = g865;
  assign g6265 = g6338;
  assign g6338 = g83;
  assign g4179 = g782;
  assign g2601 = g578;
  assign g4174 = g762;
  assign g2604 = g589;
  assign g6253 = g6297;
  assign g6297 = g29;
  assign g4172 = g754;
  assign g4181 = g790;
  assign g2608 = g582;
  assign g2610 = g584;
  assign g6281 = g6292;
  assign g6292 = g101;
  assign g2607 = g581;
  assign g2611 = g585;
  assign g6282 = g6293;
  assign g6293 = g102;
  assign g8565 = g3435;
  assign g6949 = g3435;
  assign g10459 = g10408;
  assign g10377 = g10336;
  assign g8561 = g3399;
  assign g6920 = g3399;
  assign g8331 = g8226;
  assign g8982 = g8814;
  assign g10465 = g10417;
  assign g9961 = g9931;
  assign g9451 = g9931;
  assign g8349 = g8241;
  assign g10457 = g10405;
  assign g8323 = g8214;
  assign g8352 = g8187;
  assign g8564 = g3431;
  assign g6942 = g3431;
  assign g10801 = g10712;
  assign g4171 = g2791;
  assign g10461 = g10411;
  assign g8313 = g8203;
  assign g10463 = g10414;
  assign g5659 = g3418;
  assign g8984 = g8816;
  assign g10628 = g10515;
  assign g8983 = g8815;
  assign g11206 = g10583;
  assign g8563 = g3425;
  assign g6932 = g3425;
  assign g8271 = g6919;
  assign g5816 = g6919;
  assign g11163 = g10779;
  assign g8566 = g3438;
  assign g6955 = g3438;
  assign g8562 = g3414;
  assign g6926 = g3414;
  assign g8980 = g8812;
  assign g10455 = g10402;
  assign g8328 = g8221;
  assign g8347 = g8200;
  assign g8979 = g8811;
  assign g8985 = g8818;
  assign g8340 = g8236;
  assign g10379 = g10339;
  assign g8316 = g8206;
  assign g8976 = g8817;
  assign g8978 = g8810;
  assign g8335 = g8230;
  assign g6842 = g5287;
  assign g8986 = g8819;
  assign g5658 = g3407;
  assign g8977 = g8806;
  assign g8981 = g8813;
  assign g8318 = g8210;
  assign g11489 = 1'b0;

  nnd2s1 U2440 ( .Q(n2656), .DIN1(n2684), .DIN2(g109) );
  hi1s1 U2441 ( .Q(n2710), .DIN(n2738) );
  hi1s1 U2442 ( .Q(n2741), .DIN(n2738) );
  or2s1 U2443 ( .Q(n2059), .DIN1(n2067), .DIN2(n2799) );
  hi1s1 U2444 ( .Q(n2060), .DIN(n2059) );
  hi1s1 U2445 ( .Q(n2062), .DIN(n2061) );
  nor2s1 U2446 ( .Q(n2063), .DIN1(g1696), .DIN2(g1703) );
  hi1s1 U2447 ( .Q(n2064), .DIN(g109) );
  hi1s1 U2448 ( .Q(n2067), .DIN(g109) );
  hi1s1 U2449 ( .Q(n2065), .DIN(g109) );
  hi1s1 U2450 ( .Q(n2066), .DIN(g109) );
  hi1s1 U2451 ( .Q(n2068), .DIN(n2063) );
  hi1s1 U2452 ( .Q(n2070), .DIN(n2063) );
  hi1s1 U2453 ( .Q(n2069), .DIN(n2350) );
  hi1s1 U2454 ( .Q(n2071), .DIN(n2079) );
  hi1s1 U2455 ( .Q(n2072), .DIN(g18) );
  hi1s1 U2456 ( .Q(n2075), .DIN(n2074) );
  or4s1 U2457 ( .Q(n2076), .DIN1(n3304), .DIN2(n2065), .DIN3(n3305), .DIN4(
        n3306) );
  hi1s1 U2458 ( .Q(n2077), .DIN(n2076) );
  hi1s1 U2459 ( .Q(n2078), .DIN(n2076) );
  hi1s1 U2460 ( .Q(n2079), .DIN(n2076) );
  or3s1 U2461 ( .Q(g9931), .DIN1(g30), .DIN2(g31), .DIN3(n2080) );
  hi1s1 U2462 ( .Q(n2080), .DIN(n2081) );
  nor2s1 U2463 ( .Q(g9930), .DIN1(n2072), .DIN2(n2083) );
  xor2s1 U2464 ( .Q(n2083), .DIN1(n2084), .DIN2(n1975) );
  nnd2s1 U2465 ( .Q(n2084), .DIN1(n2085), .DIN2(n2086) );
  nnd2s1 U2466 ( .Q(n2086), .DIN1(n2087), .DIN2(n2088) );
  nnd2s1 U2467 ( .Q(n2088), .DIN1(n1982), .DIN2(n2089) );
  nnd2s1 U2468 ( .Q(n2089), .DIN1(n2090), .DIN2(n2091) );
  and3s1 U2469 ( .Q(g9895), .DIN1(n2092), .DIN2(n2093), .DIN3(g18) );
  nnd2s1 U2470 ( .Q(n2093), .DIN1(n2094), .DIN2(n1948) );
  nnd3s1 U2471 ( .Q(n2092), .DIN1(n2095), .DIN2(n2096), .DIN3(g1834) );
  nnd2s1 U2472 ( .Q(n2096), .DIN1(n2097), .DIN2(n1983) );
  or2s1 U2473 ( .Q(n2097), .DIN1(n2098), .DIN2(n2099) );
  and3s1 U2474 ( .Q(g9827), .DIN1(n2100), .DIN2(n2101), .DIN3(g18) );
  nnd3s1 U2475 ( .Q(n2101), .DIN1(n2102), .DIN2(n2103), .DIN3(n1980) );
  or2s1 U2476 ( .Q(n2100), .DIN1(n2103), .DIN2(n1980) );
  nnd2s1 U2477 ( .Q(n2103), .DIN1(n2099), .DIN2(n2104) );
  nnd3s1 U2478 ( .Q(n2104), .DIN1(n2105), .DIN2(n2106), .DIN3(n2107) );
  nnd3s1 U2479 ( .Q(n2105), .DIN1(g1814), .DIN2(g1822), .DIN3(g1828) );
  nor2s1 U2480 ( .Q(g9826), .DIN1(n2108), .DIN2(n2082) );
  xor2s1 U2481 ( .Q(n2108), .DIN1(n2109), .DIN2(n1953) );
  nor2s1 U2482 ( .Q(n2109), .DIN1(n2110), .DIN2(n2111) );
  nor2s1 U2483 ( .Q(n2110), .DIN1(n2112), .DIN2(n2113) );
  nor2s1 U2484 ( .Q(g9825), .DIN1(n2114), .DIN2(n2072) );
  xor2s1 U2485 ( .Q(n2114), .DIN1(g1814), .DIN2(n2115) );
  nnd2s1 U2486 ( .Q(n2115), .DIN1(n2099), .DIN2(n2116) );
  nnd3s1 U2487 ( .Q(n2116), .DIN1(n2098), .DIN2(n2117), .DIN3(n2118) );
  hi1s1 U2488 ( .Q(n2117), .DIN(n2112) );
  nor2s1 U2489 ( .Q(n2112), .DIN1(n2119), .DIN2(g1822) );
  nnd3s1 U2490 ( .Q(g9824), .DIN1(n2120), .DIN2(n2121), .DIN3(g47) );
  nnd2s1 U2491 ( .Q(g9823), .DIN1(n2122), .DIN2(g47) );
  nnd4s1 U2492 ( .Q(g9822), .DIN1(g46), .DIN2(n2123), .DIN3(n2081), .DIN4(
        n2124) );
  nnd3s1 U2493 ( .Q(g9821), .DIN1(n2120), .DIN2(n2124), .DIN3(g46) );
  and4s1 U2494 ( .Q(n2120), .DIN1(n2125), .DIN2(n2126), .DIN3(n2081), .DIN4(
        n2127) );
  and3s1 U2495 ( .Q(n2127), .DIN1(n2128), .DIN2(n2129), .DIN3(n2130) );
  and3s1 U2496 ( .Q(g9820), .DIN1(n2131), .DIN2(n2132), .DIN3(g18) );
  nnd3s1 U2497 ( .Q(n2132), .DIN1(n2133), .DIN2(n2134), .DIN3(n1978) );
  nnd2s1 U2498 ( .Q(n2133), .DIN1(n2135), .DIN2(n2136) );
  nnd3s1 U2499 ( .Q(n2131), .DIN1(n2135), .DIN2(n2136), .DIN3(g605) );
  nnd3s1 U2500 ( .Q(n2136), .DIN1(n2137), .DIN2(n2138), .DIN3(n2139) );
  nnd2s1 U2501 ( .Q(n2138), .DIN1(n2140), .DIN2(g599) );
  nnd2s1 U2502 ( .Q(n2137), .DIN1(n2090), .DIN2(n1987) );
  nor2s1 U2503 ( .Q(g9819), .DIN1(n2141), .DIN2(n2082) );
  xor2s1 U2504 ( .Q(n2141), .DIN1(g599), .DIN2(n2142) );
  nnd2s1 U2505 ( .Q(n2142), .DIN1(n2135), .DIN2(n2143) );
  nnd2s1 U2506 ( .Q(n2143), .DIN1(n2144), .DIN2(n2145) );
  nor2s1 U2507 ( .Q(g9818), .DIN1(n2146), .DIN2(n2082) );
  xor2s1 U2508 ( .Q(n2146), .DIN1(g591), .DIN2(n2147) );
  nnd2s1 U2509 ( .Q(n2147), .DIN1(n2135), .DIN2(n2148) );
  nnd3s1 U2510 ( .Q(n2148), .DIN1(n2149), .DIN2(n2145), .DIN3(n2150) );
  nnd2s1 U2511 ( .Q(n2145), .DIN1(n2140), .DIN2(n1985) );
  nnd2s1 U2512 ( .Q(g9356), .DIN1(n2151), .DIN2(n2152) );
  nnd2s1 U2513 ( .Q(n2152), .DIN1(n2153), .DIN2(n2154) );
  xor2s1 U2514 ( .Q(n2154), .DIN1(n2155), .DIN2(n2008) );
  nnd3s1 U2515 ( .Q(n2155), .DIN1(n2156), .DIN2(n2157), .DIN3(n2158) );
  or2s1 U2516 ( .Q(n2157), .DIN1(n2159), .DIN2(g1950) );
  nnd3s1 U2517 ( .Q(n2156), .DIN1(n2160), .DIN2(n2161), .DIN3(n2159) );
  nnd2s1 U2518 ( .Q(g9355), .DIN1(n2151), .DIN2(n2162) );
  nnd2s1 U2519 ( .Q(n2162), .DIN1(n2153), .DIN2(n2163) );
  xor2s1 U2520 ( .Q(n2163), .DIN1(n2164), .DIN2(n1993) );
  nnd3s1 U2521 ( .Q(n2164), .DIN1(n2165), .DIN2(n2166), .DIN3(n2158) );
  or2s1 U2522 ( .Q(n2166), .DIN1(n2159), .DIN2(g1941) );
  nnd2s1 U2523 ( .Q(n2165), .DIN1(n2167), .DIN2(n2159) );
  nnd2s1 U2524 ( .Q(n2167), .DIN1(n2168), .DIN2(n2169) );
  nnd2s1 U2525 ( .Q(n2169), .DIN1(n2170), .DIN2(n1954) );
  nnd2s1 U2526 ( .Q(n2170), .DIN1(n2171), .DIN2(n2172) );
  nnd2s1 U2527 ( .Q(n2168), .DIN1(g1927), .DIN2(n2173) );
  nnd2s1 U2528 ( .Q(n2173), .DIN1(n2174), .DIN2(n2175) );
  nnd2s1 U2529 ( .Q(g9354), .DIN1(n2151), .DIN2(n2176) );
  nnd2s1 U2530 ( .Q(n2176), .DIN1(n2153), .DIN2(n2177) );
  xor2s1 U2531 ( .Q(n2177), .DIN1(n2178), .DIN2(n1954) );
  nnd2s1 U2532 ( .Q(n2178), .DIN1(n2158), .DIN2(n2179) );
  nnd3s1 U2533 ( .Q(n2179), .DIN1(n2180), .DIN2(n2181), .DIN3(n2182) );
  nnd2s1 U2534 ( .Q(n2182), .DIN1(g1932), .DIN2(n2183) );
  nnd2s1 U2535 ( .Q(n2181), .DIN1(n2184), .DIN2(n2172) );
  nnd2s1 U2536 ( .Q(n2180), .DIN1(n2185), .DIN2(n2175) );
  nnd2s1 U2537 ( .Q(g9353), .DIN1(n2151), .DIN2(n2186) );
  nnd2s1 U2538 ( .Q(n2186), .DIN1(n2153), .DIN2(n2187) );
  xor2s1 U2539 ( .Q(n2187), .DIN1(n2188), .DIN2(n2028) );
  nnd2s1 U2540 ( .Q(n2188), .DIN1(n2158), .DIN2(n2189) );
  nnd3s1 U2541 ( .Q(n2189), .DIN1(n2190), .DIN2(n2191), .DIN3(n2192) );
  nnd2s1 U2542 ( .Q(n2192), .DIN1(g1923), .DIN2(n2183) );
  nnd3s1 U2543 ( .Q(n2191), .DIN1(n2184), .DIN2(n1932), .DIN3(n1957) );
  nnd3s1 U2544 ( .Q(n2190), .DIN1(n2185), .DIN2(g1900), .DIN3(g1909) );
  nnd2s1 U2545 ( .Q(g9352), .DIN1(n2151), .DIN2(n2193) );
  nnd2s1 U2546 ( .Q(n2193), .DIN1(n2153), .DIN2(n2194) );
  xor2s1 U2547 ( .Q(n2194), .DIN1(n2195), .DIN2(n1957) );
  nnd2s1 U2548 ( .Q(n2195), .DIN1(n2158), .DIN2(n2196) );
  nnd3s1 U2549 ( .Q(n2196), .DIN1(n2197), .DIN2(n2198), .DIN3(n2199) );
  nnd2s1 U2550 ( .Q(n2199), .DIN1(g1914), .DIN2(n2183) );
  nnd2s1 U2551 ( .Q(n2198), .DIN1(n2184), .DIN2(n1932) );
  hi1s1 U2552 ( .Q(n2184), .DIN(n2200) );
  nnd2s1 U2553 ( .Q(n2197), .DIN1(n2185), .DIN2(g1900) );
  hi1s1 U2554 ( .Q(n2185), .DIN(n2201) );
  nnd2s1 U2555 ( .Q(g9351), .DIN1(n2151), .DIN2(n2202) );
  nnd2s1 U2556 ( .Q(n2202), .DIN1(n2153), .DIN2(n2203) );
  xor2s1 U2557 ( .Q(n2203), .DIN1(n2204), .DIN2(n1932) );
  nnd2s1 U2558 ( .Q(n2204), .DIN1(n2158), .DIN2(n2205) );
  nnd3s1 U2559 ( .Q(n2205), .DIN1(n2201), .DIN2(n2200), .DIN3(n2206) );
  nnd2s1 U2560 ( .Q(n2206), .DIN1(g1905), .DIN2(n2183) );
  nnd2s1 U2561 ( .Q(n2200), .DIN1(n2159), .DIN2(n2171) );
  nnd2s1 U2562 ( .Q(n2201), .DIN1(n2159), .DIN2(n2174) );
  nnd2s1 U2563 ( .Q(g9350), .DIN1(n2151), .DIN2(n2207) );
  nnd2s1 U2564 ( .Q(n2207), .DIN1(n2153), .DIN2(n2208) );
  xor2s1 U2565 ( .Q(n2208), .DIN1(n2209), .DIN2(n2010) );
  nnd3s1 U2566 ( .Q(n2209), .DIN1(n2210), .DIN2(n2211), .DIN3(n2158) );
  or2s1 U2567 ( .Q(n2211), .DIN1(n2159), .DIN2(g1896) );
  nnd2s1 U2568 ( .Q(n2210), .DIN1(n2159), .DIN2(n2212) );
  nnd3s1 U2569 ( .Q(n2212), .DIN1(n2213), .DIN2(n2214), .DIN3(n2215) );
  nnd2s1 U2570 ( .Q(n2215), .DIN1(g1882), .DIN2(n2216) );
  nnd2s1 U2571 ( .Q(n2214), .DIN1(n2217), .DIN2(n1956) );
  nnd2s1 U2572 ( .Q(n2213), .DIN1(g1872), .DIN2(n1935) );
  nnd2s1 U2573 ( .Q(g9349), .DIN1(n2151), .DIN2(n2218) );
  nnd2s1 U2574 ( .Q(n2218), .DIN1(n2153), .DIN2(n2219) );
  xor2s1 U2575 ( .Q(n2219), .DIN1(n2220), .DIN2(n1935) );
  nnd3s1 U2576 ( .Q(n2220), .DIN1(n2221), .DIN2(n2222), .DIN3(n2158) );
  hi1s1 U2577 ( .Q(n2158), .DIN(n2223) );
  or2s1 U2578 ( .Q(n2222), .DIN1(n2159), .DIN2(g1887) );
  nnd2s1 U2579 ( .Q(n2221), .DIN1(n2224), .DIN2(n2159) );
  xor2s1 U2580 ( .Q(n2224), .DIN1(n1956), .DIN2(n2216) );
  nnd2s1 U2581 ( .Q(g9348), .DIN1(n2151), .DIN2(n2225) );
  nnd2s1 U2582 ( .Q(n2225), .DIN1(n2153), .DIN2(n2226) );
  xor2s1 U2583 ( .Q(n2226), .DIN1(g1872), .DIN2(n2227) );
  nor2s1 U2584 ( .Q(n2227), .DIN1(n2228), .DIN2(n2223) );
  nor2s1 U2585 ( .Q(n2223), .DIN1(n2183), .DIN2(n2229) );
  nor2s1 U2586 ( .Q(n2228), .DIN1(g1878), .DIN2(n2159) );
  hi1s1 U2587 ( .Q(n2159), .DIN(n2183) );
  nnd2s1 U2588 ( .Q(n2183), .DIN1(n2230), .DIN2(n2094) );
  nnd2s1 U2589 ( .Q(n2094), .DIN1(n2095), .DIN2(g1840) );
  nnd4s1 U2590 ( .Q(n2151), .DIN1(n2231), .DIN2(n2102), .DIN3(n2098), .DIN4(
        n2232) );
  hi1s1 U2591 ( .Q(n2232), .DIN(n2153) );
  nor2s1 U2592 ( .Q(n2153), .DIN1(n2233), .DIN2(n2099) );
  hi1s1 U2593 ( .Q(n2099), .DIN(n2111) );
  nnd3s1 U2594 ( .Q(n2111), .DIN1(n2234), .DIN2(n2235), .DIN3(n2229) );
  and2s1 U2595 ( .Q(n2229), .DIN1(n2095), .DIN2(n2236) );
  nnd2s1 U2596 ( .Q(n2236), .DIN1(n2237), .DIN2(n2098) );
  or2s1 U2597 ( .Q(n2237), .DIN1(n1989), .DIN2(n2238) );
  nnd2s1 U2598 ( .Q(n2235), .DIN1(g1945), .DIN2(n2161) );
  nnd4s1 U2599 ( .Q(n2161), .DIN1(g1936), .DIN2(g1927), .DIN3(n2174), .DIN4(
        n2175) );
  and3s1 U2600 ( .Q(n2175), .DIN1(g1909), .DIN2(g1900), .DIN3(g1918) );
  and4s1 U2601 ( .Q(n2174), .DIN1(g1891), .DIN2(g1882), .DIN3(g1872), .DIN4(
        n2217) );
  nnd2s1 U2602 ( .Q(n2234), .DIN1(n2160), .DIN2(n2008) );
  nnd4s1 U2603 ( .Q(n2160), .DIN1(n2171), .DIN2(n2172), .DIN3(n1954), .DIN4(
        n1993) );
  and3s1 U2604 ( .Q(n2172), .DIN1(n1957), .DIN2(n2028), .DIN3(n1932) );
  and4s1 U2605 ( .Q(n2171), .DIN1(n2216), .DIN2(n1956), .DIN3(n1935), .DIN4(
        n2010) );
  hi1s1 U2606 ( .Q(n2216), .DIN(n2217) );
  nnd2s1 U2607 ( .Q(n2217), .DIN1(g1822), .DIN2(n2106) );
  nnd2s1 U2608 ( .Q(n2106), .DIN1(n2239), .DIN2(n1980) );
  nnd3s1 U2609 ( .Q(n2098), .DIN1(g1814), .DIN2(n1983), .DIN3(g1834) );
  nnd2s1 U2610 ( .Q(g9347), .DIN1(n2240), .DIN2(n2241) );
  nnd2s1 U2611 ( .Q(n2241), .DIN1(n2242), .DIN2(n2243) );
  xor2s1 U2612 ( .Q(n2243), .DIN1(n2244), .DIN2(n2009) );
  nnd3s1 U2613 ( .Q(n2244), .DIN1(n2245), .DIN2(n2246), .DIN3(n2247) );
  or2s1 U2614 ( .Q(n2246), .DIN1(n2248), .DIN2(g736) );
  nnd3s1 U2615 ( .Q(n2245), .DIN1(n2249), .DIN2(n2250), .DIN3(n2248) );
  nnd2s1 U2616 ( .Q(g9346), .DIN1(n2240), .DIN2(n2251) );
  nnd2s1 U2617 ( .Q(n2251), .DIN1(n2242), .DIN2(n2252) );
  xor2s1 U2618 ( .Q(n2252), .DIN1(n2253), .DIN2(n1994) );
  nnd3s1 U2619 ( .Q(n2253), .DIN1(n2254), .DIN2(n2255), .DIN3(n2247) );
  or2s1 U2620 ( .Q(n2255), .DIN1(n2248), .DIN2(g727) );
  nnd2s1 U2621 ( .Q(n2254), .DIN1(n2256), .DIN2(n2248) );
  nnd2s1 U2622 ( .Q(n2256), .DIN1(n2257), .DIN2(n2258) );
  nnd2s1 U2623 ( .Q(n2258), .DIN1(n2259), .DIN2(n1955) );
  nnd2s1 U2624 ( .Q(n2259), .DIN1(n2260), .DIN2(n2261) );
  nnd2s1 U2625 ( .Q(n2257), .DIN1(g713), .DIN2(n2262) );
  nnd2s1 U2626 ( .Q(n2262), .DIN1(n2263), .DIN2(n2264) );
  nnd2s1 U2627 ( .Q(g9345), .DIN1(n2240), .DIN2(n2265) );
  nnd2s1 U2628 ( .Q(n2265), .DIN1(n2242), .DIN2(n2266) );
  xor2s1 U2629 ( .Q(n2266), .DIN1(n2267), .DIN2(n1955) );
  nnd2s1 U2630 ( .Q(n2267), .DIN1(n2247), .DIN2(n2268) );
  nnd3s1 U2631 ( .Q(n2268), .DIN1(n2269), .DIN2(n2270), .DIN3(n2271) );
  nnd2s1 U2632 ( .Q(n2271), .DIN1(g718), .DIN2(n2272) );
  nnd2s1 U2633 ( .Q(n2270), .DIN1(n2273), .DIN2(n2261) );
  nnd2s1 U2634 ( .Q(n2269), .DIN1(n2274), .DIN2(n2264) );
  nnd2s1 U2635 ( .Q(g9344), .DIN1(n2240), .DIN2(n2275) );
  nnd2s1 U2636 ( .Q(n2275), .DIN1(n2242), .DIN2(n2276) );
  xor2s1 U2637 ( .Q(n2276), .DIN1(n2277), .DIN2(n2029) );
  nnd2s1 U2638 ( .Q(n2277), .DIN1(n2247), .DIN2(n2278) );
  nnd3s1 U2639 ( .Q(n2278), .DIN1(n2279), .DIN2(n2280), .DIN3(n2281) );
  nnd2s1 U2640 ( .Q(n2281), .DIN1(g709), .DIN2(n2272) );
  nnd3s1 U2641 ( .Q(n2280), .DIN1(n2273), .DIN2(n1933), .DIN3(n1958) );
  nnd3s1 U2642 ( .Q(n2279), .DIN1(n2274), .DIN2(g686), .DIN3(g695) );
  nnd2s1 U2643 ( .Q(g9343), .DIN1(n2240), .DIN2(n2282) );
  nnd2s1 U2644 ( .Q(n2282), .DIN1(n2242), .DIN2(n2283) );
  xor2s1 U2645 ( .Q(n2283), .DIN1(n2284), .DIN2(n1958) );
  nnd2s1 U2646 ( .Q(n2284), .DIN1(n2247), .DIN2(n2285) );
  nnd3s1 U2647 ( .Q(n2285), .DIN1(n2286), .DIN2(n2287), .DIN3(n2288) );
  nnd2s1 U2648 ( .Q(n2288), .DIN1(g700), .DIN2(n2272) );
  nnd2s1 U2649 ( .Q(n2287), .DIN1(n2273), .DIN2(n1933) );
  hi1s1 U2650 ( .Q(n2273), .DIN(n2289) );
  nnd2s1 U2651 ( .Q(n2286), .DIN1(n2274), .DIN2(g686) );
  hi1s1 U2652 ( .Q(n2274), .DIN(n2290) );
  nnd2s1 U2653 ( .Q(g9342), .DIN1(n2240), .DIN2(n2291) );
  nnd2s1 U2654 ( .Q(n2291), .DIN1(n2242), .DIN2(n2292) );
  xor2s1 U2655 ( .Q(n2292), .DIN1(n2293), .DIN2(n1933) );
  nnd2s1 U2656 ( .Q(n2293), .DIN1(n2247), .DIN2(n2294) );
  nnd3s1 U2657 ( .Q(n2294), .DIN1(n2290), .DIN2(n2289), .DIN3(n2295) );
  nnd2s1 U2658 ( .Q(n2295), .DIN1(g691), .DIN2(n2272) );
  nnd2s1 U2659 ( .Q(n2289), .DIN1(n2248), .DIN2(n2260) );
  nnd2s1 U2660 ( .Q(n2290), .DIN1(n2248), .DIN2(n2263) );
  nnd2s1 U2661 ( .Q(g9341), .DIN1(n2240), .DIN2(n2296) );
  nnd2s1 U2662 ( .Q(n2296), .DIN1(n2242), .DIN2(n2297) );
  xor2s1 U2663 ( .Q(n2297), .DIN1(n2298), .DIN2(n1968) );
  nnd3s1 U2664 ( .Q(n2298), .DIN1(n2299), .DIN2(n2300), .DIN3(n2247) );
  or2s1 U2665 ( .Q(n2300), .DIN1(n2248), .DIN2(g682) );
  nnd2s1 U2666 ( .Q(n2299), .DIN1(n2248), .DIN2(n2301) );
  nnd3s1 U2667 ( .Q(n2301), .DIN1(n2302), .DIN2(n2303), .DIN3(n2304) );
  nnd2s1 U2668 ( .Q(n2304), .DIN1(g668), .DIN2(n2305) );
  nnd2s1 U2669 ( .Q(n2303), .DIN1(n2306), .DIN2(n2039) );
  nnd2s1 U2670 ( .Q(n2302), .DIN1(g658), .DIN2(n1936) );
  nnd2s1 U2671 ( .Q(g9340), .DIN1(n2240), .DIN2(n2307) );
  nnd2s1 U2672 ( .Q(n2307), .DIN1(n2242), .DIN2(n2308) );
  xor2s1 U2673 ( .Q(n2308), .DIN1(n2309), .DIN2(n1936) );
  nnd3s1 U2674 ( .Q(n2309), .DIN1(n2310), .DIN2(n2311), .DIN3(n2247) );
  hi1s1 U2675 ( .Q(n2247), .DIN(n2312) );
  or2s1 U2676 ( .Q(n2311), .DIN1(n2248), .DIN2(g673) );
  nnd2s1 U2677 ( .Q(n2310), .DIN1(n2313), .DIN2(n2248) );
  xor2s1 U2678 ( .Q(n2313), .DIN1(n2306), .DIN2(g658) );
  nnd2s1 U2679 ( .Q(g9339), .DIN1(n2240), .DIN2(n2314) );
  nnd2s1 U2680 ( .Q(n2314), .DIN1(n2242), .DIN2(n2315) );
  xor2s1 U2681 ( .Q(n2315), .DIN1(g658), .DIN2(n2316) );
  nor2s1 U2682 ( .Q(n2316), .DIN1(n2317), .DIN2(n2312) );
  nor2s1 U2683 ( .Q(n2312), .DIN1(n2272), .DIN2(n2318) );
  nor2s1 U2684 ( .Q(n2317), .DIN1(g664), .DIN2(n2248) );
  hi1s1 U2685 ( .Q(n2248), .DIN(n2272) );
  nnd2s1 U2686 ( .Q(n2272), .DIN1(n2319), .DIN2(n2320) );
  nnd2s1 U2687 ( .Q(n2320), .DIN1(g617), .DIN2(n2087) );
  nnd4s1 U2688 ( .Q(n2240), .DIN1(n2144), .DIN2(n2134), .DIN3(n2149), .DIN4(
        n2321) );
  nnd2s1 U2689 ( .Q(g9338), .DIN1(n2085), .DIN2(n2322) );
  nnd2s1 U2690 ( .Q(n2322), .DIN1(g622), .DIN2(n2323) );
  nnd2s1 U2691 ( .Q(n2323), .DIN1(n2321), .DIN2(n2324) );
  nnd2s1 U2692 ( .Q(n2324), .DIN1(n2134), .DIN2(n2149) );
  hi1s1 U2693 ( .Q(n2321), .DIN(n2242) );
  nor2s1 U2694 ( .Q(n2242), .DIN1(n2325), .DIN2(n2135) );
  nnd3s1 U2695 ( .Q(n2085), .DIN1(n2090), .DIN2(n1987), .DIN3(n2135) );
  hi1s1 U2696 ( .Q(n2135), .DIN(n2091) );
  nnd3s1 U2697 ( .Q(n2091), .DIN1(n2326), .DIN2(n2327), .DIN3(n2318) );
  and2s1 U2698 ( .Q(n2318), .DIN1(n2087), .DIN2(n2328) );
  nnd2s1 U2699 ( .Q(n2328), .DIN1(n2329), .DIN2(n2149) );
  or2s1 U2700 ( .Q(n2329), .DIN1(n1981), .DIN2(n2330) );
  nnd2s1 U2701 ( .Q(n2327), .DIN1(g731), .DIN2(n2250) );
  nnd4s1 U2702 ( .Q(n2250), .DIN1(g722), .DIN2(g713), .DIN3(n2263), .DIN4(
        n2264) );
  and3s1 U2703 ( .Q(n2264), .DIN1(g695), .DIN2(g686), .DIN3(g704) );
  and4s1 U2704 ( .Q(n2263), .DIN1(g677), .DIN2(g668), .DIN3(g658), .DIN4(n2306) );
  nnd2s1 U2705 ( .Q(n2326), .DIN1(n2249), .DIN2(n2009) );
  nnd4s1 U2706 ( .Q(n2249), .DIN1(n2260), .DIN2(n2261), .DIN3(n1955), .DIN4(
        n1994) );
  and3s1 U2707 ( .Q(n2261), .DIN1(n1958), .DIN2(n2029), .DIN3(n1933) );
  and4s1 U2708 ( .Q(n2260), .DIN1(n2305), .DIN2(n2039), .DIN3(n1936), .DIN4(
        n1968) );
  hi1s1 U2709 ( .Q(n2305), .DIN(n2306) );
  nnd2s1 U2710 ( .Q(n2306), .DIN1(n2139), .DIN2(g599) );
  and2s1 U2711 ( .Q(n2139), .DIN1(n2331), .DIN2(n2332) );
  nnd2s1 U2712 ( .Q(n2332), .DIN1(n2333), .DIN2(n1978) );
  hi1s1 U2713 ( .Q(n2090), .DIN(n2149) );
  nnd3s1 U2714 ( .Q(n2149), .DIN1(g591), .DIN2(n1982), .DIN3(g611) );
  and2s1 U2715 ( .Q(g8993), .DIN1(g109), .DIN2(n2334) );
  xor2s1 U2716 ( .Q(n2334), .DIN1(g1428), .DIN2(n2335) );
  and2s1 U2717 ( .Q(g8992), .DIN1(g109), .DIN2(n2336) );
  xor2s1 U2718 ( .Q(n2336), .DIN1(g1403), .DIN2(n2337) );
  and2s1 U2719 ( .Q(g8991), .DIN1(g109), .DIN2(n2338) );
  xor2s1 U2720 ( .Q(n2338), .DIN1(g1432), .DIN2(n2339) );
  and2s1 U2721 ( .Q(g8990), .DIN1(g109), .DIN2(n2340) );
  xor2s1 U2722 ( .Q(n2340), .DIN1(g1436), .DIN2(n2341) );
  and2s1 U2723 ( .Q(g8989), .DIN1(g109), .DIN2(n2342) );
  xor2s1 U2724 ( .Q(n2342), .DIN1(g1440), .DIN2(n2343) );
  and2s1 U2725 ( .Q(g8988), .DIN1(g109), .DIN2(n2344) );
  xor2s1 U2726 ( .Q(n2344), .DIN1(g1444), .DIN2(n2345) );
  and2s1 U2727 ( .Q(g8987), .DIN1(g109), .DIN2(n2346) );
  xor2s1 U2728 ( .Q(n2346), .DIN1(g1448), .DIN2(n2347) );
  nnd2s1 U2729 ( .Q(g8874), .DIN1(n2348), .DIN2(n2349) );
  nnd2s1 U2730 ( .Q(n2349), .DIN1(g1636), .DIN2(n2070) );
  nnd2s1 U2731 ( .Q(n2348), .DIN1(n2063), .DIN2(n2347) );
  nnd2s1 U2732 ( .Q(n2347), .DIN1(n2351), .DIN2(n2352) );
  nnd2s1 U2733 ( .Q(n2352), .DIN1(n2353), .DIN2(n2072) );
  xor2s1 U2734 ( .Q(n2353), .DIN1(g1145), .DIN2(n2354) );
  nor2s1 U2735 ( .Q(n2354), .DIN1(n1974), .DIN2(n2355) );
  nnd2s1 U2736 ( .Q(g8873), .DIN1(n2356), .DIN2(n2357) );
  nnd2s1 U2737 ( .Q(n2357), .DIN1(g1633), .DIN2(n2068) );
  nnd2s1 U2738 ( .Q(n2356), .DIN1(n2063), .DIN2(n2345) );
  nnd2s1 U2739 ( .Q(n2345), .DIN1(n2358), .DIN2(n2359) );
  nnd2s1 U2740 ( .Q(n2359), .DIN1(n2360), .DIN2(n2082) );
  xor2s1 U2741 ( .Q(n2360), .DIN1(g1141), .DIN2(n2361) );
  nor2s1 U2742 ( .Q(n2361), .DIN1(g1101), .DIN2(n2355) );
  nnd3s1 U2743 ( .Q(n2355), .DIN1(n1976), .DIN2(n1929), .DIN3(g1110) );
  nnd2s1 U2744 ( .Q(g8872), .DIN1(n2362), .DIN2(n2363) );
  nnd2s1 U2745 ( .Q(n2363), .DIN1(g1630), .DIN2(n2069) );
  nnd2s1 U2746 ( .Q(n2362), .DIN1(n2350), .DIN2(n2343) );
  nnd2s1 U2747 ( .Q(n2343), .DIN1(n2364), .DIN2(n2365) );
  nnd2s1 U2748 ( .Q(n2365), .DIN1(n2366), .DIN2(n2082) );
  xor2s1 U2749 ( .Q(n2366), .DIN1(g1137), .DIN2(n2367) );
  nor2s1 U2750 ( .Q(n2367), .DIN1(n1974), .DIN2(n2368) );
  nnd2s1 U2751 ( .Q(g8871), .DIN1(n2369), .DIN2(n2370) );
  nnd2s1 U2752 ( .Q(n2370), .DIN1(g1627), .DIN2(n2070) );
  nnd2s1 U2753 ( .Q(n2369), .DIN1(n2063), .DIN2(n2341) );
  nnd2s1 U2754 ( .Q(n2341), .DIN1(n2371), .DIN2(n2372) );
  nnd2s1 U2755 ( .Q(n2372), .DIN1(n2373), .DIN2(n2082) );
  xor2s1 U2756 ( .Q(n2373), .DIN1(g1133), .DIN2(n2374) );
  nor2s1 U2757 ( .Q(n2374), .DIN1(g1101), .DIN2(n2368) );
  nnd3s1 U2758 ( .Q(n2368), .DIN1(g1104), .DIN2(n1949), .DIN3(g1107) );
  nnd2s1 U2759 ( .Q(g8870), .DIN1(n2375), .DIN2(n2376) );
  nnd2s1 U2760 ( .Q(n2376), .DIN1(g1624), .DIN2(n2068) );
  nnd2s1 U2761 ( .Q(n2375), .DIN1(n2063), .DIN2(n2339) );
  nnd2s1 U2762 ( .Q(n2339), .DIN1(n2377), .DIN2(n2378) );
  nnd2s1 U2763 ( .Q(n2378), .DIN1(n2379), .DIN2(n2072) );
  xor2s1 U2764 ( .Q(n2379), .DIN1(g1129), .DIN2(n2380) );
  nor2s1 U2765 ( .Q(n2380), .DIN1(n1974), .DIN2(n2381) );
  nnd2s1 U2766 ( .Q(g8869), .DIN1(n2382), .DIN2(n2383) );
  nnd2s1 U2767 ( .Q(n2383), .DIN1(g1621), .DIN2(n2069) );
  nnd2s1 U2768 ( .Q(n2382), .DIN1(n2350), .DIN2(n2337) );
  nnd2s1 U2769 ( .Q(n2337), .DIN1(n2384), .DIN2(n2385) );
  nnd2s1 U2770 ( .Q(n2385), .DIN1(n2386), .DIN2(n2082) );
  xor2s1 U2771 ( .Q(n2386), .DIN1(g1125), .DIN2(n2387) );
  nor2s1 U2772 ( .Q(n2387), .DIN1(g1101), .DIN2(n2381) );
  nnd3s1 U2773 ( .Q(n2381), .DIN1(n1976), .DIN2(n1949), .DIN3(g1107) );
  nnd2s1 U2774 ( .Q(g8868), .DIN1(n2388), .DIN2(n2389) );
  nnd2s1 U2775 ( .Q(n2389), .DIN1(g1615), .DIN2(n2070) );
  nnd2s1 U2776 ( .Q(n2388), .DIN1(n2350), .DIN2(n2335) );
  nnd2s1 U2777 ( .Q(n2335), .DIN1(n2390), .DIN2(n2391) );
  nnd2s1 U2778 ( .Q(n2391), .DIN1(n2392), .DIN2(n2072) );
  xor2s1 U2779 ( .Q(n2392), .DIN1(g1121), .DIN2(n2393) );
  nor2s1 U2780 ( .Q(n2393), .DIN1(n2394), .DIN2(n1974) );
  nnd3s1 U2781 ( .Q(g8782), .DIN1(n2395), .DIN2(n2396), .DIN3(n2134) );
  nnd2s1 U2782 ( .Q(n2396), .DIN1(g664), .DIN2(n2397) );
  nnd2s1 U2783 ( .Q(g8781), .DIN1(n2398), .DIN2(n2399) );
  nnd2s1 U2784 ( .Q(n2399), .DIN1(n2325), .DIN2(n2400) );
  nnd3s1 U2785 ( .Q(n2400), .DIN1(n2401), .DIN2(n2402), .DIN3(g4190) );
  nnd2s1 U2786 ( .Q(n2402), .DIN1(n2403), .DIN2(n2404) );
  nnd2s1 U2787 ( .Q(n2404), .DIN1(g4187), .DIN2(g4186) );
  nnd2s1 U2788 ( .Q(n2403), .DIN1(g4189), .DIN2(g4188) );
  nnd2s1 U2789 ( .Q(n2401), .DIN1(n2405), .DIN2(n2406) );
  nnd2s1 U2790 ( .Q(n2405), .DIN1(g4185), .DIN2(g4184) );
  nnd2s1 U2791 ( .Q(n2398), .DIN1(n2407), .DIN2(n2134) );
  nnd2s1 U2792 ( .Q(n2407), .DIN1(n2408), .DIN2(n2409) );
  nnd2s1 U2793 ( .Q(n2409), .DIN1(g2613), .DIN2(n2410) );
  nnd3s1 U2794 ( .Q(n2410), .DIN1(n2411), .DIN2(n2412), .DIN3(g5656) );
  nnd3s1 U2795 ( .Q(n2412), .DIN1(n2150), .DIN2(n1975), .DIN3(n2413) );
  nnd2s1 U2796 ( .Q(n2413), .DIN1(n2414), .DIN2(g591) );
  nnd2s1 U2797 ( .Q(n2414), .DIN1(g617), .DIN2(n2330) );
  xor2s1 U2798 ( .Q(n2411), .DIN1(n2415), .DIN2(n2416) );
  nnd2s1 U2799 ( .Q(n2416), .DIN1(n2417), .DIN2(n2418) );
  nnd2s1 U2800 ( .Q(n2418), .DIN1(n2333), .DIN2(g639) );
  nnd2s1 U2801 ( .Q(n2417), .DIN1(n2419), .DIN2(n1981) );
  nnd2s1 U2802 ( .Q(n2419), .DIN1(n1975), .DIN2(n2420) );
  nor2s1 U2803 ( .Q(n2415), .DIN1(n1987), .DIN2(\DFF_270/net557 ) );
  or2s1 U2804 ( .Q(n2408), .DIN1(n2331), .DIN2(g622) );
  nor2s1 U2805 ( .Q(g8780), .DIN1(n2072), .DIN2(n2421) );
  xor2s1 U2806 ( .Q(n2421), .DIN1(n2422), .DIN2(n1982) );
  nnd2s1 U2807 ( .Q(n2422), .DIN1(n2395), .DIN2(n2423) );
  or2s1 U2808 ( .Q(n2423), .DIN1(n2319), .DIN2(g617) );
  nnd4s1 U2809 ( .Q(n2319), .DIN1(n2330), .DIN2(n2087), .DIN3(g591), .DIN4(
        n1975) );
  nnd2s1 U2810 ( .Q(n2395), .DIN1(g736), .DIN2(n2424) );
  nnd3s1 U2811 ( .Q(g8695), .DIN1(n2425), .DIN2(n2426), .DIN3(n2102) );
  nnd2s1 U2812 ( .Q(n2426), .DIN1(g1878), .DIN2(n2427) );
  nor2s1 U2813 ( .Q(g8694), .DIN1(n2082), .DIN2(n2428) );
  xor2s1 U2814 ( .Q(n2428), .DIN1(n2429), .DIN2(n1983) );
  nnd2s1 U2815 ( .Q(n2429), .DIN1(n2425), .DIN2(n2430) );
  or2s1 U2816 ( .Q(n2430), .DIN1(n2230), .DIN2(g1840) );
  nnd4s1 U2817 ( .Q(n2230), .DIN1(n2238), .DIN2(n2095), .DIN3(g1814), .DIN4(
        n1948) );
  nnd2s1 U2818 ( .Q(n2425), .DIN1(g1950), .DIN2(n2431) );
  nor2s1 U2819 ( .Q(g8573), .DIN1(g5653), .DIN2(n2432) );
  xor2s1 U2820 ( .Q(n2432), .DIN1(g1806), .DIN2(n2433) );
  nnd2s1 U2821 ( .Q(n2433), .DIN1(g1801), .DIN2(n2434) );
  nor2s1 U2822 ( .Q(g8572), .DIN1(n2435), .DIN2(n2045) );
  nor2s1 U2823 ( .Q(g8571), .DIN1(n2435), .DIN2(n2046) );
  nor2s1 U2824 ( .Q(g8570), .DIN1(n2435), .DIN2(n2007) );
  nor2s1 U2825 ( .Q(g8569), .DIN1(n2435), .DIN2(n2047) );
  nnd2s1 U2826 ( .Q(n2435), .DIN1(g109), .DIN2(n2436) );
  nnd3s1 U2827 ( .Q(n2436), .DIN1(\DFF_436/net723 ), .DIN2(n2437), .DIN3(n2438) );
  and2s1 U2828 ( .Q(g8568), .DIN1(n2439), .DIN2(n2440) );
  xor2s1 U2829 ( .Q(n2439), .DIN1(n2441), .DIN2(g4190) );
  nor2s1 U2830 ( .Q(n2441), .DIN1(n2043), .DIN2(n2442) );
  and3s1 U2831 ( .Q(g8567), .DIN1(n2443), .DIN2(n2444), .DIN3(n2445) );
  nnd2s1 U2832 ( .Q(n2443), .DIN1(n2055), .DIN2(n2446) );
  nnd2s1 U2833 ( .Q(n2446), .DIN1(g786), .DIN2(n2447) );
  nor2s1 U2834 ( .Q(g8450), .DIN1(g5653), .DIN2(n2448) );
  xor2s1 U2835 ( .Q(n2448), .DIN1(g1801), .DIN2(n2449) );
  nnd2s1 U2836 ( .Q(g8449), .DIN1(n2450), .DIN2(n2451) );
  nnd2s1 U2837 ( .Q(n2451), .DIN1(g1512), .DIN2(n2068) );
  nnd2s1 U2838 ( .Q(n2450), .DIN1(n2452), .DIN2(n2063) );
  xor2s1 U2839 ( .Q(n2452), .DIN1(n2453), .DIN2(n1934) );
  nnd4s1 U2840 ( .Q(n2453), .DIN1(g1110), .DIN2(g1104), .DIN3(n1974), .DIN4(
        n1929) );
  nnd2s1 U2841 ( .Q(g8448), .DIN1(n2454), .DIN2(n2455) );
  nnd2s1 U2842 ( .Q(n2455), .DIN1(g1639), .DIN2(n2069) );
  nnd2s1 U2843 ( .Q(n2454), .DIN1(n2456), .DIN2(n2063) );
  xor2s1 U2844 ( .Q(n2456), .DIN1(g1117), .DIN2(n2457) );
  nor2s1 U2845 ( .Q(n2457), .DIN1(g1101), .DIN2(n2394) );
  nnd3s1 U2846 ( .Q(n2394), .DIN1(n1929), .DIN2(n1949), .DIN3(g1104) );
  and2s1 U2847 ( .Q(g8447), .DIN1(g109), .DIN2(n2458) );
  xor2s1 U2848 ( .Q(n2458), .DIN1(g1494), .DIN2(n2459) );
  nor2s1 U2849 ( .Q(g8446), .DIN1(n2064), .DIN2(n2460) );
  xor2s1 U2850 ( .Q(n2460), .DIN1(g1490), .DIN2(n2461) );
  nor2s1 U2851 ( .Q(g8445), .DIN1(n2066), .DIN2(n2462) );
  xor2s1 U2852 ( .Q(n2462), .DIN1(g1486), .DIN2(n2463) );
  nor2s1 U2853 ( .Q(g8444), .DIN1(n2064), .DIN2(n2464) );
  xor2s1 U2854 ( .Q(n2464), .DIN1(g1482), .DIN2(n2465) );
  and2s1 U2855 ( .Q(g8443), .DIN1(g109), .DIN2(n2466) );
  xor2s1 U2856 ( .Q(n2466), .DIN1(g1478), .DIN2(n2467) );
  and2s1 U2857 ( .Q(g8442), .DIN1(g109), .DIN2(n2468) );
  xor2s1 U2858 ( .Q(n2468), .DIN1(g1474), .DIN2(n2469) );
  and2s1 U2859 ( .Q(g8441), .DIN1(g109), .DIN2(n2470) );
  xor2s1 U2860 ( .Q(n2470), .DIN1(g1470), .DIN2(n2471) );
  and2s1 U2861 ( .Q(g8440), .DIN1(n2472), .DIN2(g109) );
  xor2s1 U2862 ( .Q(n2472), .DIN1(g1466), .DIN2(n2473) );
  and2s1 U2863 ( .Q(g8439), .DIN1(n2474), .DIN2(g109) );
  xor2s1 U2864 ( .Q(n2474), .DIN1(g1462), .DIN2(n2475) );
  nor2s1 U2865 ( .Q(g8438), .DIN1(n2476), .DIN2(n2065) );
  xor2s1 U2866 ( .Q(n2476), .DIN1(n1991), .DIN2(n2477) );
  nor2s1 U2867 ( .Q(g8437), .DIN1(n2478), .DIN2(n2479) );
  xor2s1 U2868 ( .Q(n2478), .DIN1(g4189), .DIN2(n2442) );
  nor2s1 U2869 ( .Q(g8436), .DIN1(n2480), .DIN2(n2481) );
  xor2s1 U2870 ( .Q(n2480), .DIN1(g786), .DIN2(n2482) );
  nnd2s1 U2871 ( .Q(g8435), .DIN1(n2483), .DIN2(n2484) );
  nnd2s1 U2872 ( .Q(n2484), .DIN1(n2485), .DIN2(g736) );
  nnd2s1 U2873 ( .Q(n2483), .DIN1(g727), .DIN2(n2424) );
  nnd2s1 U2874 ( .Q(g8434), .DIN1(n2486), .DIN2(n2487) );
  nnd2s1 U2875 ( .Q(n2487), .DIN1(g727), .DIN2(n2485) );
  nnd2s1 U2876 ( .Q(n2486), .DIN1(n2424), .DIN2(g718) );
  nnd2s1 U2877 ( .Q(g8433), .DIN1(n2488), .DIN2(n2489) );
  nnd2s1 U2878 ( .Q(n2489), .DIN1(n2485), .DIN2(g718) );
  nnd2s1 U2879 ( .Q(n2488), .DIN1(n2424), .DIN2(g709) );
  nnd2s1 U2880 ( .Q(g8432), .DIN1(n2490), .DIN2(n2491) );
  nnd2s1 U2881 ( .Q(n2491), .DIN1(n2485), .DIN2(g709) );
  nnd2s1 U2882 ( .Q(n2490), .DIN1(n2424), .DIN2(g700) );
  nnd2s1 U2883 ( .Q(g8431), .DIN1(n2492), .DIN2(n2493) );
  nnd2s1 U2884 ( .Q(n2493), .DIN1(n2485), .DIN2(g700) );
  nnd2s1 U2885 ( .Q(n2492), .DIN1(n2424), .DIN2(g691) );
  nnd2s1 U2886 ( .Q(g8430), .DIN1(n2494), .DIN2(n2495) );
  nnd2s1 U2887 ( .Q(n2495), .DIN1(n2485), .DIN2(g691) );
  nnd2s1 U2888 ( .Q(n2494), .DIN1(g682), .DIN2(n2424) );
  nnd2s1 U2889 ( .Q(g8429), .DIN1(n2496), .DIN2(n2497) );
  nnd2s1 U2890 ( .Q(n2497), .DIN1(g682), .DIN2(n2485) );
  nnd2s1 U2891 ( .Q(n2496), .DIN1(g673), .DIN2(n2424) );
  nnd2s1 U2892 ( .Q(g8428), .DIN1(n2498), .DIN2(n2499) );
  nnd2s1 U2893 ( .Q(n2499), .DIN1(g673), .DIN2(n2485) );
  nor2s1 U2894 ( .Q(n2485), .DIN1(n2424), .DIN2(n2325) );
  nnd2s1 U2895 ( .Q(n2498), .DIN1(g664), .DIN2(n2424) );
  hi1s1 U2896 ( .Q(n2424), .DIN(n2397) );
  nnd3s1 U2897 ( .Q(n2397), .DIN1(n2087), .DIN2(n1975), .DIN3(g617) );
  nor2s1 U2898 ( .Q(g8427), .DIN1(n2067), .DIN2(n2500) );
  xor2s1 U2899 ( .Q(n2500), .DIN1(n1937), .DIN2(g7750) );
  nor2s1 U2900 ( .Q(g8426), .DIN1(n2067), .DIN2(n2501) );
  xor2s1 U2901 ( .Q(n2501), .DIN1(n1992), .DIN2(g7752) );
  nor2s1 U2902 ( .Q(g8425), .DIN1(n2066), .DIN2(n2502) );
  xor2s1 U2903 ( .Q(n2502), .DIN1(n1959), .DIN2(g7753) );
  and2s1 U2904 ( .Q(g8424), .DIN1(g109), .DIN2(n2503) );
  xor2s1 U2905 ( .Q(n2503), .DIN1(g174), .DIN2(g7754) );
  and2s1 U2906 ( .Q(g8423), .DIN1(g109), .DIN2(n2504) );
  xor2s1 U2907 ( .Q(n2504), .DIN1(g170), .DIN2(g7755) );
  nor2s1 U2908 ( .Q(g8422), .DIN1(n2066), .DIN2(n2505) );
  xor2s1 U2909 ( .Q(n2505), .DIN1(n1960), .DIN2(g7756) );
  nor2s1 U2910 ( .Q(g8421), .DIN1(n2067), .DIN2(n2506) );
  xor2s1 U2911 ( .Q(n2506), .DIN1(n1996), .DIN2(g7757) );
  nor2s1 U2912 ( .Q(g8420), .DIN1(n2507), .DIN2(n2065) );
  xor2s1 U2913 ( .Q(n2507), .DIN1(n1961), .DIN2(g7758) );
  nor2s1 U2914 ( .Q(g8419), .DIN1(n2508), .DIN2(n2065) );
  xor2s1 U2915 ( .Q(n2508), .DIN1(n1938), .DIN2(g7759) );
  and2s1 U2916 ( .Q(g8418), .DIN1(n2509), .DIN2(g109) );
  xor2s1 U2917 ( .Q(n2509), .DIN1(g166), .DIN2(g7751) );
  nnd2s1 U2918 ( .Q(g8288), .DIN1(n2510), .DIN2(n2511) );
  nnd2s1 U2919 ( .Q(n2511), .DIN1(n2512), .DIN2(g1950) );
  nnd2s1 U2920 ( .Q(n2510), .DIN1(g1941), .DIN2(n2431) );
  nnd2s1 U2921 ( .Q(g8287), .DIN1(n2513), .DIN2(n2514) );
  nnd2s1 U2922 ( .Q(n2514), .DIN1(g1941), .DIN2(n2512) );
  nnd2s1 U2923 ( .Q(n2513), .DIN1(n2431), .DIN2(g1932) );
  nnd2s1 U2924 ( .Q(g8286), .DIN1(n2515), .DIN2(n2516) );
  nnd2s1 U2925 ( .Q(n2516), .DIN1(n2512), .DIN2(g1932) );
  nnd2s1 U2926 ( .Q(n2515), .DIN1(n2431), .DIN2(g1923) );
  nnd2s1 U2927 ( .Q(g8285), .DIN1(n2517), .DIN2(n2518) );
  nnd2s1 U2928 ( .Q(n2518), .DIN1(n2512), .DIN2(g1923) );
  nnd2s1 U2929 ( .Q(n2517), .DIN1(n2431), .DIN2(g1914) );
  nnd2s1 U2930 ( .Q(g8284), .DIN1(n2519), .DIN2(n2520) );
  nnd2s1 U2931 ( .Q(n2520), .DIN1(n2512), .DIN2(g1914) );
  nnd2s1 U2932 ( .Q(n2519), .DIN1(n2431), .DIN2(g1905) );
  nnd2s1 U2933 ( .Q(g8283), .DIN1(n2521), .DIN2(n2522) );
  nnd2s1 U2934 ( .Q(n2522), .DIN1(n2512), .DIN2(g1905) );
  nnd2s1 U2935 ( .Q(n2521), .DIN1(g1896), .DIN2(n2431) );
  nnd2s1 U2936 ( .Q(g8282), .DIN1(n2523), .DIN2(n2524) );
  nnd2s1 U2937 ( .Q(n2524), .DIN1(g1896), .DIN2(n2512) );
  nnd2s1 U2938 ( .Q(n2523), .DIN1(g1887), .DIN2(n2431) );
  nnd2s1 U2939 ( .Q(g8281), .DIN1(n2525), .DIN2(n2526) );
  nnd2s1 U2940 ( .Q(n2526), .DIN1(g1887), .DIN2(n2512) );
  nor2s1 U2941 ( .Q(n2512), .DIN1(n2431), .DIN2(n2233) );
  nnd2s1 U2942 ( .Q(n2525), .DIN1(g1878), .DIN2(n2431) );
  hi1s1 U2943 ( .Q(n2431), .DIN(n2427) );
  nnd3s1 U2944 ( .Q(n2427), .DIN1(g1840), .DIN2(n1948), .DIN3(n2095) );
  and3s1 U2945 ( .Q(g8280), .DIN1(n2449), .DIN2(n2061), .DIN3(n2527) );
  nnd2s1 U2946 ( .Q(n2527), .DIN1(n2528), .DIN2(n1952) );
  hi1s1 U2947 ( .Q(n2449), .DIN(n2434) );
  nor2s1 U2948 ( .Q(n2434), .DIN1(n1952), .DIN2(n2528) );
  nor2s1 U2949 ( .Q(g8279), .DIN1(n2529), .DIN2(n2530) );
  nor2s1 U2950 ( .Q(n2529), .DIN1(n2531), .DIN2(g1231) );
  nor2s1 U2951 ( .Q(g8278), .DIN1(n2532), .DIN2(n2530) );
  and2s1 U2952 ( .Q(n2532), .DIN1(n2533), .DIN2(n2534) );
  nnd3s1 U2953 ( .Q(n2534), .DIN1(g1223), .DIN2(n2535), .DIN3(n2536) );
  hi1s1 U2954 ( .Q(n2536), .DIN(n2537) );
  nnd2s1 U2955 ( .Q(n2533), .DIN1(g1227), .DIN2(n2538) );
  hi1s1 U2956 ( .Q(n2538), .DIN(n2531) );
  nor2s1 U2957 ( .Q(n2531), .DIN1(n2539), .DIN2(n2535) );
  nor2s1 U2958 ( .Q(g8277), .DIN1(n2540), .DIN2(n2530) );
  xor2s1 U2959 ( .Q(n2540), .DIN1(g1223), .DIN2(n2537) );
  nnd2s1 U2960 ( .Q(n2537), .DIN1(n2541), .DIN2(g1218) );
  nor2s1 U2961 ( .Q(g8276), .DIN1(n2542), .DIN2(n2530) );
  or2s1 U2962 ( .Q(n2530), .DIN1(n2067), .DIN2(g1212) );
  xor2s1 U2963 ( .Q(n2542), .DIN1(g1218), .DIN2(n2539) );
  hi1s1 U2964 ( .Q(n2539), .DIN(n2541) );
  nor2s1 U2965 ( .Q(n2541), .DIN1(n2543), .DIN2(n2544) );
  hi1s1 U2966 ( .Q(g8275), .DIN(n2545) );
  xor2s1 U2967 ( .Q(n2545), .DIN1(n2444), .DIN2(g590) );
  nnd3s1 U2968 ( .Q(n2444), .DIN1(g786), .DIN2(n2447), .DIN3(g790) );
  hi1s1 U2969 ( .Q(n2447), .DIN(n2482) );
  and3s1 U2970 ( .Q(g8274), .DIN1(n2546), .DIN2(n2442), .DIN3(n2440) );
  nnd3s1 U2971 ( .Q(n2442), .DIN1(g4188), .DIN2(g4187), .DIN3(n2547) );
  nnd2s1 U2972 ( .Q(n2546), .DIN1(n2049), .DIN2(n2548) );
  nnd2s1 U2973 ( .Q(n2548), .DIN1(n2547), .DIN2(g4187) );
  hi1s1 U2974 ( .Q(n2547), .DIN(n2549) );
  and3s1 U2975 ( .Q(g8273), .DIN1(n2550), .DIN2(n2482), .DIN3(n2445) );
  nnd3s1 U2976 ( .Q(n2482), .DIN1(g778), .DIN2(n2551), .DIN3(g782) );
  nnd2s1 U2977 ( .Q(n2550), .DIN1(n2056), .DIN2(n2552) );
  nnd2s1 U2978 ( .Q(n2552), .DIN1(g778), .DIN2(n2551) );
  hi1s1 U2979 ( .Q(n2551), .DIN(n2553) );
  nnd2s1 U2980 ( .Q(g8272), .DIN1(n2554), .DIN2(n2555) );
  or4s1 U2981 ( .Q(n2555), .DIN1(n2556), .DIN2(n2557), .DIN3(n2558), .DIN4(
        n2559) );
  nnd4s1 U2982 ( .Q(n2559), .DIN1(n1996), .DIN2(n1961), .DIN3(n1938), .DIN4(
        n1925) );
  nnd4s1 U2983 ( .Q(n2558), .DIN1(n1926), .DIN2(n1937), .DIN3(n1992), .DIN4(
        n1959) );
  nnd4s1 U2984 ( .Q(n2557), .DIN1(g182), .DIN2(g7749), .DIN3(n2560), .DIN4(
        g166) );
  nnd4s1 U2985 ( .Q(n2556), .DIN1(g170), .DIN2(g174), .DIN3(n2017), .DIN4(
        n1960) );
  nnd2s1 U2986 ( .Q(n2554), .DIN1(g123), .DIN2(g109) );
  nnd2s1 U2987 ( .Q(g8241), .DIN1(n2023), .DIN2(n2561) );
  nnd2s1 U2988 ( .Q(g8236), .DIN1(n2034), .DIN2(n2561) );
  nnd2s1 U2989 ( .Q(g8230), .DIN1(n2018), .DIN2(n2561) );
  nnd2s1 U2990 ( .Q(g8226), .DIN1(n2035), .DIN2(n2561) );
  nnd2s1 U2991 ( .Q(g8221), .DIN1(n2019), .DIN2(n2561) );
  nnd2s1 U2992 ( .Q(g8214), .DIN1(n2036), .DIN2(n2561) );
  nnd2s1 U2993 ( .Q(g8210), .DIN1(n2020), .DIN2(n2561) );
  nnd2s1 U2994 ( .Q(g8206), .DIN1(n2037), .DIN2(n2561) );
  nnd2s1 U2995 ( .Q(g8203), .DIN1(n2021), .DIN2(n2561) );
  nnd2s1 U2996 ( .Q(g8200), .DIN1(n2038), .DIN2(n2561) );
  nnd2s1 U2997 ( .Q(g8187), .DIN1(n2022), .DIN2(n2561) );
  hi1s1 U2998 ( .Q(n2561), .DIN(g82) );
  nor2s1 U2999 ( .Q(g8080), .DIN1(g5653), .DIN2(n2562) );
  and2s1 U3000 ( .Q(n2562), .DIN1(n2563), .DIN2(n2564) );
  nnd3s1 U3001 ( .Q(n2564), .DIN1(g1786), .DIN2(n2565), .DIN3(n2566) );
  nnd2s1 U3002 ( .Q(n2563), .DIN1(g1791), .DIN2(n2528) );
  or2s1 U3003 ( .Q(n2528), .DIN1(n2567), .DIN2(n2565) );
  nnd4s1 U3004 ( .Q(n2565), .DIN1(g1791), .DIN2(g1786), .DIN3(g1781), .DIN4(
        n2568) );
  nnd2s1 U3005 ( .Q(g8079), .DIN1(n2569), .DIN2(n2570) );
  or3s1 U3006 ( .Q(n2570), .DIN1(n2571), .DIN2(n2572), .DIN3(n2573) );
  nnd4s1 U3007 ( .Q(n2573), .DIN1(g1453), .DIN2(g7329), .DIN3(g1508), .DIN4(
        n2574) );
  and4s1 U3008 ( .Q(n2574), .DIN1(n2575), .DIN2(g1462), .DIN3(g1470), .DIN4(
        g1474) );
  nnd4s1 U3009 ( .Q(n2572), .DIN1(g1478), .DIN2(g1490), .DIN3(g1494), .DIN4(
        n1991) );
  or4s1 U3010 ( .Q(n2571), .DIN1(g1466), .DIN2(g1482), .DIN3(g1486), .DIN4(
        g1499) );
  nnd2s1 U3011 ( .Q(n2569), .DIN1(g4), .DIN2(g109) );
  nnd2s1 U3012 ( .Q(g8078), .DIN1(n2576), .DIN2(n2577) );
  or4s1 U3013 ( .Q(n2577), .DIN1(n2578), .DIN2(n2579), .DIN3(n2580), .DIN4(
        n2581) );
  nnd4s1 U3014 ( .Q(n2581), .DIN1(g1440), .DIN2(g1436), .DIN3(g1432), .DIN4(
        g1428) );
  or4s1 U3015 ( .Q(n2580), .DIN1(g1403), .DIN2(g1407), .DIN3(g1411), .DIN4(
        g1415) );
  nnd3s1 U3016 ( .Q(n2579), .DIN1(g1424), .DIN2(g1419), .DIN3(g1515) );
  nnd4s1 U3017 ( .Q(n2578), .DIN1(g7335), .DIN2(n2575), .DIN3(g1448), .DIN4(
        g1444) );
  nnd2s1 U3018 ( .Q(n2576), .DIN1(g1), .DIN2(g109) );
  nor2s1 U3019 ( .Q(g8077), .DIN1(n2582), .DIN2(n2479) );
  xor2s1 U3020 ( .Q(n2582), .DIN1(g4187), .DIN2(n2549) );
  nor2s1 U3021 ( .Q(g8076), .DIN1(n2583), .DIN2(n2481) );
  xor2s1 U3022 ( .Q(n2583), .DIN1(g778), .DIN2(n2553) );
  nnd2s1 U3023 ( .Q(g8067), .DIN1(n2584), .DIN2(n2585) );
  nnd2s1 U3024 ( .Q(n2585), .DIN1(g654), .DIN2(n2586) );
  nor2s1 U3025 ( .Q(g8066), .DIN1(n2587), .DIN2(n2588) );
  nor2s1 U3026 ( .Q(n2587), .DIN1(n2589), .DIN2(n2590) );
  hi1s1 U3027 ( .Q(n2590), .DIN(n2586) );
  nor2s1 U3028 ( .Q(n2589), .DIN1(n2591), .DIN2(n2026) );
  nor2s1 U3029 ( .Q(g8065), .DIN1(n2592), .DIN2(n2588) );
  hi1s1 U3030 ( .Q(n2588), .DIN(n2584) );
  nor2s1 U3031 ( .Q(n2592), .DIN1(n2593), .DIN2(n2591) );
  and2s1 U3032 ( .Q(n2593), .DIN1(n2594), .DIN2(g646) );
  nnd3s1 U3033 ( .Q(g8064), .DIN1(n2595), .DIN2(n2594), .DIN3(n2584) );
  nor2s1 U3034 ( .Q(n2584), .DIN1(n2325), .DIN2(n2087) );
  hi1s1 U3035 ( .Q(n2325), .DIN(n2134) );
  nnd2s1 U3036 ( .Q(n2595), .DIN1(g643), .DIN2(n1997) );
  nnd3s1 U3037 ( .Q(g8063), .DIN1(n2596), .DIN2(n2597), .DIN3(n2134) );
  nnd3s1 U3038 ( .Q(n2597), .DIN1(n2087), .DIN2(n2598), .DIN3(n1981) );
  nnd3s1 U3039 ( .Q(n2598), .DIN1(n2150), .DIN2(n2420), .DIN3(n2144) );
  and2s1 U3040 ( .Q(n2144), .DIN1(n2331), .DIN2(n2599) );
  nnd2s1 U3041 ( .Q(n2599), .DIN1(g599), .DIN2(n1978) );
  nnd3s1 U3042 ( .Q(n2331), .DIN1(n1951), .DIN2(n1985), .DIN3(g605) );
  hi1s1 U3043 ( .Q(n2420), .DIN(n2140) );
  nor2s1 U3044 ( .Q(n2140), .DIN1(n1978), .DIN2(n1951) );
  hi1s1 U3045 ( .Q(n2150), .DIN(n2333) );
  nor2s1 U3046 ( .Q(n2333), .DIN1(n1985), .DIN2(g591) );
  or2s1 U3047 ( .Q(n2596), .DIN1(n1981), .DIN2(n2087) );
  nor2s1 U3048 ( .Q(n2087), .DIN1(n2586), .DIN2(g654) );
  nnd2s1 U3049 ( .Q(n2586), .DIN1(n2591), .DIN2(n2026) );
  nor2s1 U3050 ( .Q(n2591), .DIN1(n2594), .DIN2(g646) );
  or2s1 U3051 ( .Q(n2594), .DIN1(n1997), .DIN2(g643) );
  nnd2s1 U3052 ( .Q(g7817), .DIN1(n2600), .DIN2(n2601) );
  nnd2s1 U3053 ( .Q(n2601), .DIN1(g1868), .DIN2(n2602) );
  nor2s1 U3054 ( .Q(g7816), .DIN1(n2603), .DIN2(n2604) );
  nor2s1 U3055 ( .Q(n2603), .DIN1(n2605), .DIN2(n2606) );
  hi1s1 U3056 ( .Q(n2606), .DIN(n2602) );
  nor2s1 U3057 ( .Q(n2605), .DIN1(n2607), .DIN2(n2027) );
  nor2s1 U3058 ( .Q(g7815), .DIN1(n2608), .DIN2(n2604) );
  hi1s1 U3059 ( .Q(n2604), .DIN(n2600) );
  nor2s1 U3060 ( .Q(n2608), .DIN1(n2609), .DIN2(n2607) );
  and2s1 U3061 ( .Q(n2609), .DIN1(n1998), .DIN2(g1861) );
  nor2s1 U3062 ( .Q(g7814), .DIN1(g5653), .DIN2(n2610) );
  xor2s1 U3063 ( .Q(n2610), .DIN1(g1786), .DIN2(n2611) );
  and3s1 U3064 ( .Q(g7813), .DIN1(n2611), .DIN2(n2061), .DIN3(n2612) );
  nnd2s1 U3065 ( .Q(n2612), .DIN1(n2613), .DIN2(n1984) );
  hi1s1 U3066 ( .Q(n2611), .DIN(n2566) );
  nor2s1 U3067 ( .Q(n2566), .DIN1(n2613), .DIN2(n1984) );
  and2s1 U3068 ( .Q(g7812), .DIN1(n2614), .DIN2(n2061) );
  nnd2s1 U3069 ( .Q(n2614), .DIN1(n2615), .DIN2(n2616) );
  nnd4s1 U3070 ( .Q(n2616), .DIN1(n2617), .DIN2(g1771), .DIN3(g1766), .DIN4(
        n2618) );
  nnd2s1 U3071 ( .Q(n2615), .DIN1(g1776), .DIN2(n2613) );
  nnd2s1 U3072 ( .Q(n2613), .DIN1(n2617), .DIN2(n2568) );
  nor2s1 U3073 ( .Q(g7811), .DIN1(g5653), .DIN2(n2619) );
  xor2s1 U3074 ( .Q(n2619), .DIN1(g1771), .DIN2(n2620) );
  nnd2s1 U3075 ( .Q(n2620), .DIN1(n2617), .DIN2(g1766) );
  nnd2s1 U3076 ( .Q(g7810), .DIN1(n2621), .DIN2(n2061) );
  xor2s1 U3077 ( .Q(n2621), .DIN1(g1766), .DIN2(n2567) );
  and3s1 U3078 ( .Q(g7809), .DIN1(n2622), .DIN2(n2042), .DIN3(g109) );
  nnd2s1 U3079 ( .Q(n2622), .DIN1(n2024), .DIN2(\DFF_452/net739 ) );
  nnd2s1 U3080 ( .Q(g7808), .DIN1(n2623), .DIN2(n2624) );
  nnd2s1 U3081 ( .Q(n2624), .DIN1(g1015), .DIN2(n2070) );
  nnd2s1 U3082 ( .Q(n2623), .DIN1(g1074), .DIN2(n2350) );
  nnd2s1 U3083 ( .Q(g7807), .DIN1(n2625), .DIN2(n2626) );
  nnd2s1 U3084 ( .Q(n2626), .DIN1(g1019), .DIN2(n2068) );
  nnd2s1 U3085 ( .Q(n2625), .DIN1(g1098), .DIN2(n2063) );
  nnd2s1 U3086 ( .Q(g7806), .DIN1(n2627), .DIN2(n2628) );
  nnd2s1 U3087 ( .Q(n2628), .DIN1(g1007), .DIN2(n2069) );
  nnd2s1 U3088 ( .Q(n2627), .DIN1(g1095), .DIN2(n2063) );
  nnd2s1 U3089 ( .Q(g7805), .DIN1(n2629), .DIN2(n2630) );
  nnd2s1 U3090 ( .Q(n2630), .DIN1(g1011), .DIN2(n2070) );
  nnd2s1 U3091 ( .Q(n2629), .DIN1(g1092), .DIN2(n2063) );
  nnd2s1 U3092 ( .Q(g7804), .DIN1(n2631), .DIN2(n2632) );
  nnd2s1 U3093 ( .Q(n2632), .DIN1(g999), .DIN2(n2068) );
  nnd2s1 U3094 ( .Q(n2631), .DIN1(g1089), .DIN2(n2350) );
  nnd2s1 U3095 ( .Q(g7803), .DIN1(n2633), .DIN2(n2634) );
  nnd2s1 U3096 ( .Q(n2634), .DIN1(g1003), .DIN2(n2069) );
  nnd2s1 U3097 ( .Q(n2633), .DIN1(g1086), .DIN2(n2063) );
  nnd2s1 U3098 ( .Q(g7802), .DIN1(n2635), .DIN2(n2636) );
  nnd2s1 U3099 ( .Q(n2636), .DIN1(g991), .DIN2(n2070) );
  nnd2s1 U3100 ( .Q(n2635), .DIN1(g1083), .DIN2(n2350) );
  nnd2s1 U3101 ( .Q(g7801), .DIN1(n2637), .DIN2(n2638) );
  nnd2s1 U3102 ( .Q(n2638), .DIN1(g995), .DIN2(n2068) );
  nnd2s1 U3103 ( .Q(n2637), .DIN1(g1080), .DIN2(n2350) );
  nnd2s1 U3104 ( .Q(g7800), .DIN1(n2639), .DIN2(n2640) );
  nnd2s1 U3105 ( .Q(n2640), .DIN1(g1032), .DIN2(n2069) );
  nnd2s1 U3106 ( .Q(n2639), .DIN1(g1077), .DIN2(n2350) );
  nnd2s1 U3107 ( .Q(g7799), .DIN1(n2641), .DIN2(n2642) );
  nnd2s1 U3108 ( .Q(n2642), .DIN1(g1023), .DIN2(n2070) );
  nnd2s1 U3109 ( .Q(n2641), .DIN1(g1071), .DIN2(n2063) );
  nnd2s1 U3110 ( .Q(g7798), .DIN1(n2643), .DIN2(n2644) );
  nnd2s1 U3111 ( .Q(n2644), .DIN1(g1027), .DIN2(n2068) );
  nnd2s1 U3112 ( .Q(n2643), .DIN1(g1068), .DIN2(n2350) );
  and3s1 U3113 ( .Q(g7786), .DIN1(n2645), .DIN2(n2549), .DIN3(n2440) );
  nnd3s1 U3114 ( .Q(n2549), .DIN1(g4185), .DIN2(g4186), .DIN3(n2646) );
  nnd2s1 U3115 ( .Q(n2645), .DIN1(n2050), .DIN2(n2647) );
  nnd2s1 U3116 ( .Q(n2647), .DIN1(n2646), .DIN2(g4185) );
  and3s1 U3117 ( .Q(g7785), .DIN1(n2648), .DIN2(n2553), .DIN3(n2445) );
  nnd3s1 U3118 ( .Q(n2553), .DIN1(g770), .DIN2(n2649), .DIN3(g774) );
  nnd2s1 U3119 ( .Q(n2648), .DIN1(n2057), .DIN2(n2650) );
  nnd2s1 U3120 ( .Q(n2650), .DIN1(g770), .DIN2(n2649) );
  hi1s1 U3121 ( .Q(n2649), .DIN(n2651) );
  nnd2s1 U3122 ( .Q(g7784), .DIN1(n2034), .DIN2(n2652) );
  nor2s1 U3123 ( .Q(g7783), .DIN1(n2653), .DIN2(n2018) );
  nnd2s1 U3124 ( .Q(g7782), .DIN1(n2035), .DIN2(n2652) );
  nor2s1 U3125 ( .Q(g7781), .DIN1(n2653), .DIN2(n2019) );
  nnd2s1 U3126 ( .Q(g7780), .DIN1(n2036), .DIN2(n2652) );
  nor2s1 U3127 ( .Q(g7779), .DIN1(n2653), .DIN2(n2020) );
  nnd2s1 U3128 ( .Q(g7778), .DIN1(n2037), .DIN2(n2652) );
  nor2s1 U3129 ( .Q(g7777), .DIN1(n2653), .DIN2(n2021) );
  nor2s1 U3130 ( .Q(g7776), .DIN1(n2653), .DIN2(n2022) );
  nor2s1 U3131 ( .Q(g7775), .DIN1(n2653), .DIN2(n2023) );
  nnd2s1 U3132 ( .Q(g7774), .DIN1(n2038), .DIN2(n2652) );
  nnd2s1 U3133 ( .Q(g7773), .DIN1(n2654), .DIN2(n2655) );
  nnd2s1 U3134 ( .Q(n2655), .DIN1(g143), .DIN2(n2656) );
  nnd2s1 U3135 ( .Q(n2654), .DIN1(n2657), .DIN2(g302) );
  nnd2s1 U3136 ( .Q(g7772), .DIN1(n2658), .DIN2(n2659) );
  nnd2s1 U3137 ( .Q(n2659), .DIN1(g166), .DIN2(n2656) );
  nnd2s1 U3138 ( .Q(n2658), .DIN1(n2657), .DIN2(g299) );
  nnd2s1 U3139 ( .Q(g7771), .DIN1(n2660), .DIN2(n2661) );
  nnd2s1 U3140 ( .Q(n2661), .DIN1(g139), .DIN2(n2656) );
  nnd2s1 U3141 ( .Q(n2660), .DIN1(n2657), .DIN2(g296) );
  nnd2s1 U3142 ( .Q(g7770), .DIN1(n2662), .DIN2(n2663) );
  nnd2s1 U3143 ( .Q(n2663), .DIN1(g135), .DIN2(n2656) );
  nnd2s1 U3144 ( .Q(n2662), .DIN1(n2657), .DIN2(g293) );
  nnd2s1 U3145 ( .Q(g7769), .DIN1(n2664), .DIN2(n2665) );
  nnd2s1 U3146 ( .Q(n2665), .DIN1(g131), .DIN2(n2656) );
  nnd2s1 U3147 ( .Q(n2664), .DIN1(n2657), .DIN2(g290) );
  nnd2s1 U3148 ( .Q(g7768), .DIN1(n2666), .DIN2(n2667) );
  nnd2s1 U3149 ( .Q(n2667), .DIN1(g127), .DIN2(n2656) );
  nnd2s1 U3150 ( .Q(n2666), .DIN1(n2657), .DIN2(g287) );
  nnd2s1 U3151 ( .Q(g7767), .DIN1(n2668), .DIN2(n2669) );
  nnd2s1 U3152 ( .Q(n2669), .DIN1(g170), .DIN2(n2656) );
  nnd2s1 U3153 ( .Q(n2668), .DIN1(n2657), .DIN2(g284) );
  nnd2s1 U3154 ( .Q(g7766), .DIN1(n2670), .DIN2(n2671) );
  nnd2s1 U3155 ( .Q(n2671), .DIN1(g174), .DIN2(n2656) );
  nnd2s1 U3156 ( .Q(n2670), .DIN1(n2657), .DIN2(g281) );
  nnd2s1 U3157 ( .Q(g7765), .DIN1(n2672), .DIN2(n2673) );
  nnd2s1 U3158 ( .Q(n2673), .DIN1(g162), .DIN2(n2656) );
  nnd2s1 U3159 ( .Q(n2672), .DIN1(n2657), .DIN2(g278) );
  nnd2s1 U3160 ( .Q(g7764), .DIN1(n2674), .DIN2(n2675) );
  nnd2s1 U3161 ( .Q(n2675), .DIN1(g158), .DIN2(n2656) );
  nnd2s1 U3162 ( .Q(n2674), .DIN1(n2657), .DIN2(g275) );
  nnd2s1 U3163 ( .Q(g7763), .DIN1(n2676), .DIN2(n2677) );
  nnd2s1 U3164 ( .Q(n2677), .DIN1(g153), .DIN2(n2656) );
  nnd2s1 U3165 ( .Q(n2676), .DIN1(n2657), .DIN2(g272) );
  nnd2s1 U3166 ( .Q(g7762), .DIN1(n2678), .DIN2(n2679) );
  nnd2s1 U3167 ( .Q(n2679), .DIN1(g148), .DIN2(n2656) );
  nnd2s1 U3168 ( .Q(n2678), .DIN1(n2657), .DIN2(g269) );
  nnd2s1 U3169 ( .Q(g7761), .DIN1(n2680), .DIN2(n2681) );
  nnd2s1 U3170 ( .Q(n2681), .DIN1(g178), .DIN2(n2656) );
  nnd2s1 U3171 ( .Q(n2680), .DIN1(n2657), .DIN2(g266) );
  nnd2s1 U3172 ( .Q(g7760), .DIN1(n2682), .DIN2(n2683) );
  nnd2s1 U3173 ( .Q(n2683), .DIN1(g182), .DIN2(n2656) );
  nnd2s1 U3174 ( .Q(n2682), .DIN1(n2657), .DIN2(g263) );
  hi1s1 U3175 ( .Q(n2657), .DIN(n2656) );
  nnd2s1 U3176 ( .Q(n2684), .DIN1(n2560), .DIN2(n2017) );
  nnd2s1 U3177 ( .Q(g7759), .DIN1(n2685), .DIN2(n2686) );
  nnd2s1 U3178 ( .Q(n2686), .DIN1(g575), .DIN2(n2072) );
  nnd2s1 U3179 ( .Q(g7758), .DIN1(n2687), .DIN2(n2688) );
  nnd2s1 U3180 ( .Q(n2688), .DIN1(g572), .DIN2(n2072) );
  nnd2s1 U3181 ( .Q(g7757), .DIN1(n2351), .DIN2(n2689) );
  nnd2s1 U3182 ( .Q(n2689), .DIN1(g569), .DIN2(n2082) );
  nnd2s1 U3183 ( .Q(g7756), .DIN1(n2358), .DIN2(n2690) );
  nnd2s1 U3184 ( .Q(n2690), .DIN1(g566), .DIN2(n2072) );
  nnd2s1 U3185 ( .Q(g7755), .DIN1(n2364), .DIN2(n2691) );
  nnd2s1 U3186 ( .Q(n2691), .DIN1(g563), .DIN2(n2082) );
  nnd2s1 U3187 ( .Q(g7754), .DIN1(n2371), .DIN2(n2692) );
  nnd2s1 U3188 ( .Q(n2692), .DIN1(g560), .DIN2(n2082) );
  nnd2s1 U3189 ( .Q(g7753), .DIN1(n2377), .DIN2(n2693) );
  nnd2s1 U3190 ( .Q(n2693), .DIN1(g557), .DIN2(n2072) );
  nnd2s1 U3191 ( .Q(g7752), .DIN1(n2384), .DIN2(n2694) );
  nnd2s1 U3192 ( .Q(n2694), .DIN1(g554), .DIN2(n2072) );
  nnd2s1 U3193 ( .Q(g7751), .DIN1(n2695), .DIN2(n2696) );
  nnd2s1 U3194 ( .Q(n2696), .DIN1(g549), .DIN2(n2082) );
  nnd2s1 U3195 ( .Q(g7750), .DIN1(n2390), .DIN2(n2697) );
  nnd2s1 U3196 ( .Q(n2697), .DIN1(g546), .DIN2(n2072) );
  and2s1 U3197 ( .Q(g7749), .DIN1(g178), .DIN2(g109) );
  nnd2s1 U3198 ( .Q(g7746), .DIN1(n2698), .DIN2(n2699) );
  nnd2s1 U3199 ( .Q(n2699), .DIN1(n2700), .DIN2(g7748) );
  nor2s1 U3200 ( .Q(g7748), .DIN1(n1926), .DIN2(n2065) );
  xor2s1 U3201 ( .Q(n2700), .DIN1(n2701), .DIN2(n1925) );
  nnd3s1 U3202 ( .Q(n2698), .DIN1(n2702), .DIN2(n2703), .DIN3(n1926) );
  nnd2s1 U3203 ( .Q(n2703), .DIN1(n2701), .DIN2(n2704) );
  nnd2s1 U3204 ( .Q(n2704), .DIN1(g109), .DIN2(n1925) );
  or2s1 U3205 ( .Q(n2702), .DIN1(n2701), .DIN2(g7747) );
  nor2s1 U3206 ( .Q(g7747), .DIN1(n1925), .DIN2(n2065) );
  xor2s1 U3207 ( .Q(n2701), .DIN1(g153), .DIN2(g182) );
  nnd2s1 U3208 ( .Q(g7745), .DIN1(n2705), .DIN2(n2706) );
  nnd2s1 U3209 ( .Q(n2706), .DIN1(g119), .DIN2(g109) );
  nnd2s1 U3210 ( .Q(g7366), .DIN1(n2707), .DIN2(n1998) );
  nnd2s1 U3211 ( .Q(g7365), .DIN1(n2708), .DIN2(n2709) );
  nnd2s1 U3212 ( .Q(n2709), .DIN1(g1448), .DIN2(n2710) );
  nnd2s1 U3213 ( .Q(n2708), .DIN1(n2711), .DIN2(g1607) );
  nnd2s1 U3214 ( .Q(g7364), .DIN1(n2712), .DIN2(n2713) );
  nnd2s1 U3215 ( .Q(n2713), .DIN1(g1444), .DIN2(n2710) );
  nnd2s1 U3216 ( .Q(n2712), .DIN1(n2711), .DIN2(g1604) );
  nnd2s1 U3217 ( .Q(g7363), .DIN1(n2714), .DIN2(n2715) );
  nnd2s1 U3218 ( .Q(n2715), .DIN1(g1440), .DIN2(n2710) );
  nnd2s1 U3219 ( .Q(n2714), .DIN1(n2711), .DIN2(g1601) );
  nnd2s1 U3220 ( .Q(g7362), .DIN1(n2716), .DIN2(n2717) );
  nnd2s1 U3221 ( .Q(n2717), .DIN1(g1436), .DIN2(n2710) );
  nnd2s1 U3222 ( .Q(n2716), .DIN1(n2711), .DIN2(g1598) );
  nnd2s1 U3223 ( .Q(g7361), .DIN1(n2718), .DIN2(n2719) );
  nnd2s1 U3224 ( .Q(n2719), .DIN1(g1432), .DIN2(n2710) );
  nnd2s1 U3225 ( .Q(n2718), .DIN1(n2711), .DIN2(g1595) );
  nnd2s1 U3226 ( .Q(g7360), .DIN1(n2720), .DIN2(n2721) );
  nnd2s1 U3227 ( .Q(n2721), .DIN1(g1403), .DIN2(n2710) );
  nnd2s1 U3228 ( .Q(n2720), .DIN1(n2711), .DIN2(g1592) );
  nnd2s1 U3229 ( .Q(g7359), .DIN1(n2722), .DIN2(n2723) );
  nnd2s1 U3230 ( .Q(n2723), .DIN1(g1428), .DIN2(n2710) );
  nnd2s1 U3231 ( .Q(n2722), .DIN1(n2711), .DIN2(g1589) );
  nnd2s1 U3232 ( .Q(g7358), .DIN1(n2724), .DIN2(n2725) );
  nnd2s1 U3233 ( .Q(n2725), .DIN1(g1407), .DIN2(n2710) );
  nnd2s1 U3234 ( .Q(n2724), .DIN1(n2711), .DIN2(g1586) );
  nnd2s1 U3235 ( .Q(g7357), .DIN1(n2726), .DIN2(n2727) );
  nnd2s1 U3236 ( .Q(n2727), .DIN1(g1424), .DIN2(n2710) );
  nnd2s1 U3237 ( .Q(n2726), .DIN1(n2711), .DIN2(g1583) );
  nnd2s1 U3238 ( .Q(g7356), .DIN1(n2728), .DIN2(n2729) );
  nnd2s1 U3239 ( .Q(n2729), .DIN1(g1411), .DIN2(n2710) );
  nnd2s1 U3240 ( .Q(n2728), .DIN1(n2711), .DIN2(g1580) );
  nnd2s1 U3241 ( .Q(g7355), .DIN1(n2730), .DIN2(n2731) );
  nnd2s1 U3242 ( .Q(n2731), .DIN1(g1419), .DIN2(n2710) );
  nnd2s1 U3243 ( .Q(n2730), .DIN1(n2711), .DIN2(g1577) );
  nnd2s1 U3244 ( .Q(g7354), .DIN1(n2732), .DIN2(n2733) );
  nnd2s1 U3245 ( .Q(n2733), .DIN1(g1515), .DIN2(n2710) );
  nnd2s1 U3246 ( .Q(n2732), .DIN1(n2711), .DIN2(g1574) );
  nnd2s1 U3247 ( .Q(g7353), .DIN1(n2734), .DIN2(n2735) );
  nnd2s1 U3248 ( .Q(n2735), .DIN1(g1520), .DIN2(n2710) );
  nnd2s1 U3249 ( .Q(n2734), .DIN1(n2711), .DIN2(g1571) );
  nnd2s1 U3250 ( .Q(g7352), .DIN1(n2736), .DIN2(n2737) );
  nnd2s1 U3251 ( .Q(n2737), .DIN1(g1415), .DIN2(n2710) );
  nnd2s1 U3252 ( .Q(n2736), .DIN1(n2711), .DIN2(g1567) );
  hi1s1 U3253 ( .Q(n2711), .DIN(n2710) );
  nnd2s1 U3254 ( .Q(g7351), .DIN1(n2739), .DIN2(n2740) );
  nnd2s1 U3255 ( .Q(n2740), .DIN1(g1453), .DIN2(n2741) );
  nnd2s1 U3256 ( .Q(n2739), .DIN1(n2742), .DIN2(g1564) );
  nnd2s1 U3257 ( .Q(g7350), .DIN1(n2743), .DIN2(n2744) );
  nnd2s1 U3258 ( .Q(n2744), .DIN1(g1458), .DIN2(n2741) );
  nnd2s1 U3259 ( .Q(n2743), .DIN1(n2742), .DIN2(g1561) );
  nnd2s1 U3260 ( .Q(g7349), .DIN1(n2745), .DIN2(n2746) );
  nnd2s1 U3261 ( .Q(n2746), .DIN1(g1462), .DIN2(n2741) );
  nnd2s1 U3262 ( .Q(n2745), .DIN1(n2742), .DIN2(g1558) );
  nnd2s1 U3263 ( .Q(g7348), .DIN1(n2747), .DIN2(n2748) );
  nnd2s1 U3264 ( .Q(n2748), .DIN1(g1466), .DIN2(n2741) );
  nnd2s1 U3265 ( .Q(n2747), .DIN1(n2742), .DIN2(g1555) );
  nnd2s1 U3266 ( .Q(g7347), .DIN1(n2749), .DIN2(n2750) );
  nnd2s1 U3267 ( .Q(n2750), .DIN1(g1470), .DIN2(n2741) );
  nnd2s1 U3268 ( .Q(n2749), .DIN1(n2742), .DIN2(g1552) );
  nnd2s1 U3269 ( .Q(g7346), .DIN1(n2751), .DIN2(n2752) );
  nnd2s1 U3270 ( .Q(n2752), .DIN1(g1474), .DIN2(n2741) );
  nnd2s1 U3271 ( .Q(n2751), .DIN1(n2742), .DIN2(g1549) );
  nnd2s1 U3272 ( .Q(g7345), .DIN1(n2753), .DIN2(n2754) );
  nnd2s1 U3273 ( .Q(n2754), .DIN1(g1478), .DIN2(n2741) );
  nnd2s1 U3274 ( .Q(n2753), .DIN1(n2742), .DIN2(g1546) );
  nnd2s1 U3275 ( .Q(g7344), .DIN1(n2755), .DIN2(n2756) );
  nnd2s1 U3276 ( .Q(n2756), .DIN1(g1482), .DIN2(n2741) );
  nnd2s1 U3277 ( .Q(n2755), .DIN1(n2742), .DIN2(g1543) );
  nnd2s1 U3278 ( .Q(g7343), .DIN1(n2757), .DIN2(n2758) );
  nnd2s1 U3279 ( .Q(n2758), .DIN1(g1486), .DIN2(n2741) );
  nnd2s1 U3280 ( .Q(n2757), .DIN1(n2742), .DIN2(g1540) );
  nnd2s1 U3281 ( .Q(g7342), .DIN1(n2759), .DIN2(n2760) );
  nnd2s1 U3282 ( .Q(n2760), .DIN1(g1490), .DIN2(n2741) );
  nnd2s1 U3283 ( .Q(n2759), .DIN1(n2742), .DIN2(g1537) );
  nnd2s1 U3284 ( .Q(g7341), .DIN1(n2761), .DIN2(n2762) );
  nnd2s1 U3285 ( .Q(n2762), .DIN1(g1494), .DIN2(n2741) );
  nnd2s1 U3286 ( .Q(n2761), .DIN1(n2742), .DIN2(g1534) );
  nnd2s1 U3287 ( .Q(g7340), .DIN1(n2763), .DIN2(n2764) );
  nnd2s1 U3288 ( .Q(n2764), .DIN1(g1499), .DIN2(n2741) );
  nnd2s1 U3289 ( .Q(n2763), .DIN1(n2742), .DIN2(g1531) );
  nnd2s1 U3290 ( .Q(g7339), .DIN1(n2765), .DIN2(n2766) );
  nnd2s1 U3291 ( .Q(n2766), .DIN1(g1504), .DIN2(n2741) );
  nnd2s1 U3292 ( .Q(n2765), .DIN1(n2742), .DIN2(g1528) );
  nnd2s1 U3293 ( .Q(g7338), .DIN1(n2767), .DIN2(n2768) );
  nnd2s1 U3294 ( .Q(n2768), .DIN1(g1508), .DIN2(n2741) );
  nnd2s1 U3295 ( .Q(n2767), .DIN1(n2742), .DIN2(g1524) );
  hi1s1 U3296 ( .Q(n2742), .DIN(n2741) );
  nor2s1 U3297 ( .Q(n2738), .DIN1(n2064), .DIN2(n2575) );
  nor2s1 U3298 ( .Q(n2575), .DIN1(n2769), .DIN2(g12) );
  hi1s1 U3299 ( .Q(n2769), .DIN(n2560) );
  nnd2s1 U3300 ( .Q(g7337), .DIN1(n2705), .DIN2(n2770) );
  nnd2s1 U3301 ( .Q(n2770), .DIN1(g12), .DIN2(g109) );
  nnd2s1 U3302 ( .Q(g7336), .DIN1(n2705), .DIN2(n2771) );
  nnd2s1 U3303 ( .Q(n2771), .DIN1(g9), .DIN2(g109) );
  nnd2s1 U3304 ( .Q(n2705), .DIN1(n2560), .DIN2(g109) );
  nor2s1 U3305 ( .Q(n2560), .DIN1(n2042), .DIN2(n2072) );
  and2s1 U3306 ( .Q(g7335), .DIN1(g1520), .DIN2(g109) );
  and2s1 U3307 ( .Q(g7334), .DIN1(g109), .DIN2(g1515) );
  and2s1 U3308 ( .Q(g7333), .DIN1(g109), .DIN2(g1419) );
  and2s1 U3309 ( .Q(g7332), .DIN1(g109), .DIN2(g1411) );
  and2s1 U3310 ( .Q(g7331), .DIN1(g109), .DIN2(g1424) );
  and2s1 U3311 ( .Q(g7330), .DIN1(g109), .DIN2(g1407) );
  and2s1 U3312 ( .Q(g7329), .DIN1(g1504), .DIN2(g109) );
  and2s1 U3313 ( .Q(g7328), .DIN1(g109), .DIN2(g1499) );
  nnd2s1 U3314 ( .Q(g7326), .DIN1(n2772), .DIN2(n2773) );
  nnd2s1 U3315 ( .Q(n2773), .DIN1(g7327), .DIN2(n2774) );
  hi1s1 U3316 ( .Q(n2774), .DIN(n2775) );
  nor2s1 U3317 ( .Q(g7327), .DIN1(n2012), .DIN2(n2065) );
  nnd3s1 U3318 ( .Q(n2772), .DIN1(g109), .DIN2(n2012), .DIN3(n2775) );
  xor2s1 U3319 ( .Q(n2775), .DIN1(n2776), .DIN2(g1494) );
  xor2s1 U3320 ( .Q(n2776), .DIN1(g1508), .DIN2(g1499) );
  nor2s1 U3321 ( .Q(g7325), .DIN1(n2064), .DIN2(n1973) );
  nor2s1 U3322 ( .Q(g7324), .DIN1(n2066), .DIN2(n1963) );
  and2s1 U3323 ( .Q(g7323), .DIN1(g109), .DIN2(g1397) );
  nor2s1 U3324 ( .Q(g7322), .DIN1(n2066), .DIN2(n1946) );
  nor2s1 U3325 ( .Q(g7321), .DIN1(n2777), .DIN2(n2024) );
  hi1s1 U3326 ( .Q(g7320), .DIN(n2777) );
  nnd2s1 U3327 ( .Q(n2777), .DIN1(g6825), .DIN2(n2778) );
  and2s1 U3328 ( .Q(g7319), .DIN1(g109), .DIN2(g1365) );
  nor2s1 U3329 ( .Q(g7318), .DIN1(n2041), .DIN2(n2065) );
  nor2s1 U3330 ( .Q(g7317), .DIN1(n2066), .DIN2(n1964) );
  nor2s1 U3331 ( .Q(g7316), .DIN1(n2064), .DIN2(n2001) );
  nor2s1 U3332 ( .Q(g7315), .DIN1(n2064), .DIN2(n2004) );
  nor2s1 U3333 ( .Q(g7314), .DIN1(n2067), .DIN2(n1962) );
  nor2s1 U3334 ( .Q(g7313), .DIN1(n2064), .DIN2(n1941) );
  nor2s1 U3335 ( .Q(g7312), .DIN1(n2066), .DIN2(n1972) );
  nor2s1 U3336 ( .Q(g7311), .DIN1(n2066), .DIN2(n2040) );
  nor2s1 U3337 ( .Q(g7310), .DIN1(n2067), .DIN2(n2003) );
  nor2s1 U3338 ( .Q(g7309), .DIN1(n2067), .DIN2(n1940) );
  nor2s1 U3339 ( .Q(g7308), .DIN1(n2067), .DIN2(n1947) );
  nor2s1 U3340 ( .Q(g7307), .DIN1(n2067), .DIN2(n1939) );
  and2s1 U3341 ( .Q(g7306), .DIN1(g109), .DIN2(g1362) );
  nor2s1 U3342 ( .Q(g7305), .DIN1(n2067), .DIN2(n2002) );
  nnd3s1 U3343 ( .Q(g7304), .DIN1(n2779), .DIN2(n2780), .DIN3(n2781) );
  nnd3s1 U3344 ( .Q(n2781), .DIN1(n2782), .DIN2(n1931), .DIN3(g6825) );
  nnd3s1 U3345 ( .Q(n2780), .DIN1(g6836), .DIN2(n2783), .DIN3(g201) );
  nnd2s1 U3346 ( .Q(n2779), .DIN1(n2784), .DIN2(n1995) );
  nnd2s1 U3347 ( .Q(n2784), .DIN1(n2785), .DIN2(n2786) );
  nnd2s1 U3348 ( .Q(n2786), .DIN1(g6836), .DIN2(n2782) );
  nnd3s1 U3349 ( .Q(n2785), .DIN1(g109), .DIN2(n1931), .DIN3(n2783) );
  hi1s1 U3350 ( .Q(n2783), .DIN(n2782) );
  xor2s1 U3351 ( .Q(n2782), .DIN1(n2787), .DIN2(g1389) );
  nor2s1 U3352 ( .Q(n2787), .DIN1(n2788), .DIN2(g1386) );
  and2s1 U3353 ( .Q(n2788), .DIN1(n1995), .DIN2(n2778) );
  nor4s1 U3354 ( .Q(n2778), .DIN1(n2789), .DIN2(n2790), .DIN3(n2791), .DIN4(
        n2792) );
  nnd4s1 U3355 ( .Q(n2792), .DIN1(n2001), .DIN2(n1962), .DIN3(n1931), .DIN4(
        n2793) );
  and3s1 U3356 ( .Q(n2793), .DIN1(n2041), .DIN2(n1946), .DIN3(n1973) );
  nnd4s1 U3357 ( .Q(n2791), .DIN1(n2002), .DIN2(n1963), .DIN3(n1939), .DIN4(
        n2794) );
  and3s1 U3358 ( .Q(n2794), .DIN1(n2040), .DIN2(n1947), .DIN3(n1972) );
  nnd4s1 U3359 ( .Q(n2790), .DIN1(n2003), .DIN2(n1965), .DIN3(n1940), .DIN4(
        n2795) );
  nor2s1 U3360 ( .Q(n2795), .DIN1(g1365), .DIN2(g1362) );
  nnd4s1 U3361 ( .Q(n2789), .DIN1(n2004), .DIN2(n1964), .DIN3(n1941), .DIN4(
        n2796) );
  nor3s1 U3362 ( .Q(n2796), .DIN1(g1389), .DIN2(g1397), .DIN3(g1386) );
  nnd2s1 U3363 ( .Q(g7303), .DIN1(n2797), .DIN2(n2798) );
  nnd2s1 U3364 ( .Q(n2798), .DIN1(g1270), .DIN2(n2060) );
  nnd2s1 U3365 ( .Q(n2797), .DIN1(g1265), .DIN2(n2799) );
  nnd2s1 U3366 ( .Q(g7302), .DIN1(n2800), .DIN2(n2801) );
  nnd2s1 U3367 ( .Q(n2801), .DIN1(g1265), .DIN2(n2060) );
  nnd2s1 U3368 ( .Q(n2800), .DIN1(g1260), .DIN2(n2799) );
  nnd2s1 U3369 ( .Q(g7301), .DIN1(n2802), .DIN2(n2803) );
  nnd2s1 U3370 ( .Q(n2803), .DIN1(g1260), .DIN2(n2060) );
  nnd2s1 U3371 ( .Q(n2802), .DIN1(g1255), .DIN2(n2799) );
  nnd2s1 U3372 ( .Q(g7300), .DIN1(n2804), .DIN2(n2805) );
  nnd2s1 U3373 ( .Q(n2805), .DIN1(g1255), .DIN2(n2060) );
  nnd2s1 U3374 ( .Q(n2804), .DIN1(g1250), .DIN2(n2799) );
  nnd2s1 U3375 ( .Q(g7299), .DIN1(n2806), .DIN2(n2807) );
  nnd2s1 U3376 ( .Q(n2807), .DIN1(g1250), .DIN2(n2060) );
  nnd2s1 U3377 ( .Q(n2806), .DIN1(g1245), .DIN2(n2799) );
  nnd2s1 U3378 ( .Q(g7298), .DIN1(n2808), .DIN2(n2809) );
  nnd2s1 U3379 ( .Q(n2809), .DIN1(g1245), .DIN2(n2060) );
  nnd2s1 U3380 ( .Q(n2808), .DIN1(g1240), .DIN2(n2799) );
  nnd2s1 U3381 ( .Q(g7297), .DIN1(n2810), .DIN2(n2811) );
  nnd2s1 U3382 ( .Q(n2811), .DIN1(g1240), .DIN2(n2060) );
  nnd2s1 U3383 ( .Q(n2810), .DIN1(g1235), .DIN2(n2799) );
  nnd2s1 U3384 ( .Q(g7296), .DIN1(n2812), .DIN2(n2813) );
  nnd2s1 U3385 ( .Q(n2813), .DIN1(g1235), .DIN2(n2060) );
  nnd2s1 U3386 ( .Q(n2812), .DIN1(g1275), .DIN2(n2799) );
  nnd2s1 U3387 ( .Q(g7295), .DIN1(n2814), .DIN2(n2815) );
  nnd2s1 U3388 ( .Q(n2815), .DIN1(g1280), .DIN2(n2060) );
  nnd2s1 U3389 ( .Q(n2814), .DIN1(g1284), .DIN2(n2799) );
  nnd2s1 U3390 ( .Q(g7294), .DIN1(n2816), .DIN2(n2817) );
  nnd2s1 U3391 ( .Q(n2817), .DIN1(g1284), .DIN2(n2060) );
  nnd2s1 U3392 ( .Q(n2816), .DIN1(g1292), .DIN2(n2799) );
  nnd2s1 U3393 ( .Q(g7293), .DIN1(n2818), .DIN2(n2819) );
  nnd2s1 U3394 ( .Q(n2819), .DIN1(g1292), .DIN2(n2060) );
  nnd2s1 U3395 ( .Q(n2818), .DIN1(g1296), .DIN2(n2799) );
  nnd2s1 U3396 ( .Q(g7292), .DIN1(n2820), .DIN2(n2821) );
  nnd2s1 U3397 ( .Q(n2821), .DIN1(g1296), .DIN2(n2060) );
  nnd2s1 U3398 ( .Q(n2820), .DIN1(g1300), .DIN2(n2799) );
  nnd2s1 U3399 ( .Q(g7291), .DIN1(n2822), .DIN2(n2823) );
  nnd2s1 U3400 ( .Q(n2823), .DIN1(g1300), .DIN2(n2060) );
  nnd2s1 U3401 ( .Q(n2822), .DIN1(g1304), .DIN2(n2799) );
  nnd2s1 U3402 ( .Q(g7290), .DIN1(n2824), .DIN2(n2825) );
  nnd2s1 U3403 ( .Q(n2825), .DIN1(g1304), .DIN2(n2060) );
  nnd2s1 U3404 ( .Q(n2824), .DIN1(g1270), .DIN2(n2799) );
  and2s1 U3405 ( .Q(g7289), .DIN1(n2826), .DIN2(n2440) );
  xor2s1 U3406 ( .Q(n2826), .DIN1(n2646), .DIN2(g4185) );
  nor2s1 U3407 ( .Q(g7288), .DIN1(n2827), .DIN2(n2481) );
  xor2s1 U3408 ( .Q(n2827), .DIN1(g770), .DIN2(n2651) );
  nnd2s1 U3409 ( .Q(g7287), .DIN1(n2828), .DIN2(n1997) );
  nor2s1 U3410 ( .Q(g7285), .DIN1(n2829), .DIN2(n2830) );
  nor2s1 U3411 ( .Q(n2830), .DIN1(n2066), .DIN2(n2437) );
  hi1s1 U3412 ( .Q(n2437), .DIN(g881) );
  hi1s1 U3413 ( .Q(n2829), .DIN(n2438) );
  and2s1 U3414 ( .Q(g6845), .DIN1(n2567), .DIN2(g1610) );
  nnd2s1 U3415 ( .Q(g6844), .DIN1(n2831), .DIN2(n2832) );
  nnd3s1 U3416 ( .Q(n2832), .DIN1(g1707), .DIN2(g1700), .DIN3(n2074) );
  nnd2s1 U3417 ( .Q(n2831), .DIN1(g4907), .DIN2(n2075) );
  nor3s1 U3418 ( .Q(g6843), .DIN1(n2350), .DIN2(g4901), .DIN3(n2833) );
  and2s1 U3419 ( .Q(g6837), .DIN1(g109), .DIN2(g1389) );
  nor2s1 U3420 ( .Q(g6836), .DIN1(n1931), .DIN2(n2065) );
  nor2s1 U3421 ( .Q(g6835), .DIN1(n2066), .DIN2(n1965) );
  nor2s1 U3422 ( .Q(g6825), .DIN1(n1995), .DIN2(n2065) );
  nor2s1 U3423 ( .Q(g6818), .DIN1(n2834), .DIN2(n2835) );
  nor2s1 U3424 ( .Q(n2835), .DIN1(n2067), .DIN2(n2011) );
  nor2s1 U3425 ( .Q(g6817), .DIN1(n1949), .DIN2(n2836) );
  nor2s1 U3426 ( .Q(g6816), .DIN1(n1929), .DIN2(n2836) );
  nor2s1 U3427 ( .Q(g6815), .DIN1(n1976), .DIN2(n2836) );
  nor2s1 U3428 ( .Q(g6814), .DIN1(n1974), .DIN2(n2836) );
  nnd2s1 U3429 ( .Q(n2836), .DIN1(g109), .DIN2(\DFF_126/net413 ) );
  nnd2s1 U3430 ( .Q(g6813), .DIN1(n2837), .DIN2(n2838) );
  nnd2s1 U3431 ( .Q(n2838), .DIN1(g1074), .DIN2(n2839) );
  nnd2s1 U3432 ( .Q(n2837), .DIN1(g342), .DIN2(n2840) );
  nnd2s1 U3433 ( .Q(g6812), .DIN1(n2841), .DIN2(n2842) );
  nnd2s1 U3434 ( .Q(n2842), .DIN1(g1098), .DIN2(n2839) );
  nnd2s1 U3435 ( .Q(n2841), .DIN1(g366), .DIN2(n2840) );
  nnd2s1 U3436 ( .Q(g6811), .DIN1(n2843), .DIN2(n2844) );
  nnd2s1 U3437 ( .Q(n2844), .DIN1(g1095), .DIN2(n2839) );
  nnd2s1 U3438 ( .Q(n2843), .DIN1(g363), .DIN2(n2840) );
  nnd2s1 U3439 ( .Q(g6810), .DIN1(n2845), .DIN2(n2846) );
  nnd2s1 U3440 ( .Q(n2846), .DIN1(g1092), .DIN2(n2839) );
  nnd2s1 U3441 ( .Q(n2845), .DIN1(g360), .DIN2(n2840) );
  nnd2s1 U3442 ( .Q(g6809), .DIN1(n2847), .DIN2(n2848) );
  nnd2s1 U3443 ( .Q(n2848), .DIN1(g1089), .DIN2(n2839) );
  nnd2s1 U3444 ( .Q(n2847), .DIN1(g357), .DIN2(n2840) );
  nnd2s1 U3445 ( .Q(g6808), .DIN1(n2849), .DIN2(n2850) );
  nnd2s1 U3446 ( .Q(n2850), .DIN1(g1086), .DIN2(n2839) );
  nnd2s1 U3447 ( .Q(n2849), .DIN1(g354), .DIN2(n2840) );
  nnd2s1 U3448 ( .Q(g6807), .DIN1(n2851), .DIN2(n2852) );
  nnd2s1 U3449 ( .Q(n2852), .DIN1(g1083), .DIN2(n2839) );
  nnd2s1 U3450 ( .Q(n2851), .DIN1(g351), .DIN2(n2840) );
  nnd2s1 U3451 ( .Q(g6806), .DIN1(n2853), .DIN2(n2854) );
  nnd2s1 U3452 ( .Q(n2854), .DIN1(g1080), .DIN2(n2839) );
  nnd2s1 U3453 ( .Q(n2853), .DIN1(g348), .DIN2(n2840) );
  nnd2s1 U3454 ( .Q(g6805), .DIN1(n2855), .DIN2(n2856) );
  nnd2s1 U3455 ( .Q(n2856), .DIN1(g1077), .DIN2(n2839) );
  nnd2s1 U3456 ( .Q(n2855), .DIN1(g345), .DIN2(n2840) );
  nnd2s1 U3457 ( .Q(g6804), .DIN1(n2857), .DIN2(n2858) );
  nnd2s1 U3458 ( .Q(n2858), .DIN1(g1071), .DIN2(n2839) );
  nnd2s1 U3459 ( .Q(n2857), .DIN1(g339), .DIN2(n2840) );
  nnd2s1 U3460 ( .Q(g6803), .DIN1(n2859), .DIN2(n2860) );
  nnd2s1 U3461 ( .Q(n2860), .DIN1(g1068), .DIN2(n2839) );
  nnd2s1 U3462 ( .Q(n2859), .DIN1(g336), .DIN2(n2840) );
  nor2s1 U3463 ( .Q(g6802), .DIN1(n2646), .DIN2(n2861) );
  nor2s1 U3464 ( .Q(n2861), .DIN1(n2862), .DIN2(n2863) );
  nor2s1 U3465 ( .Q(n2863), .DIN1(g6800), .DIN2(n1990) );
  nor2s1 U3466 ( .Q(n2862), .DIN1(n1999), .DIN2(n2479) );
  nor2s1 U3467 ( .Q(n2646), .DIN1(n2406), .DIN2(n1999) );
  nnd2s1 U3468 ( .Q(n2406), .DIN1(g4183), .DIN2(g4182) );
  nnd2s1 U3469 ( .Q(g6801), .DIN1(n2864), .DIN2(n2440) );
  xor2s1 U3470 ( .Q(n2864), .DIN1(n1990), .DIN2(g4182) );
  nnd2s1 U3471 ( .Q(g6800), .DIN1(n2440), .DIN2(g4182) );
  hi1s1 U3472 ( .Q(n2440), .DIN(n2479) );
  nnd3s1 U3473 ( .Q(n2479), .DIN1(g2639), .DIN2(g109), .DIN3(g745) );
  and3s1 U3474 ( .Q(g6799), .DIN1(n2865), .DIN2(n2651), .DIN3(n2445) );
  nnd3s1 U3475 ( .Q(n2651), .DIN1(g762), .DIN2(g758), .DIN3(g766) );
  nnd2s1 U3476 ( .Q(n2865), .DIN1(n2058), .DIN2(n2866) );
  nnd2s1 U3477 ( .Q(n2866), .DIN1(g762), .DIN2(g758) );
  nnd2s1 U3478 ( .Q(g6798), .DIN1(n2867), .DIN2(n2868) );
  nnd3s1 U3479 ( .Q(n2868), .DIN1(n2445), .DIN2(g758), .DIN3(n2051) );
  nnd2s1 U3480 ( .Q(n2867), .DIN1(g6797), .DIN2(g762) );
  nor2s1 U3481 ( .Q(g6797), .DIN1(n2481), .DIN2(g758) );
  hi1s1 U3482 ( .Q(n2481), .DIN(n2445) );
  nor2s1 U3483 ( .Q(n2445), .DIN1(n2064), .DIN2(g590) );
  nor4s1 U3484 ( .Q(g6339), .DIN1(n2869), .DIN2(n2870), .DIN3(n2025), .DIN4(
        n1952) );
  nnd3s1 U3485 ( .Q(n2870), .DIN1(n2568), .DIN2(n1984), .DIN3(g1786) );
  hi1s1 U3486 ( .Q(n2568), .DIN(n2618) );
  nnd3s1 U3487 ( .Q(n2618), .DIN1(g1771), .DIN2(g1766), .DIN3(g1776) );
  nnd4s1 U3488 ( .Q(n2869), .DIN1(g1707), .DIN2(g1690), .DIN3(g1806), .DIN4(
        g1801) );
  nnd2s1 U3489 ( .Q(g6337), .DIN1(n2871), .DIN2(n2872) );
  nnd2s1 U3490 ( .Q(n2872), .DIN1(g1718), .DIN2(n2069) );
  nnd2s1 U3491 ( .Q(n2871), .DIN1(g5653), .DIN2(n2350) );
  nnd2s1 U3492 ( .Q(g6336), .DIN1(n2873), .DIN2(n2874) );
  nnd2s1 U3493 ( .Q(n2874), .DIN1(g5653), .DIN2(n2070) );
  nnd2s1 U3494 ( .Q(n2873), .DIN1(g1710), .DIN2(n2350) );
  and2s1 U3495 ( .Q(g6330), .DIN1(n2068), .DIN2(g1357) );
  nor2s1 U3496 ( .Q(g6313), .DIN1(n2064), .DIN2(n1934) );
  nor2s1 U3497 ( .Q(g6312), .DIN1(n2066), .DIN2(n1970) );
  nor2s1 U3498 ( .Q(g6311), .DIN1(n2067), .DIN2(n1944) );
  nor2s1 U3499 ( .Q(g6310), .DIN1(n2064), .DIN2(n2013) );
  nor2s1 U3500 ( .Q(g6309), .DIN1(n2064), .DIN2(n1971) );
  nor2s1 U3501 ( .Q(g6308), .DIN1(n2066), .DIN2(n1945) );
  nor2s1 U3502 ( .Q(g6307), .DIN1(n2067), .DIN2(n2014) );
  nor2s1 U3503 ( .Q(g6306), .DIN1(n2015), .DIN2(n2065) );
  nor2s1 U3504 ( .Q(g6305), .DIN1(n2065), .DIN2(n2016) );
  nor2s1 U3505 ( .Q(g6304), .DIN1(n2067), .DIN2(n1988) );
  nor2s1 U3506 ( .Q(g6303), .DIN1(n2064), .DIN2(n2005) );
  nor2s1 U3507 ( .Q(g6302), .DIN1(n2066), .DIN2(n1966) );
  nor2s1 U3508 ( .Q(g6301), .DIN1(n2067), .DIN2(n1942) );
  nor2s1 U3509 ( .Q(g6300), .DIN1(n2064), .DIN2(n1927) );
  nor2s1 U3510 ( .Q(g6299), .DIN1(n2066), .DIN2(n1969) );
  nor2s1 U3511 ( .Q(g5673), .DIN1(g4906), .DIN2(\DFF_489/net776 ) );
  nor2s1 U3512 ( .Q(g5671), .DIN1(g4906), .DIN2(\DFF_330/net617 ) );
  nor2s1 U3513 ( .Q(g5670), .DIN1(g4906), .DIN2(\DFF_385/net672 ) );
  nnd2s1 U3514 ( .Q(g5669), .DIN1(n2875), .DIN2(n2876) );
  nnd2s1 U3515 ( .Q(n2876), .DIN1(g1762), .DIN2(n2877) );
  nnd2s1 U3516 ( .Q(n2875), .DIN1(n2878), .DIN2(g1806) );
  nnd2s1 U3517 ( .Q(g5668), .DIN1(n2879), .DIN2(n2880) );
  nnd2s1 U3518 ( .Q(n2880), .DIN1(g1759), .DIN2(n2877) );
  nnd2s1 U3519 ( .Q(n2879), .DIN1(n2878), .DIN2(g1801) );
  nnd2s1 U3520 ( .Q(g5667), .DIN1(n2881), .DIN2(n2882) );
  nnd2s1 U3521 ( .Q(n2882), .DIN1(g1756), .DIN2(n2877) );
  nnd2s1 U3522 ( .Q(n2881), .DIN1(n2878), .DIN2(g1796) );
  nnd2s1 U3523 ( .Q(g5666), .DIN1(n2883), .DIN2(n2884) );
  nnd2s1 U3524 ( .Q(n2884), .DIN1(g1753), .DIN2(n2877) );
  nnd2s1 U3525 ( .Q(n2883), .DIN1(n2878), .DIN2(g1791) );
  nnd2s1 U3526 ( .Q(g5665), .DIN1(n2885), .DIN2(n2886) );
  nnd2s1 U3527 ( .Q(n2886), .DIN1(g1750), .DIN2(n2877) );
  nnd2s1 U3528 ( .Q(n2885), .DIN1(n2878), .DIN2(g1786) );
  nnd2s1 U3529 ( .Q(g5664), .DIN1(n2887), .DIN2(n2888) );
  nnd2s1 U3530 ( .Q(n2888), .DIN1(g1747), .DIN2(n2877) );
  nnd2s1 U3531 ( .Q(n2887), .DIN1(n2878), .DIN2(g1781) );
  nnd2s1 U3532 ( .Q(g5663), .DIN1(n2889), .DIN2(n2890) );
  nnd2s1 U3533 ( .Q(n2890), .DIN1(g1744), .DIN2(n2877) );
  nnd2s1 U3534 ( .Q(n2889), .DIN1(n2878), .DIN2(g1776) );
  nnd2s1 U3535 ( .Q(g5662), .DIN1(n2891), .DIN2(n2892) );
  nnd2s1 U3536 ( .Q(n2892), .DIN1(g1741), .DIN2(n2877) );
  nnd2s1 U3537 ( .Q(n2891), .DIN1(n2878), .DIN2(g1771) );
  nnd2s1 U3538 ( .Q(g5661), .DIN1(n2893), .DIN2(n2894) );
  nnd2s1 U3539 ( .Q(n2894), .DIN1(g1738), .DIN2(n2877) );
  nnd2s1 U3540 ( .Q(n2893), .DIN1(n2878), .DIN2(g1766) );
  hi1s1 U3541 ( .Q(n2878), .DIN(n2877) );
  or2s1 U3542 ( .Q(g5660), .DIN1(g1289), .DIN2(g1212) );
  nor2s1 U3543 ( .Q(g5657), .DIN1(g4894), .DIN2(\DFF_157/net444 ) );
  and2s1 U3544 ( .Q(g5656), .DIN1(g632), .DIN2(n2828) );
  hi1s1 U3545 ( .Q(n2828), .DIN(g4894) );
  nor2s1 U3546 ( .Q(g5655), .DIN1(g4894), .DIN2(\DFF_136/net423 ) );
  nor2s1 U3547 ( .Q(g5654), .DIN1(g4894), .DIN2(\DFF_336/net623 ) );
  nor2s1 U3548 ( .Q(g5287), .DIN1(g1696), .DIN2(g4901) );
  nor2s1 U3549 ( .Q(g4907), .DIN1(g4217), .DIN2(g1707) );
  nnd2s1 U3550 ( .Q(g4901), .DIN1(g1700), .DIN2(\DFF_275/net562 ) );
  and4s1 U3551 ( .Q(g4897), .DIN1(g928), .DIN2(g932), .DIN3(g936), .DIN4(g940)
         );
  nnd2s1 U3552 ( .Q(g4895), .DIN1(n2895), .DIN2(n2896) );
  nnd2s1 U3553 ( .Q(n2896), .DIN1(n2653), .DIN2(g2639) );
  nnd2s1 U3554 ( .Q(n2895), .DIN1(g754), .DIN2(g2791) );
  nnd2s1 U3555 ( .Q(g4894), .DIN1(n2134), .DIN2(n2897) );
  nnd2s1 U3556 ( .Q(n2897), .DIN1(g611), .DIN2(n1951) );
  nnd3s1 U3557 ( .Q(n2134), .DIN1(n1951), .DIN2(n1975), .DIN3(n2330) );
  nor2s1 U3558 ( .Q(n2330), .DIN1(g599), .DIN2(g605) );
  hi1s1 U3559 ( .Q(g4217), .DIN(g1700) );
  nnd2s1 U3560 ( .Q(g3438), .DIN1(n2898), .DIN2(n2899) );
  nnd2s1 U3561 ( .Q(n2899), .DIN1(g1669), .DIN2(n2074) );
  nnd2s1 U3562 ( .Q(n2898), .DIN1(g1687), .DIN2(g1690) );
  nnd2s1 U3563 ( .Q(g3435), .DIN1(n2900), .DIN2(n2901) );
  nnd2s1 U3564 ( .Q(n2901), .DIN1(g1666), .DIN2(n2074) );
  nnd2s1 U3565 ( .Q(n2900), .DIN1(g1684), .DIN2(g1690) );
  nnd2s1 U3566 ( .Q(g3431), .DIN1(n2902), .DIN2(n2903) );
  nnd2s1 U3567 ( .Q(n2903), .DIN1(g1663), .DIN2(n2074) );
  nnd2s1 U3568 ( .Q(n2902), .DIN1(g1681), .DIN2(g1690) );
  nnd2s1 U3569 ( .Q(g3425), .DIN1(n2904), .DIN2(n2905) );
  nnd2s1 U3570 ( .Q(n2905), .DIN1(g1660), .DIN2(n2074) );
  nnd2s1 U3571 ( .Q(n2904), .DIN1(g1678), .DIN2(g1690) );
  and3s1 U3572 ( .Q(g3418), .DIN1(g743), .DIN2(g109), .DIN3(g744) );
  nnd2s1 U3573 ( .Q(g3414), .DIN1(n2906), .DIN2(n2907) );
  nnd2s1 U3574 ( .Q(n2907), .DIN1(g1657), .DIN2(n2074) );
  nnd2s1 U3575 ( .Q(n2906), .DIN1(g1675), .DIN2(g1690) );
  and3s1 U3576 ( .Q(g3407), .DIN1(g741), .DIN2(g109), .DIN3(g742) );
  nnd2s1 U3577 ( .Q(g3399), .DIN1(n2908), .DIN2(n2909) );
  nnd2s1 U3578 ( .Q(n2909), .DIN1(g1654), .DIN2(n2074) );
  nnd2s1 U3579 ( .Q(n2908), .DIN1(g1672), .DIN2(g1690) );
  nor2s1 U3580 ( .Q(g3329), .DIN1(g1737), .DIN2(g1610) );
  hi1s1 U3581 ( .Q(g3327), .DIN(g23) );
  and2s1 U3582 ( .Q(g2791), .DIN1(g2639), .DIN2(n2910) );
  nor2s1 U3583 ( .Q(g11657), .DIN1(n2911), .DIN2(n2912) );
  and2s1 U3584 ( .Q(n2911), .DIN1(n2913), .DIN2(n2914) );
  or3s1 U3585 ( .Q(n2914), .DIN1(n2000), .DIN2(g4898), .DIN3(n2915) );
  nnd2s1 U3586 ( .Q(n2913), .DIN1(g1351), .DIN2(n2916) );
  nnd2s1 U3587 ( .Q(n2916), .DIN1(g4898), .DIN2(g11593) );
  and4s1 U3588 ( .Q(g4898), .DIN1(g1351), .DIN2(g1346), .DIN3(g1341), .DIN4(
        g1336) );
  nor2s1 U3589 ( .Q(g11656), .DIN1(n2917), .DIN2(n2912) );
  xor2s1 U3590 ( .Q(n2917), .DIN1(g1346), .DIN2(n2915) );
  nnd2s1 U3591 ( .Q(n2915), .DIN1(n2918), .DIN2(g1341) );
  hi1s1 U3592 ( .Q(n2918), .DIN(n2919) );
  nor2s1 U3593 ( .Q(g11655), .DIN1(n2920), .DIN2(n2912) );
  xor2s1 U3594 ( .Q(n2920), .DIN1(n2919), .DIN2(g1341) );
  nnd2s1 U3595 ( .Q(n2919), .DIN1(g11593), .DIN2(g1336) );
  nor2s1 U3596 ( .Q(g11654), .DIN1(n2921), .DIN2(n2912) );
  nnd2s1 U3597 ( .Q(n2912), .DIN1(g109), .DIN2(n2922) );
  nnd3s1 U3598 ( .Q(n2922), .DIN1(n2923), .DIN2(n2011), .DIN3(g1212) );
  xor2s1 U3599 ( .Q(n2921), .DIN1(g1336), .DIN2(n2924) );
  nnd2s1 U3600 ( .Q(g11653), .DIN1(n2925), .DIN2(n2926) );
  nnd2s1 U3601 ( .Q(n2926), .DIN1(g336), .DIN2(n2652) );
  nnd2s1 U3602 ( .Q(n2925), .DIN1(n2927), .DIN2(n2653) );
  nnd2s1 U3603 ( .Q(n2927), .DIN1(n2928), .DIN2(n2929) );
  nnd2s1 U3604 ( .Q(n2929), .DIN1(n2930), .DIN2(n2931) );
  nnd2s1 U3605 ( .Q(n2928), .DIN1(n2932), .DIN2(n2933) );
  nnd2s1 U3606 ( .Q(g11642), .DIN1(n2934), .DIN2(n2935) );
  nnd2s1 U3607 ( .Q(n2935), .DIN1(g345), .DIN2(n2652) );
  nnd2s1 U3608 ( .Q(n2934), .DIN1(n2936), .DIN2(n2653) );
  xor2s1 U3609 ( .Q(n2936), .DIN1(n2933), .DIN2(n2930) );
  xor2s1 U3610 ( .Q(n2930), .DIN1(n2937), .DIN2(n2938) );
  xor2s1 U3611 ( .Q(n2937), .DIN1(n2939), .DIN2(n2940) );
  xor2s1 U3612 ( .Q(n2940), .DIN1(n2941), .DIN2(n2942) );
  xor2s1 U3613 ( .Q(n2942), .DIN1(n2943), .DIN2(n2944) );
  xor2s1 U3614 ( .Q(n2941), .DIN1(n2945), .DIN2(n2946) );
  xor2s1 U3615 ( .Q(n2939), .DIN1(n2947), .DIN2(n2948) );
  xor2s1 U3616 ( .Q(n2948), .DIN1(n2949), .DIN2(n2950) );
  xor2s1 U3617 ( .Q(n2947), .DIN1(n2951), .DIN2(n2952) );
  and2s1 U3618 ( .Q(n2933), .DIN1(n2953), .DIN2(n2954) );
  or2s1 U3619 ( .Q(n2954), .DIN1(n2955), .DIN2(n2077) );
  xor2s1 U3620 ( .Q(n2955), .DIN1(n2956), .DIN2(n2957) );
  nnd4s1 U3621 ( .Q(n2957), .DIN1(g456), .DIN2(n1930), .DIN3(n1977), .DIN4(
        n1950) );
  nnd2s1 U3622 ( .Q(n2953), .DIN1(g305), .DIN2(n2078) );
  nnd2s1 U3623 ( .Q(g11635), .DIN1(n2958), .DIN2(n2959) );
  nnd2s1 U3624 ( .Q(n2959), .DIN1(g1333), .DIN2(n2960) );
  nnd2s1 U3625 ( .Q(n2958), .DIN1(n2961), .DIN2(g1806) );
  nnd2s1 U3626 ( .Q(g11634), .DIN1(n2962), .DIN2(n2963) );
  nnd2s1 U3627 ( .Q(n2963), .DIN1(g1330), .DIN2(n2960) );
  nnd2s1 U3628 ( .Q(n2962), .DIN1(n2961), .DIN2(g1801) );
  nnd2s1 U3629 ( .Q(g11633), .DIN1(n2964), .DIN2(n2965) );
  nnd2s1 U3630 ( .Q(n2965), .DIN1(g1327), .DIN2(n2960) );
  nnd2s1 U3631 ( .Q(n2964), .DIN1(n2961), .DIN2(g1796) );
  nnd2s1 U3632 ( .Q(g11632), .DIN1(n2966), .DIN2(n2967) );
  nnd2s1 U3633 ( .Q(n2967), .DIN1(g1324), .DIN2(n2960) );
  nnd2s1 U3634 ( .Q(n2966), .DIN1(n2961), .DIN2(g1791) );
  nnd2s1 U3635 ( .Q(g11631), .DIN1(n2968), .DIN2(n2969) );
  nnd2s1 U3636 ( .Q(n2969), .DIN1(g1321), .DIN2(n2960) );
  nnd2s1 U3637 ( .Q(n2968), .DIN1(n2961), .DIN2(g1786) );
  nnd2s1 U3638 ( .Q(g11630), .DIN1(n2970), .DIN2(n2971) );
  nnd2s1 U3639 ( .Q(n2971), .DIN1(g1318), .DIN2(n2960) );
  nnd2s1 U3640 ( .Q(n2970), .DIN1(n2961), .DIN2(g1781) );
  nnd2s1 U3641 ( .Q(g11629), .DIN1(n2972), .DIN2(n2973) );
  nnd2s1 U3642 ( .Q(n2973), .DIN1(g1314), .DIN2(n2960) );
  nnd2s1 U3643 ( .Q(n2972), .DIN1(n2961), .DIN2(g1776) );
  nnd2s1 U3644 ( .Q(g11628), .DIN1(n2974), .DIN2(n2975) );
  nnd2s1 U3645 ( .Q(n2975), .DIN1(g1311), .DIN2(n2960) );
  nnd2s1 U3646 ( .Q(n2974), .DIN1(n2961), .DIN2(g1771) );
  nnd2s1 U3647 ( .Q(g11627), .DIN1(n2976), .DIN2(n2977) );
  nnd2s1 U3648 ( .Q(n2977), .DIN1(g1308), .DIN2(n2960) );
  nnd2s1 U3649 ( .Q(n2976), .DIN1(n2961), .DIN2(g1766) );
  hi1s1 U3650 ( .Q(n2961), .DIN(n2960) );
  nnd2s1 U3651 ( .Q(n2960), .DIN1(g1317), .DIN2(g11593) );
  nnd2s1 U3652 ( .Q(g11611), .DIN1(n2978), .DIN2(n2979) );
  nnd2s1 U3653 ( .Q(n2979), .DIN1(g1618), .DIN2(n2070) );
  nnd2s1 U3654 ( .Q(n2978), .DIN1(n2980), .DIN2(n2063) );
  xor2s1 U3655 ( .Q(n2980), .DIN1(n2981), .DIN2(n2982) );
  xor2s1 U3656 ( .Q(n2982), .DIN1(g1610), .DIN2(n2983) );
  nnd2s1 U3657 ( .Q(n2983), .DIN1(n2984), .DIN2(n2985) );
  nnd2s1 U3658 ( .Q(n2985), .DIN1(n2986), .DIN2(n2987) );
  nnd2s1 U3659 ( .Q(n2986), .DIN1(n2988), .DIN2(n2989) );
  or2s1 U3660 ( .Q(n2989), .DIN1(n2990), .DIN2(g1149) );
  nnd2s1 U3661 ( .Q(n2988), .DIN1(g1153), .DIN2(g1149) );
  nnd2s1 U3662 ( .Q(n2984), .DIN1(n2991), .DIN2(n2992) );
  nnd2s1 U3663 ( .Q(n2992), .DIN1(n2993), .DIN2(n2994) );
  nnd2s1 U3664 ( .Q(n2994), .DIN1(g1149), .DIN2(n1988) );
  nnd2s1 U3665 ( .Q(n2993), .DIN1(n2990), .DIN2(n2016) );
  nnd2s1 U3666 ( .Q(n2990), .DIN1(n1988), .DIN2(n2995) );
  or4s1 U3667 ( .Q(n2995), .DIN1(n2996), .DIN2(n2997), .DIN3(n2998), .DIN4(
        n2999) );
  nnd3s1 U3668 ( .Q(n2999), .DIN1(n1944), .DIN2(n1970), .DIN3(n2013) );
  nnd4s1 U3669 ( .Q(n2998), .DIN1(n2005), .DIN2(n1966), .DIN3(n1942), .DIN4(
        n1927) );
  nnd3s1 U3670 ( .Q(n2997), .DIN1(n1969), .DIN2(n2015), .DIN3(n1934) );
  nnd3s1 U3671 ( .Q(n2996), .DIN1(n1945), .DIN2(n1971), .DIN3(n2014) );
  hi1s1 U3672 ( .Q(n2991), .DIN(n2987) );
  nnd4s1 U3673 ( .Q(n2987), .DIN1(g1101), .DIN2(n1976), .DIN3(n1929), .DIN4(
        n1949) );
  nor2s1 U3674 ( .Q(g11594), .DIN1(n3000), .DIN2(n2065) );
  xor2s1 U3675 ( .Q(n3000), .DIN1(n3001), .DIN2(n3002) );
  xor2s1 U3676 ( .Q(n3002), .DIN1(g1415), .DIN2(n2981) );
  and2s1 U3677 ( .Q(n2981), .DIN1(n3003), .DIN2(n3004) );
  nnd2s1 U3678 ( .Q(n3004), .DIN1(n3005), .DIN2(n2072) );
  nnd2s1 U3679 ( .Q(n3005), .DIN1(n3006), .DIN2(n3007) );
  or2s1 U3680 ( .Q(n3007), .DIN1(n3008), .DIN2(g1811) );
  nnd2s1 U3681 ( .Q(n3006), .DIN1(n3009), .DIN2(n3008) );
  nnd4s1 U3682 ( .Q(n3008), .DIN1(n2006), .DIN2(n1967), .DIN3(n1943), .DIN4(
        n1928) );
  nnd2s1 U3683 ( .Q(n3009), .DIN1(n3010), .DIN2(n3011) );
  nnd2s1 U3684 ( .Q(n3003), .DIN1(g201), .DIN2(g18) );
  xor2s1 U3685 ( .Q(n3001), .DIN1(g1419), .DIN2(n3012) );
  xor2s1 U3686 ( .Q(n3012), .DIN1(g1515), .DIN2(g1448) );
  hi1s1 U3687 ( .Q(g11593), .DIN(n2924) );
  nnd3s1 U3688 ( .Q(n2924), .DIN1(n2799), .DIN2(n3013), .DIN3(n2544) );
  or4s1 U3689 ( .Q(n3013), .DIN1(n3014), .DIN2(n3015), .DIN3(n3016), .DIN4(
        n3017) );
  nnd4s1 U3690 ( .Q(n3017), .DIN1(n3018), .DIN2(n3019), .DIN3(n3020), .DIN4(
        n3021) );
  nor2s1 U3691 ( .Q(n3021), .DIN1(n3022), .DIN2(n3023) );
  xor2s1 U3692 ( .Q(n3023), .DIN1(g1265), .DIN2(g1015) );
  xor2s1 U3693 ( .Q(n3022), .DIN1(g1250), .DIN2(g1011) );
  hi1s1 U3694 ( .Q(n3020), .DIN(n3024) );
  xor2s1 U3695 ( .Q(n3024), .DIN1(g1240), .DIN2(g1003) );
  hi1s1 U3696 ( .Q(n3019), .DIN(n3025) );
  xor2s1 U3697 ( .Q(n3025), .DIN1(g1255), .DIN2(g1007) );
  xor2s1 U3698 ( .Q(n3018), .DIN1(n3026), .DIN2(n3027) );
  or3s1 U3699 ( .Q(n3016), .DIN1(n3028), .DIN2(n3029), .DIN3(n3030) );
  xor2s1 U3700 ( .Q(n3030), .DIN1(g1270), .DIN2(g1023) );
  xor2s1 U3701 ( .Q(n3029), .DIN1(g1235), .DIN2(g991) );
  xor2s1 U3702 ( .Q(n3028), .DIN1(g1260), .DIN2(g1019) );
  xor2s1 U3703 ( .Q(n3015), .DIN1(g995), .DIN2(g1275) );
  xor2s1 U3704 ( .Q(n3014), .DIN1(g999), .DIN2(g1245) );
  nnd2s1 U3705 ( .Q(g11513), .DIN1(n3031), .DIN2(n3032) );
  nnd2s1 U3706 ( .Q(n3032), .DIN1(g342), .DIN2(n2652) );
  nnd2s1 U3707 ( .Q(n3031), .DIN1(n2943), .DIN2(n2653) );
  nnd2s1 U3708 ( .Q(n2943), .DIN1(n3033), .DIN2(n3034) );
  nnd2s1 U3709 ( .Q(n3034), .DIN1(n3035), .DIN2(n2071) );
  xor2s1 U3710 ( .Q(n3035), .DIN1(g516), .DIN2(n3037) );
  nor2s1 U3711 ( .Q(n3037), .DIN1(n2073), .DIN2(n3038) );
  nnd2s1 U3712 ( .Q(n3033), .DIN1(g309), .DIN2(n2079) );
  nnd2s1 U3713 ( .Q(g11512), .DIN1(n3039), .DIN2(n3040) );
  nnd2s1 U3714 ( .Q(n3040), .DIN1(g366), .DIN2(n2652) );
  nnd2s1 U3715 ( .Q(n3039), .DIN1(n2944), .DIN2(n2653) );
  nnd2s1 U3716 ( .Q(n2944), .DIN1(n3041), .DIN2(n3042) );
  nnd2s1 U3717 ( .Q(n3042), .DIN1(n3043), .DIN2(n3036) );
  xor2s1 U3718 ( .Q(n3043), .DIN1(g511), .DIN2(n3044) );
  nor2s1 U3719 ( .Q(n3044), .DIN1(g456), .DIN2(n3038) );
  nnd3s1 U3720 ( .Q(n3038), .DIN1(n1930), .DIN2(n1977), .DIN3(g471) );
  nnd2s1 U3721 ( .Q(n3041), .DIN1(g333), .DIN2(n2078) );
  nnd2s1 U3722 ( .Q(g11511), .DIN1(n3045), .DIN2(n3046) );
  nnd2s1 U3723 ( .Q(n3046), .DIN1(g363), .DIN2(n2652) );
  nnd2s1 U3724 ( .Q(n3045), .DIN1(n2945), .DIN2(n2653) );
  nnd2s1 U3725 ( .Q(n2945), .DIN1(n3047), .DIN2(n3048) );
  nnd2s1 U3726 ( .Q(n3048), .DIN1(n3049), .DIN2(n2071) );
  xor2s1 U3727 ( .Q(n3049), .DIN1(g506), .DIN2(n3050) );
  nor2s1 U3728 ( .Q(n3050), .DIN1(g471), .DIN2(n3051) );
  nnd2s1 U3729 ( .Q(n3047), .DIN1(g330), .DIN2(n2079) );
  nnd2s1 U3730 ( .Q(g11510), .DIN1(n3052), .DIN2(n3053) );
  nnd2s1 U3731 ( .Q(n3053), .DIN1(g360), .DIN2(n2652) );
  nnd2s1 U3732 ( .Q(n3052), .DIN1(n2946), .DIN2(n2653) );
  nnd2s1 U3733 ( .Q(n2946), .DIN1(n3054), .DIN2(n3055) );
  or2s1 U3734 ( .Q(n3055), .DIN1(n3056), .DIN2(n2078) );
  xor2s1 U3735 ( .Q(n3056), .DIN1(n3057), .DIN2(g501) );
  nnd3s1 U3736 ( .Q(n3057), .DIN1(n3058), .DIN2(n1950), .DIN3(g466) );
  nnd2s1 U3737 ( .Q(n3054), .DIN1(g327), .DIN2(n2078) );
  nnd2s1 U3738 ( .Q(g11509), .DIN1(n3059), .DIN2(n3060) );
  nnd2s1 U3739 ( .Q(n3060), .DIN1(g357), .DIN2(n2652) );
  nnd2s1 U3740 ( .Q(n3059), .DIN1(n2949), .DIN2(n2653) );
  nnd2s1 U3741 ( .Q(n2949), .DIN1(n3061), .DIN2(n3062) );
  nnd2s1 U3742 ( .Q(n3062), .DIN1(n3063), .DIN2(n3036) );
  xor2s1 U3743 ( .Q(n3063), .DIN1(g496), .DIN2(n3064) );
  nor2s1 U3744 ( .Q(n3064), .DIN1(n2073), .DIN2(n3065) );
  nnd2s1 U3745 ( .Q(n3061), .DIN1(g324), .DIN2(n2077) );
  nnd2s1 U3746 ( .Q(g11508), .DIN1(n3066), .DIN2(n3067) );
  nnd2s1 U3747 ( .Q(n3067), .DIN1(g354), .DIN2(n2652) );
  nnd2s1 U3748 ( .Q(n3066), .DIN1(n2950), .DIN2(n2653) );
  nnd2s1 U3749 ( .Q(n2950), .DIN1(n3068), .DIN2(n3069) );
  nnd2s1 U3750 ( .Q(n3069), .DIN1(n3070), .DIN2(n2076) );
  xor2s1 U3751 ( .Q(n3070), .DIN1(g491), .DIN2(n3071) );
  nor2s1 U3752 ( .Q(n3071), .DIN1(g456), .DIN2(n3065) );
  nnd3s1 U3753 ( .Q(n3065), .DIN1(n1930), .DIN2(n1950), .DIN3(g466) );
  nnd2s1 U3754 ( .Q(n3068), .DIN1(g321), .DIN2(n2079) );
  nnd2s1 U3755 ( .Q(g11507), .DIN1(n3072), .DIN2(n3073) );
  nnd2s1 U3756 ( .Q(n3073), .DIN1(g351), .DIN2(n2652) );
  nnd2s1 U3757 ( .Q(n3072), .DIN1(n2951), .DIN2(n2653) );
  nnd2s1 U3758 ( .Q(n2951), .DIN1(n3074), .DIN2(n3075) );
  nnd2s1 U3759 ( .Q(n3075), .DIN1(n3076), .DIN2(n2071) );
  xor2s1 U3760 ( .Q(n3076), .DIN1(g486), .DIN2(n3077) );
  nor2s1 U3761 ( .Q(n3077), .DIN1(n2073), .DIN2(n3078) );
  nnd2s1 U3762 ( .Q(n3074), .DIN1(g318), .DIN2(n2077) );
  nnd2s1 U3763 ( .Q(g11506), .DIN1(n3079), .DIN2(n3080) );
  nnd2s1 U3764 ( .Q(n3080), .DIN1(g348), .DIN2(n2652) );
  nnd2s1 U3765 ( .Q(n3079), .DIN1(n2952), .DIN2(n2653) );
  nnd2s1 U3766 ( .Q(n2952), .DIN1(n3081), .DIN2(n3082) );
  nnd2s1 U3767 ( .Q(n3082), .DIN1(n3083), .DIN2(n2071) );
  xor2s1 U3768 ( .Q(n3083), .DIN1(g481), .DIN2(n3084) );
  nor2s1 U3769 ( .Q(n3084), .DIN1(g456), .DIN2(n3078) );
  nnd3s1 U3770 ( .Q(n3078), .DIN1(n1977), .DIN2(n1950), .DIN3(g461) );
  nnd2s1 U3771 ( .Q(n3081), .DIN1(g315), .DIN2(n2078) );
  nnd2s1 U3772 ( .Q(g11505), .DIN1(n3085), .DIN2(n3086) );
  nnd2s1 U3773 ( .Q(n3086), .DIN1(g339), .DIN2(n2652) );
  hi1s1 U3774 ( .Q(n2652), .DIN(n2653) );
  nnd2s1 U3775 ( .Q(n3085), .DIN1(n2938), .DIN2(n2653) );
  nor2s1 U3776 ( .Q(n2653), .DIN1(n2910), .DIN2(g754) );
  hi1s1 U3777 ( .Q(n2910), .DIN(g750) );
  nnd2s1 U3778 ( .Q(n2938), .DIN1(n3087), .DIN2(n3088) );
  or2s1 U3779 ( .Q(n3088), .DIN1(n3089), .DIN2(n2077) );
  xor2s1 U3780 ( .Q(n3089), .DIN1(n3090), .DIN2(g476) );
  nnd3s1 U3781 ( .Q(n3090), .DIN1(n3058), .DIN2(n1977), .DIN3(g471) );
  nnd2s1 U3782 ( .Q(n3087), .DIN1(g312), .DIN2(n2077) );
  nor2s1 U3783 ( .Q(g11473), .DIN1(n3091), .DIN2(n3092) );
  and2s1 U3784 ( .Q(n3092), .DIN1(n3093), .DIN2(n3094) );
  nnd3s1 U3785 ( .Q(n3094), .DIN1(g981), .DIN2(n3095), .DIN3(n3096) );
  nnd2s1 U3786 ( .Q(n3093), .DIN1(g986), .DIN2(n3097) );
  nnd2s1 U3787 ( .Q(n3097), .DIN1(g4896), .DIN2(g11179) );
  hi1s1 U3788 ( .Q(g4896), .DIN(n3095) );
  nnd4s1 U3789 ( .Q(n3095), .DIN1(g986), .DIN2(g981), .DIN3(g976), .DIN4(g971)
         );
  nor2s1 U3790 ( .Q(g11472), .DIN1(n3098), .DIN2(n3091) );
  hi1s1 U3791 ( .Q(n3098), .DIN(n3099) );
  xor2s1 U3792 ( .Q(n3099), .DIN1(g981), .DIN2(n3096) );
  nor2s1 U3793 ( .Q(n3096), .DIN1(n3100), .DIN2(n2044) );
  nor2s1 U3794 ( .Q(g11471), .DIN1(n3101), .DIN2(n3091) );
  xor2s1 U3795 ( .Q(n3101), .DIN1(g976), .DIN2(n3100) );
  nnd2s1 U3796 ( .Q(n3100), .DIN1(g11179), .DIN2(g971) );
  nor2s1 U3797 ( .Q(g11470), .DIN1(n3102), .DIN2(n3091) );
  nnd2s1 U3798 ( .Q(n3091), .DIN1(g109), .DIN2(n3103) );
  nnd3s1 U3799 ( .Q(n3103), .DIN1(n3104), .DIN2(n3105), .DIN3(g869) );
  xor2s1 U3800 ( .Q(n3102), .DIN1(g971), .DIN2(n3106) );
  nor2s1 U3801 ( .Q(g11469), .DIN1(n3107), .DIN2(n3108) );
  nor2s1 U3802 ( .Q(n3107), .DIN1(n3109), .DIN2(g471) );
  nor2s1 U3803 ( .Q(n3109), .DIN1(n3051), .DIN2(n3110) );
  and2s1 U3804 ( .Q(g11468), .DIN1(n3111), .DIN2(n3112) );
  nnd2s1 U3805 ( .Q(n3112), .DIN1(n3113), .DIN2(n3114) );
  nnd4s1 U3806 ( .Q(n3114), .DIN1(n3115), .DIN2(g461), .DIN3(g456), .DIN4(
        n3051) );
  nnd2s1 U3807 ( .Q(n3113), .DIN1(g466), .DIN2(n3116) );
  nnd2s1 U3808 ( .Q(n3116), .DIN1(n3115), .DIN2(n3117) );
  and2s1 U3809 ( .Q(g11467), .DIN1(n3111), .DIN2(n3118) );
  nnd3s1 U3810 ( .Q(n3118), .DIN1(n3119), .DIN2(n3120), .DIN3(n3121) );
  hi1s1 U3811 ( .Q(n3121), .DIN(n3058) );
  nor2s1 U3812 ( .Q(n3058), .DIN1(n1930), .DIN2(g456) );
  nnd2s1 U3813 ( .Q(n3120), .DIN1(g461), .DIN2(n3110) );
  nnd3s1 U3814 ( .Q(n3119), .DIN1(g456), .DIN2(n1930), .DIN3(n3115) );
  hi1s1 U3815 ( .Q(n3111), .DIN(n3108) );
  nor2s1 U3816 ( .Q(g11466), .DIN1(n3122), .DIN2(n3108) );
  nnd2s1 U3817 ( .Q(n3108), .DIN1(g109), .DIN2(\DFF_441/net728 ) );
  xor2s1 U3818 ( .Q(n3122), .DIN1(n2073), .DIN2(n3115) );
  hi1s1 U3819 ( .Q(n3115), .DIN(n3110) );
  nnd2s1 U3820 ( .Q(n3110), .DIN1(n3036), .DIN2(n3123) );
  nnd2s1 U3821 ( .Q(n3123), .DIN1(n3117), .DIN2(g471) );
  hi1s1 U3822 ( .Q(n3117), .DIN(n3051) );
  nnd3s1 U3823 ( .Q(n3051), .DIN1(g461), .DIN2(g456), .DIN3(g466) );
  nnd2s1 U3824 ( .Q(g11443), .DIN1(n3124), .DIN2(n3125) );
  nnd2s1 U3825 ( .Q(n3125), .DIN1(g1275), .DIN2(n2060) );
  nnd2s1 U3826 ( .Q(n3124), .DIN1(n2799), .DIN2(n3027) );
  nnd2s1 U3827 ( .Q(n3027), .DIN1(n3126), .DIN2(n3127) );
  or2s1 U3828 ( .Q(n3127), .DIN1(n3026), .DIN2(n2544) );
  xor2s1 U3829 ( .Q(n3026), .DIN1(g1027), .DIN2(n3128) );
  nnd2s1 U3830 ( .Q(n3128), .DIN1(g1032), .DIN2(n2931) );
  nnd2s1 U3831 ( .Q(n3126), .DIN1(n3129), .DIN2(n2544) );
  nor2s1 U3832 ( .Q(n2544), .DIN1(n2048), .DIN2(n2535) );
  nnd3s1 U3833 ( .Q(n2535), .DIN1(g1223), .DIN2(g1218), .DIN3(g1227) );
  nnd2s1 U3834 ( .Q(n3129), .DIN1(n3130), .DIN2(n3131) );
  nnd2s1 U3835 ( .Q(n3131), .DIN1(g1280), .DIN2(n2031) );
  nnd2s1 U3836 ( .Q(n3130), .DIN1(n3132), .DIN2(n2052) );
  nnd2s1 U3837 ( .Q(n3132), .DIN1(n2031), .DIN2(n3133) );
  or4s1 U3838 ( .Q(n3133), .DIN1(n3134), .DIN2(n3135), .DIN3(n3136), .DIN4(
        n3137) );
  or3s1 U3839 ( .Q(n3137), .DIN1(g1270), .DIN2(g1275), .DIN3(g1265) );
  or4s1 U3840 ( .Q(n3136), .DIN1(g1292), .DIN2(g1296), .DIN3(g1300), .DIN4(
        g1304) );
  or3s1 U3841 ( .Q(n3135), .DIN1(g1240), .DIN2(g1245), .DIN3(g1235) );
  or3s1 U3842 ( .Q(n3134), .DIN1(g1255), .DIN2(g1260), .DIN3(g1250) );
  hi1s1 U3843 ( .Q(n2799), .DIN(n2543) );
  nnd3s1 U3844 ( .Q(n2543), .DIN1(n2063), .DIN2(n2061), .DIN3(g1289) );
  nor2s1 U3845 ( .Q(g11442), .DIN1(n3138), .DIN2(n3139) );
  nor2s1 U3846 ( .Q(n3138), .DIN1(n3140), .DIN2(g382) );
  nor2s1 U3847 ( .Q(n3140), .DIN1(n3141), .DIN2(n3142) );
  and2s1 U3848 ( .Q(g11441), .DIN1(n3143), .DIN2(n3144) );
  nnd2s1 U3849 ( .Q(n3144), .DIN1(n3145), .DIN2(n3146) );
  nnd4s1 U3850 ( .Q(n3146), .DIN1(n3147), .DIN2(g374), .DIN3(g369), .DIN4(
        n3141) );
  nnd2s1 U3851 ( .Q(n3145), .DIN1(g378), .DIN2(n3148) );
  nnd2s1 U3852 ( .Q(n3148), .DIN1(n3147), .DIN2(n3149) );
  and2s1 U3853 ( .Q(g11440), .DIN1(n3150), .DIN2(n3143) );
  xor2s1 U3854 ( .Q(n3150), .DIN1(n3151), .DIN2(g374) );
  and2s1 U3855 ( .Q(n3151), .DIN1(g369), .DIN2(n3147) );
  nor2s1 U3856 ( .Q(g11439), .DIN1(n3152), .DIN2(n3139) );
  hi1s1 U3857 ( .Q(n3139), .DIN(n3143) );
  nor2s1 U3858 ( .Q(n3143), .DIN1(n2064), .DIN2(g869) );
  xor2s1 U3859 ( .Q(n3152), .DIN1(g369), .DIN2(n3142) );
  hi1s1 U3860 ( .Q(n3142), .DIN(n3147) );
  nor2s1 U3861 ( .Q(n3147), .DIN1(n2078), .DIN2(n3153) );
  nnd3s1 U3862 ( .Q(g11409), .DIN1(n3154), .DIN2(n3155), .DIN3(n3156) );
  nnd3s1 U3863 ( .Q(n3156), .DIN1(n3157), .DIN2(n3158), .DIN3(n2233) );
  nnd3s1 U3864 ( .Q(n3158), .DIN1(n3159), .DIN2(n3160), .DIN3(n2074) );
  nnd2s1 U3865 ( .Q(n3160), .DIN1(n3161), .DIN2(n3162) );
  nnd2s1 U3866 ( .Q(n3162), .DIN1(g1771), .DIN2(g1766) );
  nnd2s1 U3867 ( .Q(n3161), .DIN1(g1781), .DIN2(g1776) );
  nnd2s1 U3868 ( .Q(n3159), .DIN1(n3163), .DIN2(n3164) );
  nnd2s1 U3869 ( .Q(n3164), .DIN1(g1791), .DIN2(g1786) );
  nnd2s1 U3870 ( .Q(n3163), .DIN1(g1801), .DIN2(g1796) );
  nnd3s1 U3871 ( .Q(n3157), .DIN1(n3165), .DIN2(n3166), .DIN3(g1690) );
  nnd2s1 U3872 ( .Q(n3166), .DIN1(n3167), .DIN2(n3168) );
  nnd2s1 U3873 ( .Q(n3168), .DIN1(g10775), .DIN2(g10774) );
  nnd2s1 U3874 ( .Q(n3167), .DIN1(g10871), .DIN2(g10872) );
  nnd2s1 U3875 ( .Q(n3165), .DIN1(n3169), .DIN2(n3170) );
  nnd2s1 U3876 ( .Q(n3170), .DIN1(g10867), .DIN2(g10868) );
  nnd2s1 U3877 ( .Q(n3169), .DIN1(g10869), .DIN2(g10870) );
  nnd3s1 U3878 ( .Q(n3155), .DIN1(n2095), .DIN2(n3171), .DIN3(n1989) );
  nnd3s1 U3879 ( .Q(n3171), .DIN1(n2118), .DIN2(n2119), .DIN3(n2231) );
  hi1s1 U3880 ( .Q(n2231), .DIN(n2113) );
  nnd2s1 U3881 ( .Q(n2113), .DIN1(n2107), .DIN2(n3172) );
  nnd2s1 U3882 ( .Q(n3172), .DIN1(g1822), .DIN2(n1980) );
  hi1s1 U3883 ( .Q(n2118), .DIN(n2239) );
  nnd2s1 U3884 ( .Q(n3154), .DIN1(n2600), .DIN2(g1857) );
  nor2s1 U3885 ( .Q(n2600), .DIN1(n2233), .DIN2(n2095) );
  nor2s1 U3886 ( .Q(n2095), .DIN1(n2602), .DIN2(g1868) );
  nnd2s1 U3887 ( .Q(n2602), .DIN1(n2607), .DIN2(n2027) );
  nor2s1 U3888 ( .Q(n2607), .DIN1(n1998), .DIN2(g1861) );
  nnd2s1 U3889 ( .Q(g11408), .DIN1(n3173), .DIN2(n3174) );
  nnd2s1 U3890 ( .Q(n3174), .DIN1(n3175), .DIN2(n2102) );
  nnd2s1 U3891 ( .Q(n3175), .DIN1(n2107), .DIN2(n3176) );
  nnd2s1 U3892 ( .Q(n3176), .DIN1(g2731), .DIN2(n3177) );
  nnd3s1 U3893 ( .Q(n3177), .DIN1(g5672), .DIN2(n3178), .DIN3(n3179) );
  xor2s1 U3894 ( .Q(n3179), .DIN1(n3180), .DIN2(n3181) );
  nnd2s1 U3895 ( .Q(n3180), .DIN1(n3182), .DIN2(n3183) );
  nnd2s1 U3896 ( .Q(n3183), .DIN1(n2239), .DIN2(g1857) );
  nor2s1 U3897 ( .Q(n2239), .DIN1(n1953), .DIN2(g1814) );
  nnd2s1 U3898 ( .Q(n3182), .DIN1(n3184), .DIN2(n1989) );
  nnd2s1 U3899 ( .Q(n3184), .DIN1(n1948), .DIN2(n2119) );
  nnd2s1 U3900 ( .Q(n2119), .DIN1(g1828), .DIN2(g1814) );
  nnd3s1 U3901 ( .Q(n3178), .DIN1(g1840), .DIN2(n1948), .DIN3(n2238) );
  and2s1 U3902 ( .Q(g5672), .DIN1(g1850), .DIN2(n2707) );
  hi1s1 U3903 ( .Q(n2707), .DIN(g4906) );
  nnd2s1 U3904 ( .Q(g4906), .DIN1(n2102), .DIN2(n3185) );
  nnd2s1 U3905 ( .Q(n3185), .DIN1(g1834), .DIN2(n1986) );
  nnd3s1 U3906 ( .Q(n2107), .DIN1(n1986), .DIN2(n1953), .DIN3(g1828) );
  nnd2s1 U3907 ( .Q(n3173), .DIN1(n3186), .DIN2(n2233) );
  hi1s1 U3908 ( .Q(n2233), .DIN(n2102) );
  nnd3s1 U3909 ( .Q(n2102), .DIN1(n1986), .DIN2(n1948), .DIN3(n2238) );
  nor2s1 U3910 ( .Q(n2238), .DIN1(g1822), .DIN2(g1828) );
  nnd2s1 U3911 ( .Q(n3186), .DIN1(n3187), .DIN2(n3188) );
  or2s1 U3912 ( .Q(n3188), .DIN1(n2075), .DIN2(g1806) );
  nnd2s1 U3913 ( .Q(n3187), .DIN1(g1690), .DIN2(n3189) );
  nnd2s1 U3914 ( .Q(g11406), .DIN1(n3190), .DIN2(n3191) );
  nnd2s1 U3915 ( .Q(n3191), .DIN1(g968), .DIN2(n3192) );
  nnd2s1 U3916 ( .Q(n3190), .DIN1(g861), .DIN2(n3193) );
  nnd2s1 U3917 ( .Q(g11405), .DIN1(n3194), .DIN2(n3195) );
  nnd2s1 U3918 ( .Q(n3195), .DIN1(g965), .DIN2(n3192) );
  nnd2s1 U3919 ( .Q(n3194), .DIN1(g857), .DIN2(n3193) );
  nnd2s1 U3920 ( .Q(g11404), .DIN1(n3196), .DIN2(n3197) );
  nnd2s1 U3921 ( .Q(n3197), .DIN1(g962), .DIN2(n3192) );
  nnd2s1 U3922 ( .Q(n3196), .DIN1(g853), .DIN2(n3193) );
  nnd2s1 U3923 ( .Q(g11403), .DIN1(n3198), .DIN2(n3199) );
  nnd2s1 U3924 ( .Q(n3199), .DIN1(g959), .DIN2(n3192) );
  nnd2s1 U3925 ( .Q(n3198), .DIN1(g849), .DIN2(n3193) );
  nnd2s1 U3926 ( .Q(g11402), .DIN1(n3200), .DIN2(n3201) );
  nnd2s1 U3927 ( .Q(n3201), .DIN1(g956), .DIN2(n3192) );
  nnd2s1 U3928 ( .Q(n3200), .DIN1(g845), .DIN2(n3193) );
  nnd2s1 U3929 ( .Q(g11401), .DIN1(n3202), .DIN2(n3203) );
  nnd2s1 U3930 ( .Q(n3203), .DIN1(g953), .DIN2(n3192) );
  nnd2s1 U3931 ( .Q(n3202), .DIN1(g841), .DIN2(n3193) );
  nnd2s1 U3932 ( .Q(g11400), .DIN1(n3204), .DIN2(n3205) );
  nnd2s1 U3933 ( .Q(n3205), .DIN1(g950), .DIN2(n3192) );
  nnd2s1 U3934 ( .Q(n3204), .DIN1(g837), .DIN2(n3193) );
  nnd2s1 U3935 ( .Q(g11399), .DIN1(n3206), .DIN2(n3207) );
  nnd2s1 U3936 ( .Q(n3207), .DIN1(g947), .DIN2(n3192) );
  nnd2s1 U3937 ( .Q(n3206), .DIN1(g833), .DIN2(n3193) );
  nnd2s1 U3938 ( .Q(g11398), .DIN1(n3208), .DIN2(n3209) );
  nnd2s1 U3939 ( .Q(n3209), .DIN1(g944), .DIN2(n3192) );
  nnd2s1 U3940 ( .Q(n3208), .DIN1(g829), .DIN2(n3193) );
  hi1s1 U3941 ( .Q(n3193), .DIN(n3192) );
  nnd3s1 U3942 ( .Q(n3192), .DIN1(n3210), .DIN2(n3105), .DIN3(g11179) );
  or2s1 U3943 ( .Q(n3210), .DIN1(n3104), .DIN2(n2066) );
  hi1s1 U3944 ( .Q(g11397), .DIN(n3211) );
  nnd2s1 U3945 ( .Q(g11338), .DIN1(n3212), .DIN2(n3213) );
  nnd2s1 U3946 ( .Q(n3213), .DIN1(g516), .DIN2(n2071) );
  nnd2s1 U3947 ( .Q(n3212), .DIN1(g476), .DIN2(n2078) );
  nnd2s1 U3948 ( .Q(g11337), .DIN1(n3214), .DIN2(n3215) );
  nnd2s1 U3949 ( .Q(n3215), .DIN1(g511), .DIN2(n3036) );
  nnd2s1 U3950 ( .Q(n3214), .DIN1(g516), .DIN2(n2079) );
  nnd2s1 U3951 ( .Q(g11336), .DIN1(n3216), .DIN2(n3217) );
  nnd2s1 U3952 ( .Q(n3217), .DIN1(g506), .DIN2(n2076) );
  nnd2s1 U3953 ( .Q(n3216), .DIN1(g511), .DIN2(n2077) );
  nnd2s1 U3954 ( .Q(g11335), .DIN1(n3218), .DIN2(n3219) );
  nnd2s1 U3955 ( .Q(n3219), .DIN1(g501), .DIN2(n2071) );
  nnd2s1 U3956 ( .Q(n3218), .DIN1(g506), .DIN2(n2078) );
  nnd2s1 U3957 ( .Q(g11334), .DIN1(n3220), .DIN2(n3221) );
  nnd2s1 U3958 ( .Q(n3221), .DIN1(g496), .DIN2(n3036) );
  nnd2s1 U3959 ( .Q(n3220), .DIN1(g501), .DIN2(n2079) );
  nnd2s1 U3960 ( .Q(g11333), .DIN1(n3222), .DIN2(n3223) );
  nnd2s1 U3961 ( .Q(n3223), .DIN1(g491), .DIN2(n2071) );
  nnd2s1 U3962 ( .Q(n3222), .DIN1(g496), .DIN2(n2079) );
  nnd2s1 U3963 ( .Q(g11332), .DIN1(n3224), .DIN2(n3225) );
  nnd2s1 U3964 ( .Q(n3225), .DIN1(g486), .DIN2(n3036) );
  nnd2s1 U3965 ( .Q(n3224), .DIN1(g491), .DIN2(n2077) );
  nnd2s1 U3966 ( .Q(g11331), .DIN1(n3226), .DIN2(n3227) );
  nnd2s1 U3967 ( .Q(n3227), .DIN1(g481), .DIN2(n3036) );
  nnd2s1 U3968 ( .Q(n3226), .DIN1(g486), .DIN2(n2077) );
  nnd2s1 U3969 ( .Q(g11330), .DIN1(n3228), .DIN2(n3229) );
  nnd2s1 U3970 ( .Q(n3229), .DIN1(g525), .DIN2(n2076) );
  nnd2s1 U3971 ( .Q(n3228), .DIN1(g521), .DIN2(n2078) );
  nnd2s1 U3972 ( .Q(g11329), .DIN1(n3230), .DIN2(n3231) );
  nnd2s1 U3973 ( .Q(n3231), .DIN1(g530), .DIN2(n2071) );
  nnd2s1 U3974 ( .Q(n3230), .DIN1(n2077), .DIN2(g525) );
  nnd2s1 U3975 ( .Q(g11328), .DIN1(n3232), .DIN2(n3233) );
  nnd2s1 U3976 ( .Q(n3233), .DIN1(g534), .DIN2(n3036) );
  nnd2s1 U3977 ( .Q(n3232), .DIN1(g530), .DIN2(n2078) );
  nnd2s1 U3978 ( .Q(g11327), .DIN1(n3234), .DIN2(n3235) );
  nnd2s1 U3979 ( .Q(n3235), .DIN1(g538), .DIN2(n2076) );
  nnd2s1 U3980 ( .Q(n3234), .DIN1(g534), .DIN2(n2078) );
  nnd2s1 U3981 ( .Q(g11326), .DIN1(n3236), .DIN2(n3237) );
  nnd2s1 U3982 ( .Q(n3237), .DIN1(g542), .DIN2(n2071) );
  nnd2s1 U3983 ( .Q(n3236), .DIN1(g538), .DIN2(n2077) );
  nnd2s1 U3984 ( .Q(g11325), .DIN1(n3238), .DIN2(n3239) );
  nnd2s1 U3985 ( .Q(n3239), .DIN1(g476), .DIN2(n2071) );
  nnd2s1 U3986 ( .Q(n3238), .DIN1(g542), .DIN2(n2078) );
  nnd2s1 U3987 ( .Q(g11324), .DIN1(n3240), .DIN2(n3241) );
  nnd2s1 U3988 ( .Q(n3241), .DIN1(n2956), .DIN2(n2076) );
  nnd2s1 U3989 ( .Q(n2956), .DIN1(n3242), .DIN2(n3243) );
  nnd2s1 U3990 ( .Q(n3243), .DIN1(g521), .DIN2(n2032) );
  nnd2s1 U3991 ( .Q(n3242), .DIN1(n3244), .DIN2(n2053) );
  nnd2s1 U3992 ( .Q(n3244), .DIN1(n2032), .DIN2(n3245) );
  or4s1 U3993 ( .Q(n3245), .DIN1(n3246), .DIN2(n3247), .DIN3(n3248), .DIN4(
        n3249) );
  or3s1 U3994 ( .Q(n3249), .DIN1(g511), .DIN2(g516), .DIN3(g506) );
  or4s1 U3995 ( .Q(n3248), .DIN1(g530), .DIN2(g534), .DIN3(g538), .DIN4(g542)
         );
  or3s1 U3996 ( .Q(n3247), .DIN1(g481), .DIN2(g486), .DIN3(g476) );
  or3s1 U3997 ( .Q(n3246), .DIN1(g496), .DIN2(g501), .DIN3(g491) );
  nnd2s1 U3998 ( .Q(n3240), .DIN1(g481), .DIN2(n2079) );
  nnd2s1 U3999 ( .Q(g11270), .DIN1(n3250), .DIN2(n3251) );
  nnd2s1 U4000 ( .Q(n3251), .DIN1(g416), .DIN2(n2071) );
  nnd2s1 U4001 ( .Q(n3250), .DIN1(g421), .DIN2(n2077) );
  nnd2s1 U4002 ( .Q(g11269), .DIN1(n3252), .DIN2(n3253) );
  nnd2s1 U4003 ( .Q(n3253), .DIN1(g411), .DIN2(n2071) );
  nnd2s1 U4004 ( .Q(n3252), .DIN1(g416), .DIN2(n2077) );
  nnd2s1 U4005 ( .Q(g11268), .DIN1(n3254), .DIN2(n3255) );
  nnd2s1 U4006 ( .Q(n3255), .DIN1(g406), .DIN2(n3036) );
  nnd2s1 U4007 ( .Q(n3254), .DIN1(g411), .DIN2(n2078) );
  nnd2s1 U4008 ( .Q(g11267), .DIN1(n3256), .DIN2(n3257) );
  nnd2s1 U4009 ( .Q(n3257), .DIN1(g401), .DIN2(n2076) );
  nnd2s1 U4010 ( .Q(n3256), .DIN1(g406), .DIN2(n2079) );
  nnd2s1 U4011 ( .Q(g11266), .DIN1(n3258), .DIN2(n3259) );
  nnd2s1 U4012 ( .Q(n3259), .DIN1(g396), .DIN2(n3036) );
  nnd2s1 U4013 ( .Q(n3258), .DIN1(g401), .DIN2(n2079) );
  nnd2s1 U4014 ( .Q(g11265), .DIN1(n3260), .DIN2(n3261) );
  nnd2s1 U4015 ( .Q(n3261), .DIN1(g391), .DIN2(n3036) );
  nnd2s1 U4016 ( .Q(n3260), .DIN1(g396), .DIN2(n2077) );
  nnd2s1 U4017 ( .Q(g11264), .DIN1(n3262), .DIN2(n3263) );
  nnd2s1 U4018 ( .Q(n3263), .DIN1(g386), .DIN2(n3036) );
  nnd2s1 U4019 ( .Q(n3262), .DIN1(g391), .DIN2(n2078) );
  nnd2s1 U4020 ( .Q(g11263), .DIN1(n3264), .DIN2(n3265) );
  nnd2s1 U4021 ( .Q(n3265), .DIN1(g426), .DIN2(n2076) );
  nnd2s1 U4022 ( .Q(n3264), .DIN1(g386), .DIN2(n2077) );
  nnd2s1 U4023 ( .Q(g11262), .DIN1(n3266), .DIN2(n3267) );
  nnd2s1 U4024 ( .Q(n3267), .DIN1(g435), .DIN2(n2071) );
  nnd2s1 U4025 ( .Q(n3266), .DIN1(g431), .DIN2(n2077) );
  nnd2s1 U4026 ( .Q(g11261), .DIN1(n3268), .DIN2(n3269) );
  nnd2s1 U4027 ( .Q(n3269), .DIN1(g440), .DIN2(n2076) );
  nnd2s1 U4028 ( .Q(n3268), .DIN1(n2079), .DIN2(g435) );
  nnd2s1 U4029 ( .Q(g11260), .DIN1(n3270), .DIN2(n3271) );
  nnd2s1 U4030 ( .Q(n3271), .DIN1(g444), .DIN2(n3036) );
  nnd2s1 U4031 ( .Q(n3270), .DIN1(g440), .DIN2(n2079) );
  nnd2s1 U4032 ( .Q(g11259), .DIN1(n3272), .DIN2(n3273) );
  nnd2s1 U4033 ( .Q(n3273), .DIN1(g448), .DIN2(n2076) );
  nnd2s1 U4034 ( .Q(n3272), .DIN1(g444), .DIN2(n2077) );
  nnd2s1 U4035 ( .Q(g11258), .DIN1(n3274), .DIN2(n3275) );
  nnd2s1 U4036 ( .Q(n3275), .DIN1(g452), .DIN2(n2071) );
  nnd2s1 U4037 ( .Q(n3274), .DIN1(g448), .DIN2(n2079) );
  nnd2s1 U4038 ( .Q(g11257), .DIN1(n3276), .DIN2(n3277) );
  nnd2s1 U4039 ( .Q(n3277), .DIN1(g421), .DIN2(n3036) );
  nnd2s1 U4040 ( .Q(n3276), .DIN1(g452), .DIN2(n2078) );
  nnd2s1 U4041 ( .Q(g11256), .DIN1(n3278), .DIN2(n3279) );
  nnd2s1 U4042 ( .Q(n3279), .DIN1(n3280), .DIN2(n3036) );
  nnd2s1 U4043 ( .Q(n3278), .DIN1(g426), .DIN2(n2079) );
  nnd2s1 U4044 ( .Q(g11185), .DIN1(n3281), .DIN2(n3282) );
  nnd2s1 U4045 ( .Q(n3282), .DIN1(g1811), .DIN2(n2567) );
  hi1s1 U4046 ( .Q(n2567), .DIN(n2617) );
  nnd2s1 U4047 ( .Q(n3281), .DIN1(n2617), .DIN2(n3283) );
  nnd4s1 U4048 ( .Q(n3283), .DIN1(g10870), .DIN2(n3010), .DIN3(n3284), .DIN4(
        n3285) );
  and3s1 U4049 ( .Q(n3285), .DIN1(n3286), .DIN2(n3287), .DIN3(n3189) );
  nor2s1 U4050 ( .Q(g11184), .DIN1(n2617), .DIN2(n1967) );
  nor2s1 U4051 ( .Q(g11183), .DIN1(n2617), .DIN2(n2006) );
  nor2s1 U4052 ( .Q(g11182), .DIN1(n2617), .DIN2(n1928) );
  nor2s1 U4053 ( .Q(g11181), .DIN1(n2617), .DIN2(n1943) );
  nor2s1 U4054 ( .Q(n2617), .DIN1(n3288), .DIN2(g1703) );
  nnd2s1 U4055 ( .Q(g11180), .DIN1(n3289), .DIN2(n3290) );
  nnd2s1 U4056 ( .Q(n3290), .DIN1(g105), .DIN2(n2068) );
  nnd2s1 U4057 ( .Q(n3289), .DIN1(n2350), .DIN2(n3291) );
  or2s1 U4058 ( .Q(n3291), .DIN1(n3292), .DIN2(n2932) );
  hi1s1 U4059 ( .Q(n2932), .DIN(n2931) );
  nnd2s1 U4060 ( .Q(n2931), .DIN1(n3010), .DIN2(n3293) );
  nnd2s1 U4061 ( .Q(n3010), .DIN1(n2122), .DIN2(n2124) );
  and3s1 U4062 ( .Q(n2122), .DIN1(n2081), .DIN2(n2121), .DIN3(n2123) );
  and4s1 U4063 ( .Q(n2123), .DIN1(n3294), .DIN2(n2130), .DIN3(n2128), .DIN4(
        n2129) );
  xor2s1 U4064 ( .Q(n3292), .DIN1(n3295), .DIN2(n3296) );
  xor2s1 U4065 ( .Q(n3296), .DIN1(g991), .DIN2(g1019) );
  xor2s1 U4066 ( .Q(n3295), .DIN1(n3297), .DIN2(n3298) );
  xor2s1 U4067 ( .Q(n3298), .DIN1(n3299), .DIN2(n3300) );
  xor2s1 U4068 ( .Q(n3300), .DIN1(g1007), .DIN2(g1003) );
  xor2s1 U4069 ( .Q(n3299), .DIN1(g1015), .DIN2(g1011) );
  xor2s1 U4070 ( .Q(n3297), .DIN1(n3301), .DIN2(n3302) );
  xor2s1 U4071 ( .Q(n3302), .DIN1(g1027), .DIN2(g1023) );
  xor2s1 U4072 ( .Q(n3301), .DIN1(g999), .DIN2(g995) );
  hi1s1 U4073 ( .Q(g11179), .DIN(n3106) );
  nnd3s1 U4074 ( .Q(n3106), .DIN1(n3303), .DIN2(n2071), .DIN3(n3153) );
  hi1s1 U4075 ( .Q(n3036), .DIN(n2079) );
  or4s1 U4076 ( .Q(n3306), .DIN1(g845), .DIN2(g849), .DIN3(g841), .DIN4(n3307)
         );
  or3s1 U4077 ( .Q(n3307), .DIN1(g857), .DIN2(g861), .DIN3(g853) );
  or3s1 U4078 ( .Q(n3305), .DIN1(g833), .DIN2(g837), .DIN3(g829) );
  nor2s1 U4079 ( .Q(n3304), .DIN1(n3308), .DIN2(n3309) );
  nnd4s1 U4080 ( .Q(n3309), .DIN1(n3293), .DIN2(n3310), .DIN3(n3189), .DIN4(
        n3286) );
  nnd4s1 U4081 ( .Q(n3308), .DIN1(n3287), .DIN2(n3311), .DIN3(n3312), .DIN4(
        n3011) );
  or4s1 U4082 ( .Q(n3303), .DIN1(n3313), .DIN2(n3314), .DIN3(n3315), .DIN4(
        n3316) );
  or4s1 U4083 ( .Q(n3316), .DIN1(n3317), .DIN2(n3318), .DIN3(n3319), .DIN4(
        n3320) );
  or2s1 U4084 ( .Q(n3320), .DIN1(n3321), .DIN2(n3322) );
  xor2s1 U4085 ( .Q(n3322), .DIN1(g386), .DIN2(g318) );
  xor2s1 U4086 ( .Q(n3321), .DIN1(g426), .DIN2(g315) );
  xor2s1 U4087 ( .Q(n3319), .DIN1(g416), .DIN2(g309) );
  xor2s1 U4088 ( .Q(n3318), .DIN1(g421), .DIN2(g312) );
  xor2s1 U4089 ( .Q(n3317), .DIN1(g305), .DIN2(n3280) );
  nnd2s1 U4090 ( .Q(n3280), .DIN1(n3323), .DIN2(n3324) );
  nnd2s1 U4091 ( .Q(n3324), .DIN1(g305), .DIN2(n3325) );
  nnd2s1 U4092 ( .Q(n3323), .DIN1(n3326), .DIN2(n3153) );
  hi1s1 U4093 ( .Q(n3153), .DIN(n3325) );
  nnd2s1 U4094 ( .Q(n3325), .DIN1(g382), .DIN2(n3149) );
  hi1s1 U4095 ( .Q(n3149), .DIN(n3141) );
  nnd3s1 U4096 ( .Q(n3141), .DIN1(g374), .DIN2(g369), .DIN3(g378) );
  nnd2s1 U4097 ( .Q(n3326), .DIN1(n3327), .DIN2(n3328) );
  nnd2s1 U4098 ( .Q(n3328), .DIN1(g431), .DIN2(n2033) );
  nnd2s1 U4099 ( .Q(n3327), .DIN1(n3329), .DIN2(n2054) );
  nnd2s1 U4100 ( .Q(n3329), .DIN1(n2033), .DIN2(n3330) );
  or4s1 U4101 ( .Q(n3330), .DIN1(n3331), .DIN2(n3332), .DIN3(n3333), .DIN4(
        n3334) );
  or3s1 U4102 ( .Q(n3334), .DIN1(g421), .DIN2(g426), .DIN3(g416) );
  or4s1 U4103 ( .Q(n3333), .DIN1(g440), .DIN2(g444), .DIN3(g448), .DIN4(g452)
         );
  or3s1 U4104 ( .Q(n3332), .DIN1(g391), .DIN2(g396), .DIN3(g386) );
  or3s1 U4105 ( .Q(n3331), .DIN1(g406), .DIN2(g411), .DIN3(g401) );
  or3s1 U4106 ( .Q(n3315), .DIN1(n3335), .DIN2(n3336), .DIN3(n3337) );
  xor2s1 U4107 ( .Q(n3337), .DIN1(g396), .DIN2(g324) );
  xor2s1 U4108 ( .Q(n3336), .DIN1(g401), .DIN2(g327) );
  xor2s1 U4109 ( .Q(n3335), .DIN1(g391), .DIN2(g321) );
  xor2s1 U4110 ( .Q(n3314), .DIN1(g411), .DIN2(g333) );
  xor2s1 U4111 ( .Q(n3313), .DIN1(g406), .DIN2(g330) );
  nnd2s1 U4112 ( .Q(g11052), .DIN1(n3338), .DIN2(n3339) );
  nnd2s1 U4113 ( .Q(n3339), .DIN1(g575), .DIN2(n2069) );
  nnd2s1 U4114 ( .Q(n3338), .DIN1(n2063), .DIN2(n3340) );
  nnd2s1 U4115 ( .Q(g11051), .DIN1(n3341), .DIN2(n3342) );
  nnd2s1 U4116 ( .Q(n3342), .DIN1(g566), .DIN2(n2070) );
  nnd2s1 U4117 ( .Q(g11050), .DIN1(n3343), .DIN2(n3344) );
  nnd2s1 U4118 ( .Q(n3344), .DIN1(g563), .DIN2(n2068) );
  nnd2s1 U4119 ( .Q(g11049), .DIN1(n3345), .DIN2(n3346) );
  nnd2s1 U4120 ( .Q(n3346), .DIN1(g560), .DIN2(n2069) );
  nnd2s1 U4121 ( .Q(g11048), .DIN1(n3347), .DIN2(n3348) );
  nnd2s1 U4122 ( .Q(n3348), .DIN1(g557), .DIN2(n2069) );
  nnd2s1 U4123 ( .Q(g11047), .DIN1(n3349), .DIN2(n3350) );
  nnd2s1 U4124 ( .Q(n3350), .DIN1(g554), .DIN2(n2068) );
  nnd2s1 U4125 ( .Q(g11044), .DIN1(n3351), .DIN2(n3352) );
  nnd2s1 U4126 ( .Q(n3352), .DIN1(g549), .DIN2(n2069) );
  nnd2s1 U4127 ( .Q(n3351), .DIN1(n2350), .DIN2(n3353) );
  nnd2s1 U4128 ( .Q(g11043), .DIN1(n3354), .DIN2(n3355) );
  nnd2s1 U4129 ( .Q(n3355), .DIN1(g546), .DIN2(n2068) );
  nnd2s1 U4130 ( .Q(g11042), .DIN1(n3341), .DIN2(n3356) );
  nnd2s1 U4131 ( .Q(n3356), .DIN1(g1687), .DIN2(n2070) );
  nnd2s1 U4132 ( .Q(n3341), .DIN1(n2350), .DIN2(n3357) );
  nnd2s1 U4133 ( .Q(n3357), .DIN1(n3358), .DIN2(n3359) );
  nnd2s1 U4134 ( .Q(n3359), .DIN1(n3360), .DIN2(n2469) );
  nnd2s1 U4135 ( .Q(n2469), .DIN1(n2358), .DIN2(n3361) );
  nnd2s1 U4136 ( .Q(n3361), .DIN1(g1627), .DIN2(n2082) );
  nnd2s1 U4137 ( .Q(n2358), .DIN1(g231), .DIN2(g18) );
  nnd2s1 U4138 ( .Q(n3358), .DIN1(n3362), .DIN2(n3363) );
  nnd2s1 U4139 ( .Q(n3363), .DIN1(g109), .DIN2(n3011) );
  nnd2s1 U4140 ( .Q(g11041), .DIN1(n3343), .DIN2(n3364) );
  nnd2s1 U4141 ( .Q(n3364), .DIN1(g1684), .DIN2(n2068) );
  nnd2s1 U4142 ( .Q(n3343), .DIN1(n2063), .DIN2(n3365) );
  nnd2s1 U4143 ( .Q(n3365), .DIN1(n3366), .DIN2(n3367) );
  nnd2s1 U4144 ( .Q(n3367), .DIN1(n3360), .DIN2(n2467) );
  nnd2s1 U4145 ( .Q(n2467), .DIN1(n2364), .DIN2(n3368) );
  nnd2s1 U4146 ( .Q(n3368), .DIN1(g1624), .DIN2(n2072) );
  nnd2s1 U4147 ( .Q(n2364), .DIN1(g225), .DIN2(g18) );
  nnd2s1 U4148 ( .Q(n3366), .DIN1(n3362), .DIN2(n3181) );
  nnd2s1 U4149 ( .Q(g11040), .DIN1(n3345), .DIN2(n3369) );
  nnd2s1 U4150 ( .Q(n3369), .DIN1(g1681), .DIN2(n2070) );
  nnd4s1 U4151 ( .Q(n3345), .DIN1(n2063), .DIN2(n3370), .DIN3(n3371), .DIN4(
        n3372) );
  nnd2s1 U4152 ( .Q(n3372), .DIN1(n3373), .DIN2(n3311) );
  nnd2s1 U4153 ( .Q(n3371), .DIN1(n2465), .DIN2(n3360) );
  and2s1 U4154 ( .Q(n2465), .DIN1(n2371), .DIN2(n3374) );
  nnd2s1 U4155 ( .Q(n3374), .DIN1(g1621), .DIN2(n2082) );
  nnd2s1 U4156 ( .Q(n2371), .DIN1(g219), .DIN2(g18) );
  nnd2s1 U4157 ( .Q(g11039), .DIN1(n3347), .DIN2(n3375) );
  nnd2s1 U4158 ( .Q(n3375), .DIN1(g1678), .DIN2(n2070) );
  nnd4s1 U4159 ( .Q(n3347), .DIN1(n2350), .DIN2(n3370), .DIN3(n3376), .DIN4(
        n3377) );
  nnd2s1 U4160 ( .Q(n3377), .DIN1(n3373), .DIN2(n3287) );
  nnd2s1 U4161 ( .Q(n3376), .DIN1(n2463), .DIN2(n3360) );
  and2s1 U4162 ( .Q(n2463), .DIN1(n2377), .DIN2(n3378) );
  nnd2s1 U4163 ( .Q(n3378), .DIN1(g1615), .DIN2(n2082) );
  nnd2s1 U4164 ( .Q(n2377), .DIN1(g213), .DIN2(g18) );
  nnd2s1 U4165 ( .Q(g11038), .DIN1(n3349), .DIN2(n3379) );
  nnd2s1 U4166 ( .Q(n3379), .DIN1(g1675), .DIN2(n2068) );
  nnd3s1 U4167 ( .Q(n3349), .DIN1(n3380), .DIN2(n3381), .DIN3(n2350) );
  nnd3s1 U4168 ( .Q(n3381), .DIN1(g109), .DIN2(n3286), .DIN3(n3362) );
  nnd2s1 U4169 ( .Q(n3380), .DIN1(n3360), .DIN2(n2461) );
  and2s1 U4170 ( .Q(n2461), .DIN1(n2384), .DIN2(n3382) );
  nnd2s1 U4171 ( .Q(n3382), .DIN1(g1639), .DIN2(n2082) );
  nnd2s1 U4172 ( .Q(n2384), .DIN1(g207), .DIN2(g18) );
  nnd2s1 U4173 ( .Q(g11037), .DIN1(n3354), .DIN2(n3383) );
  nnd2s1 U4174 ( .Q(n3383), .DIN1(g1672), .DIN2(n2069) );
  nnd2s1 U4175 ( .Q(n3354), .DIN1(n2063), .DIN2(n3384) );
  nnd2s1 U4176 ( .Q(n3384), .DIN1(n3385), .DIN2(n3386) );
  nnd3s1 U4177 ( .Q(n3386), .DIN1(g109), .DIN2(g10867), .DIN3(n3362) );
  nnd2s1 U4178 ( .Q(n3385), .DIN1(n3360), .DIN2(n2459) );
  nnd2s1 U4179 ( .Q(n2459), .DIN1(n2390), .DIN2(n3387) );
  nnd2s1 U4180 ( .Q(n3387), .DIN1(g1618), .DIN2(n2072) );
  nnd2s1 U4181 ( .Q(n2390), .DIN1(g186), .DIN2(g18) );
  nnd2s1 U4182 ( .Q(g11036), .DIN1(n3388), .DIN2(n3389) );
  nnd2s1 U4183 ( .Q(n3389), .DIN1(g1669), .DIN2(n2839) );
  nnd3s1 U4184 ( .Q(n3388), .DIN1(n3362), .DIN2(n3390), .DIN3(n2840) );
  nnd2s1 U4185 ( .Q(n3390), .DIN1(g109), .DIN2(n3311) );
  nnd2s1 U4186 ( .Q(g11035), .DIN1(n3391), .DIN2(n3392) );
  nnd2s1 U4187 ( .Q(n3392), .DIN1(g1666), .DIN2(n2839) );
  nnd2s1 U4188 ( .Q(n3391), .DIN1(n2840), .DIN2(n3393) );
  nnd2s1 U4189 ( .Q(n3393), .DIN1(n1979), .DIN2(n3394) );
  nnd2s1 U4190 ( .Q(n3394), .DIN1(n3395), .DIN2(g10869) );
  nnd2s1 U4191 ( .Q(g11034), .DIN1(n3396), .DIN2(n3397) );
  nnd2s1 U4192 ( .Q(n3397), .DIN1(g1663), .DIN2(n2839) );
  nnd2s1 U4193 ( .Q(n3396), .DIN1(n2840), .DIN2(n3353) );
  nnd3s1 U4194 ( .Q(n3353), .DIN1(n3398), .DIN2(n1979), .DIN3(n3399) );
  nnd2s1 U4195 ( .Q(n3399), .DIN1(n3360), .DIN2(n2477) );
  nnd2s1 U4196 ( .Q(n2477), .DIN1(n2695), .DIN2(n3400) );
  nnd2s1 U4197 ( .Q(n3400), .DIN1(g1512), .DIN2(n2082) );
  nnd2s1 U4198 ( .Q(n2695), .DIN1(g192), .DIN2(g18) );
  nnd2s1 U4199 ( .Q(n3398), .DIN1(n3395), .DIN2(g10868) );
  nnd2s1 U4200 ( .Q(g11033), .DIN1(n3401), .DIN2(n3402) );
  nnd2s1 U4201 ( .Q(n3402), .DIN1(g1660), .DIN2(n2839) );
  nnd2s1 U4202 ( .Q(n3401), .DIN1(n2840), .DIN2(n3340) );
  nnd3s1 U4203 ( .Q(n3340), .DIN1(n3403), .DIN2(n3404), .DIN3(n3370) );
  nnd2s1 U4204 ( .Q(n3370), .DIN1(n3405), .DIN2(n3373) );
  nnd2s1 U4205 ( .Q(n3405), .DIN1(g109), .DIN2(n1979) );
  nnd2s1 U4206 ( .Q(n3404), .DIN1(g10867), .DIN2(n3373) );
  hi1s1 U4207 ( .Q(n3373), .DIN(n3360) );
  nnd2s1 U4208 ( .Q(n3403), .DIN1(n2475), .DIN2(n3360) );
  nnd2s1 U4209 ( .Q(n2475), .DIN1(n2685), .DIN2(n3406) );
  nnd2s1 U4210 ( .Q(n3406), .DIN1(g1636), .DIN2(n2072) );
  nnd2s1 U4211 ( .Q(n2685), .DIN1(g248), .DIN2(g18) );
  nnd2s1 U4212 ( .Q(g10882), .DIN1(n3407), .DIN2(n3408) );
  nnd2s1 U4213 ( .Q(n3408), .DIN1(g1733), .DIN2(n3409) );
  nnd2s1 U4214 ( .Q(n3407), .DIN1(n2833), .DIN2(n3181) );
  hi1s1 U4215 ( .Q(n3181), .DIN(n3284) );
  nor2s1 U4216 ( .Q(n3284), .DIN1(n2064), .DIN2(g10871) );
  hi1s1 U4217 ( .Q(n2833), .DIN(n3409) );
  nnd2s1 U4218 ( .Q(g10881), .DIN1(n3410), .DIN2(n3411) );
  nnd2s1 U4219 ( .Q(n3411), .DIN1(n3412), .DIN2(g10870) );
  nnd2s1 U4220 ( .Q(n3410), .DIN1(g1730), .DIN2(n3409) );
  nnd2s1 U4221 ( .Q(g10880), .DIN1(n3413), .DIN2(n3414) );
  nnd2s1 U4222 ( .Q(n3414), .DIN1(n3412), .DIN2(g10869) );
  nnd2s1 U4223 ( .Q(n3413), .DIN1(g1727), .DIN2(n3409) );
  nnd2s1 U4224 ( .Q(g10879), .DIN1(n3415), .DIN2(n3416) );
  nnd2s1 U4225 ( .Q(n3416), .DIN1(n3412), .DIN2(g10868) );
  nnd2s1 U4226 ( .Q(n3415), .DIN1(g1724), .DIN2(n3409) );
  nnd2s1 U4227 ( .Q(g10878), .DIN1(n3417), .DIN2(n3418) );
  nnd2s1 U4228 ( .Q(n3418), .DIN1(n3412), .DIN2(g10867) );
  nor2s1 U4229 ( .Q(n3412), .DIN1(n3409), .DIN2(n2065) );
  nnd2s1 U4230 ( .Q(n3417), .DIN1(g1721), .DIN2(n3409) );
  nnd2s1 U4231 ( .Q(n3409), .DIN1(g1703), .DIN2(g1696) );
  nnd2s1 U4232 ( .Q(g10877), .DIN1(n3419), .DIN2(n3420) );
  nnd2s1 U4233 ( .Q(n3420), .DIN1(g572), .DIN2(n2069) );
  nnd2s1 U4234 ( .Q(n3419), .DIN1(n2063), .DIN2(n3421) );
  nnd2s1 U4235 ( .Q(g10876), .DIN1(n3422), .DIN2(n3423) );
  nnd2s1 U4236 ( .Q(n3423), .DIN1(g569), .DIN2(n2069) );
  nnd2s1 U4237 ( .Q(n3422), .DIN1(n2350), .DIN2(n3424) );
  nor2s1 U4238 ( .Q(n2350), .DIN1(g1696), .DIN2(g1703) );
  nnd2s1 U4239 ( .Q(g10875), .DIN1(n3425), .DIN2(n3426) );
  nnd2s1 U4240 ( .Q(n3426), .DIN1(g1657), .DIN2(n2839) );
  nnd2s1 U4241 ( .Q(n3425), .DIN1(n2840), .DIN2(n3421) );
  nnd3s1 U4242 ( .Q(n3421), .DIN1(n3427), .DIN2(n1979), .DIN3(n3428) );
  nnd2s1 U4243 ( .Q(n3428), .DIN1(n3360), .DIN2(n2473) );
  nnd2s1 U4244 ( .Q(n2473), .DIN1(n2687), .DIN2(n3429) );
  nnd2s1 U4245 ( .Q(n3429), .DIN1(g1633), .DIN2(n2082) );
  nnd2s1 U4246 ( .Q(n2687), .DIN1(g243), .DIN2(g18) );
  nnd2s1 U4247 ( .Q(n3427), .DIN1(n3395), .DIN2(g10775) );
  nor2s1 U4248 ( .Q(n3395), .DIN1(n2066), .DIN2(n3360) );
  nnd2s1 U4249 ( .Q(g10874), .DIN1(n3430), .DIN2(n3431) );
  nnd2s1 U4250 ( .Q(n3431), .DIN1(g1654), .DIN2(n2839) );
  nnd2s1 U4251 ( .Q(n3430), .DIN1(n2840), .DIN2(n3424) );
  nnd2s1 U4252 ( .Q(n3424), .DIN1(n3432), .DIN2(n3433) );
  nnd2s1 U4253 ( .Q(n3433), .DIN1(n3362), .DIN2(n3434) );
  nnd2s1 U4254 ( .Q(n3434), .DIN1(g109), .DIN2(n3293) );
  nor2s1 U4255 ( .Q(n3362), .DIN1(n3360), .DIN2(g1718) );
  nnd2s1 U4256 ( .Q(n3432), .DIN1(n3360), .DIN2(n2471) );
  nnd2s1 U4257 ( .Q(n2471), .DIN1(n2351), .DIN2(n3435) );
  nnd2s1 U4258 ( .Q(n3435), .DIN1(g1630), .DIN2(n2072) );
  hi1s1 U4259 ( .Q(n2082), .DIN(g18) );
  nnd2s1 U4260 ( .Q(n2351), .DIN1(g237), .DIN2(g18) );
  nor2s1 U4261 ( .Q(n3360), .DIN1(g1357), .DIN2(g1718) );
  hi1s1 U4262 ( .Q(n2840), .DIN(n2839) );
  nnd2s1 U4263 ( .Q(n2839), .DIN1(g1703), .DIN2(n3288) );
  hi1s1 U4264 ( .Q(n3288), .DIN(g1696) );
  hi1s1 U4265 ( .Q(g10872), .DIN(n3011) );
  hi1s1 U4266 ( .Q(g10869), .DIN(n3287) );
  xor2s1 U4267 ( .Q(g10779), .DIN1(n3211), .DIN2(n3436) );
  nnd2s1 U4268 ( .Q(g10712), .DIN1(n3437), .DIN2(n3211) );
  nnd2s1 U4269 ( .Q(n3211), .DIN1(n3438), .DIN2(n3439) );
  nnd2s1 U4270 ( .Q(n3439), .DIN1(n3440), .DIN2(n3441) );
  nnd2s1 U4271 ( .Q(n3441), .DIN1(n3442), .DIN2(n2030) );
  hi1s1 U4272 ( .Q(n3440), .DIN(n3443) );
  nnd3s1 U4273 ( .Q(n3438), .DIN1(n3442), .DIN2(n2030), .DIN3(n3443) );
  xor2s1 U4274 ( .Q(n3443), .DIN1(n3444), .DIN2(n3445) );
  xor2s1 U4275 ( .Q(n3445), .DIN1(n3446), .DIN2(n3447) );
  xor2s1 U4276 ( .Q(n3447), .DIN1(g10867), .DIN2(n3286) );
  xor2s1 U4277 ( .Q(n3446), .DIN1(n3287), .DIN2(g10870) );
  xor2s1 U4278 ( .Q(n3444), .DIN1(n3448), .DIN2(n3449) );
  xor2s1 U4279 ( .Q(n3449), .DIN1(g10871), .DIN2(n3310) );
  xor2s1 U4280 ( .Q(n3448), .DIN1(n3011), .DIN2(n3293) );
  nor2s1 U4281 ( .Q(g10583), .DIN1(n3450), .DIN2(n3436) );
  nnd2s1 U4282 ( .Q(n3436), .DIN1(n3451), .DIN2(n3452) );
  nnd2s1 U4283 ( .Q(n3452), .DIN1(g109), .DIN2(n3453) );
  nnd4s1 U4284 ( .Q(n3453), .DIN1(n3454), .DIN2(n3455), .DIN3(n3456), .DIN4(
        n3457) );
  nnd2s1 U4285 ( .Q(n3457), .DIN1(n2834), .DIN2(g10871) );
  hi1s1 U4286 ( .Q(g10871), .DIN(n3312) );
  hi1s1 U4287 ( .Q(n2834), .DIN(n2923) );
  nnd3s1 U4288 ( .Q(n2923), .DIN1(g109), .DIN2(\DFF_194/net481 ), .DIN3(g3069)
         );
  nnd2s1 U4289 ( .Q(n3456), .DIN1(g865), .DIN2(g10775) );
  hi1s1 U4290 ( .Q(g10775), .DIN(n3310) );
  nnd2s1 U4291 ( .Q(n3455), .DIN1(g108), .DIN2(g10870) );
  hi1s1 U4292 ( .Q(g10870), .DIN(n3311) );
  or2s1 U4293 ( .Q(n3454), .DIN1(n3011), .DIN2(g105) );
  nnd2s1 U4294 ( .Q(n3451), .DIN1(g6846), .DIN2(g10774) );
  nor2s1 U4295 ( .Q(g6846), .DIN1(n2877), .DIN2(n2065) );
  nnd2s1 U4296 ( .Q(n2877), .DIN1(g1765), .DIN2(g1610) );
  hi1s1 U4297 ( .Q(n3450), .DIN(g10515) );
  nnd2s1 U4298 ( .Q(g10515), .DIN1(g109), .DIN2(n3458) );
  nnd4s1 U4299 ( .Q(n3458), .DIN1(n3459), .DIN2(n3460), .DIN3(n3461), .DIN4(
        n3462) );
  or2s1 U4300 ( .Q(n3462), .DIN1(n3105), .DIN2(n3311) );
  nnd2s1 U4301 ( .Q(n3105), .DIN1(g757), .DIN2(g109) );
  nor2s1 U4302 ( .Q(n3461), .DIN1(n3463), .DIN2(n3464) );
  nor2s1 U4303 ( .Q(n3464), .DIN1(n3287), .DIN2(n2438) );
  nnd3s1 U4304 ( .Q(n2438), .DIN1(g109), .DIN2(\DFF_121/net408 ), .DIN3(g2986)
         );
  nor2s1 U4305 ( .Q(n3463), .DIN1(n3312), .DIN2(n3104) );
  nnd2s1 U4306 ( .Q(n3104), .DIN1(g3007), .DIN2(\DFF_93/net380 ) );
  nnd2s1 U4307 ( .Q(n3460), .DIN1(g877), .DIN2(g10867) );
  hi1s1 U4308 ( .Q(g10867), .DIN(n3189) );
  nnd2s1 U4309 ( .Q(n3459), .DIN1(g881), .DIN2(g10868) );
  hi1s1 U4310 ( .Q(g10868), .DIN(n3286) );
  nnd2s1 U4311 ( .Q(g10417), .DIN1(n3437), .DIN2(n3011) );
  nor4s1 U4312 ( .Q(n3011), .DIN1(n3465), .DIN2(n3466), .DIN3(n3467), .DIN4(
        n3468) );
  nnd3s1 U4313 ( .Q(n3468), .DIN1(n3469), .DIN2(n3470), .DIN3(n3471) );
  nnd2s1 U4314 ( .Q(n3471), .DIN1(n3472), .DIN2(g1607) );
  nnd2s1 U4315 ( .Q(n3470), .DIN1(g913), .DIN2(n3473) );
  nnd2s1 U4316 ( .Q(n3469), .DIN1(n3474), .DIN2(g1583) );
  nnd4s1 U4317 ( .Q(n3467), .DIN1(n3475), .DIN2(n3476), .DIN3(n3477), .DIN4(
        n3478) );
  nnd2s1 U4318 ( .Q(n3478), .DIN1(n3479), .DIN2(n3480) );
  nnd2s1 U4319 ( .Q(n3477), .DIN1(g1330), .DIN2(n3481) );
  nnd2s1 U4320 ( .Q(n3476), .DIN1(g1185), .DIN2(n3482) );
  nnd2s1 U4321 ( .Q(n3475), .DIN1(g965), .DIN2(n3483) );
  nnd3s1 U4322 ( .Q(n3466), .DIN1(n3484), .DIN2(n3485), .DIN3(n3486) );
  nnd2s1 U4323 ( .Q(n3486), .DIN1(g38), .DIN2(n3442) );
  nnd2s1 U4324 ( .Q(n3485), .DIN1(n3487), .DIN2(g302) );
  nnd2s1 U4325 ( .Q(n3484), .DIN1(n3488), .DIN2(g1759) );
  nnd3s1 U4326 ( .Q(n3465), .DIN1(n3489), .DIN2(n3490), .DIN3(n3491) );
  nnd2s1 U4327 ( .Q(n3491), .DIN1(n3492), .DIN2(g278) );
  nnd2s1 U4328 ( .Q(n3490), .DIN1(n3493), .DIN2(g1540) );
  nnd2s1 U4329 ( .Q(n3489), .DIN1(n3494), .DIN2(g1564) );
  nnd2s1 U4330 ( .Q(g10414), .DIN1(n3437), .DIN2(n3312) );
  nor4s1 U4331 ( .Q(n3312), .DIN1(n3495), .DIN2(n3496), .DIN3(n3497), .DIN4(
        n3498) );
  nnd4s1 U4332 ( .Q(n3498), .DIN1(n3499), .DIN2(n3500), .DIN3(n3501), .DIN4(
        n3502) );
  nnd2s1 U4333 ( .Q(n3502), .DIN1(n3474), .DIN2(g1580) );
  nnd2s1 U4334 ( .Q(n3501), .DIN1(n3472), .DIN2(g1604) );
  nnd2s1 U4335 ( .Q(n3500), .DIN1(n3493), .DIN2(g1537) );
  nnd2s1 U4336 ( .Q(n3499), .DIN1(n3494), .DIN2(g1561) );
  nnd4s1 U4337 ( .Q(n3497), .DIN1(n3503), .DIN2(n3504), .DIN3(n3505), .DIN4(
        n3506) );
  nnd2s1 U4338 ( .Q(n3506), .DIN1(g1327), .DIN2(n3481) );
  nnd2s1 U4339 ( .Q(n3505), .DIN1(g1182), .DIN2(n3482) );
  nnd2s1 U4340 ( .Q(n3504), .DIN1(g962), .DIN2(n3483) );
  nnd2s1 U4341 ( .Q(n3503), .DIN1(g910), .DIN2(n3473) );
  nnd4s1 U4342 ( .Q(n3496), .DIN1(n3507), .DIN2(n3508), .DIN3(n3509), .DIN4(
        n3510) );
  nnd4s1 U4343 ( .Q(n3510), .DIN1(n3511), .DIN2(n3480), .DIN3(n3479), .DIN4(
        n3512) );
  nnd2s1 U4344 ( .Q(n3509), .DIN1(g16), .DIN2(n3513) );
  nnd2s1 U4345 ( .Q(n3508), .DIN1(g37), .DIN2(n3442) );
  nnd2s1 U4346 ( .Q(n3507), .DIN1(g7), .DIN2(n3514) );
  nnd4s1 U4347 ( .Q(n3495), .DIN1(n3515), .DIN2(n3516), .DIN3(n3517), .DIN4(
        n3518) );
  nnd2s1 U4348 ( .Q(n3518), .DIN1(n3492), .DIN2(g275) );
  nnd2s1 U4349 ( .Q(n3517), .DIN1(n3487), .DIN2(g299) );
  nnd2s1 U4350 ( .Q(n3516), .DIN1(g1733), .DIN2(n3519) );
  nnd2s1 U4351 ( .Q(n3515), .DIN1(n3488), .DIN2(g1756) );
  nnd2s1 U4352 ( .Q(g10411), .DIN1(n3437), .DIN2(n3311) );
  nor4s1 U4353 ( .Q(n3311), .DIN1(n3520), .DIN2(n3521), .DIN3(n3522), .DIN4(
        n3523) );
  nnd4s1 U4354 ( .Q(n3523), .DIN1(n3524), .DIN2(n3525), .DIN3(n3526), .DIN4(
        n3527) );
  and2s1 U4355 ( .Q(n3527), .DIN1(n3528), .DIN2(n3529) );
  nnd2s1 U4356 ( .Q(n3529), .DIN1(n3530), .DIN2(g986) );
  nnd2s1 U4357 ( .Q(n3528), .DIN1(g907), .DIN2(n3473) );
  nnd2s1 U4358 ( .Q(n3526), .DIN1(g959), .DIN2(n3483) );
  nnd2s1 U4359 ( .Q(n3525), .DIN1(g1324), .DIN2(n3481) );
  nnd2s1 U4360 ( .Q(n3524), .DIN1(g1179), .DIN2(n3482) );
  nnd4s1 U4361 ( .Q(n3522), .DIN1(n3531), .DIN2(n3532), .DIN3(n3533), .DIN4(
        n3534) );
  and3s1 U4362 ( .Q(n3534), .DIN1(n3535), .DIN2(n3536), .DIN3(n3537) );
  nnd2s1 U4363 ( .Q(n3537), .DIN1(n3538), .DIN2(g940) );
  nnd2s1 U4364 ( .Q(n3536), .DIN1(g17), .DIN2(n3513) );
  nnd2s1 U4365 ( .Q(n3535), .DIN1(g895), .DIN2(n3539) );
  nnd2s1 U4366 ( .Q(n3533), .DIN1(g8), .DIN2(n3514) );
  nnd2s1 U4367 ( .Q(n3531), .DIN1(g1203), .DIN2(n3540) );
  nnd4s1 U4368 ( .Q(n3521), .DIN1(n3541), .DIN2(n3542), .DIN3(n3543), .DIN4(
        n3544) );
  nor2s1 U4369 ( .Q(n3544), .DIN1(n3545), .DIN2(n3546) );
  nor2s1 U4370 ( .Q(n3546), .DIN1(n3547), .DIN2(\DFF_228/net515 ) );
  and2s1 U4371 ( .Q(n3545), .DIN1(g1753), .DIN2(n3488) );
  nnd2s1 U4372 ( .Q(n3543), .DIN1(g1730), .DIN2(n3519) );
  nnd2s1 U4373 ( .Q(n3542), .DIN1(n3492), .DIN2(g272) );
  nnd2s1 U4374 ( .Q(n3541), .DIN1(n3487), .DIN2(g296) );
  nnd4s1 U4375 ( .Q(n3520), .DIN1(n3548), .DIN2(n3549), .DIN3(n3550), .DIN4(
        n3551) );
  nnd2s1 U4376 ( .Q(n3551), .DIN1(n3472), .DIN2(g1601) );
  nor2s1 U4377 ( .Q(n3550), .DIN1(n3552), .DIN2(n3553) );
  and2s1 U4378 ( .Q(n3553), .DIN1(g1577), .DIN2(n3474) );
  and2s1 U4379 ( .Q(n3552), .DIN1(g1351), .DIN2(n3554) );
  nnd2s1 U4380 ( .Q(n3549), .DIN1(n3493), .DIN2(g1534) );
  nnd2s1 U4381 ( .Q(n3548), .DIN1(n3494), .DIN2(g1558) );
  nnd2s1 U4382 ( .Q(g10408), .DIN1(n3437), .DIN2(n3287) );
  nor4s1 U4383 ( .Q(n3287), .DIN1(n3555), .DIN2(n3556), .DIN3(n3557), .DIN4(
        n3558) );
  nnd4s1 U4384 ( .Q(n3558), .DIN1(n3559), .DIN2(n3560), .DIN3(n3561), .DIN4(
        n3562) );
  and2s1 U4385 ( .Q(n3562), .DIN1(n3563), .DIN2(n3564) );
  nnd2s1 U4386 ( .Q(n3564), .DIN1(n3530), .DIN2(g981) );
  nnd2s1 U4387 ( .Q(n3563), .DIN1(g904), .DIN2(n3473) );
  nnd2s1 U4388 ( .Q(n3561), .DIN1(g956), .DIN2(n3483) );
  nnd2s1 U4389 ( .Q(n3560), .DIN1(g1321), .DIN2(n3481) );
  nnd2s1 U4390 ( .Q(n3559), .DIN1(g1176), .DIN2(n3482) );
  nnd4s1 U4391 ( .Q(n3557), .DIN1(n3565), .DIN2(n3532), .DIN3(n3566), .DIN4(
        n3567) );
  and3s1 U4392 ( .Q(n3567), .DIN1(n3568), .DIN2(n3569), .DIN3(n3570) );
  nnd2s1 U4393 ( .Q(n3570), .DIN1(n3538), .DIN2(g936) );
  nnd2s1 U4394 ( .Q(n3569), .DIN1(n3513), .DIN2(g9) );
  nnd2s1 U4395 ( .Q(n3568), .DIN1(g892), .DIN2(n3539) );
  nnd2s1 U4396 ( .Q(n3566), .DIN1(n3514), .DIN2(g1) );
  nnd2s1 U4397 ( .Q(n3565), .DIN1(g1200), .DIN2(n3540) );
  nnd4s1 U4398 ( .Q(n3556), .DIN1(n3571), .DIN2(n3572), .DIN3(n3573), .DIN4(
        n3574) );
  nor2s1 U4399 ( .Q(n3574), .DIN1(n3575), .DIN2(n3576) );
  nor2s1 U4400 ( .Q(n3576), .DIN1(n3547), .DIN2(\DFF_242/net529 ) );
  and2s1 U4401 ( .Q(n3575), .DIN1(g1750), .DIN2(n3488) );
  nnd2s1 U4402 ( .Q(n3573), .DIN1(g1727), .DIN2(n3519) );
  nnd2s1 U4403 ( .Q(n3572), .DIN1(n3492), .DIN2(g269) );
  nnd2s1 U4404 ( .Q(n3571), .DIN1(n3487), .DIN2(g293) );
  nnd4s1 U4405 ( .Q(n3555), .DIN1(n3577), .DIN2(n3578), .DIN3(n3579), .DIN4(
        n3580) );
  nnd2s1 U4406 ( .Q(n3580), .DIN1(n3472), .DIN2(g1598) );
  nor2s1 U4407 ( .Q(n3579), .DIN1(n3581), .DIN2(n3582) );
  and2s1 U4408 ( .Q(n3582), .DIN1(g1574), .DIN2(n3474) );
  nor2s1 U4409 ( .Q(n3581), .DIN1(n2000), .DIN2(n3583) );
  nnd2s1 U4410 ( .Q(n3578), .DIN1(n3493), .DIN2(g1531) );
  nnd2s1 U4411 ( .Q(n3577), .DIN1(n3494), .DIN2(g1555) );
  nnd2s1 U4412 ( .Q(g10405), .DIN1(n3437), .DIN2(n3286) );
  nor4s1 U4413 ( .Q(n3286), .DIN1(n3584), .DIN2(n3585), .DIN3(n3586), .DIN4(
        n3587) );
  nnd4s1 U4414 ( .Q(n3587), .DIN1(n3588), .DIN2(n3589), .DIN3(n3590), .DIN4(
        n3591) );
  nnd2s1 U4415 ( .Q(n3591), .DIN1(g1173), .DIN2(n3482) );
  nor2s1 U4416 ( .Q(n3590), .DIN1(n3592), .DIN2(n3593) );
  and2s1 U4417 ( .Q(n3593), .DIN1(n3481), .DIN2(g1318) );
  nor2s1 U4418 ( .Q(n3592), .DIN1(n2007), .DIN2(n3594) );
  nnd2s1 U4419 ( .Q(n3589), .DIN1(g953), .DIN2(n3483) );
  nnd2s1 U4420 ( .Q(n3588), .DIN1(n3530), .DIN2(g976) );
  nnd4s1 U4421 ( .Q(n3586), .DIN1(n3595), .DIN2(n3532), .DIN3(n3596), .DIN4(
        n3597) );
  and3s1 U4422 ( .Q(n3597), .DIN1(n3598), .DIN2(n3599), .DIN3(n3600) );
  nnd2s1 U4423 ( .Q(n3600), .DIN1(g889), .DIN2(n3539) );
  nnd2s1 U4424 ( .Q(n3599), .DIN1(n3514), .DIN2(g4) );
  nnd2s1 U4425 ( .Q(n3598), .DIN1(n3513), .DIN2(g12) );
  nnd2s1 U4426 ( .Q(n3596), .DIN1(g1197), .DIN2(n3540) );
  nnd2s1 U4427 ( .Q(n3595), .DIN1(g925), .DIN2(n3601) );
  nnd4s1 U4428 ( .Q(n3585), .DIN1(n3602), .DIN2(n3603), .DIN3(n3604), .DIN4(
        n3605) );
  nor2s1 U4429 ( .Q(n3605), .DIN1(n3606), .DIN2(n3607) );
  nor2s1 U4430 ( .Q(n3607), .DIN1(n3547), .DIN2(\DFF_384/net671 ) );
  and2s1 U4431 ( .Q(n3606), .DIN1(g1747), .DIN2(n3488) );
  nnd2s1 U4432 ( .Q(n3604), .DIN1(g1724), .DIN2(n3519) );
  nnd2s1 U4433 ( .Q(n3603), .DIN1(n3492), .DIN2(g266) );
  nnd2s1 U4434 ( .Q(n3602), .DIN1(n3487), .DIN2(g290) );
  nnd4s1 U4435 ( .Q(n3584), .DIN1(n3608), .DIN2(n3609), .DIN3(n3610), .DIN4(
        n3611) );
  and3s1 U4436 ( .Q(n3611), .DIN1(n3612), .DIN2(n3613), .DIN3(n3614) );
  nnd2s1 U4437 ( .Q(n3614), .DIN1(n3474), .DIN2(g1571) );
  nnd2s1 U4438 ( .Q(n3613), .DIN1(g901), .DIN2(n3473) );
  nnd2s1 U4439 ( .Q(n3612), .DIN1(n3554), .DIN2(g1341) );
  nnd2s1 U4440 ( .Q(n3610), .DIN1(n3494), .DIN2(g1552) );
  nnd2s1 U4441 ( .Q(n3609), .DIN1(n3472), .DIN2(g1595) );
  nnd2s1 U4442 ( .Q(n3608), .DIN1(n3493), .DIN2(g1528) );
  nnd2s1 U4443 ( .Q(g10402), .DIN1(n3437), .DIN2(n3189) );
  nor4s1 U4444 ( .Q(n3189), .DIN1(n3615), .DIN2(n3616), .DIN3(n3617), .DIN4(
        n3618) );
  nnd4s1 U4445 ( .Q(n3618), .DIN1(n3619), .DIN2(n3620), .DIN3(n3621), .DIN4(
        n3622) );
  and3s1 U4446 ( .Q(n3622), .DIN1(n3623), .DIN2(n3624), .DIN3(n3625) );
  nnd2s1 U4447 ( .Q(n3625), .DIN1(g1314), .DIN2(n3481) );
  nnd2s1 U4448 ( .Q(n3624), .DIN1(g886), .DIN2(n3539) );
  hi1s1 U4449 ( .Q(n3539), .DIN(n3626) );
  nnd2s1 U4450 ( .Q(n3623), .DIN1(n3538), .DIN2(g928) );
  hi1s1 U4451 ( .Q(n3538), .DIN(n3594) );
  nnd2s1 U4452 ( .Q(n3621), .DIN1(n3530), .DIN2(g971) );
  nnd2s1 U4453 ( .Q(n3620), .DIN1(g1170), .DIN2(n3482) );
  nnd2s1 U4454 ( .Q(n3619), .DIN1(g950), .DIN2(n3483) );
  nnd4s1 U4455 ( .Q(n3617), .DIN1(n3532), .DIN2(n3480), .DIN3(n3627), .DIN4(
        n3628) );
  and3s1 U4456 ( .Q(n3628), .DIN1(n3629), .DIN2(n3630), .DIN3(n3631) );
  nnd2s1 U4457 ( .Q(n3631), .DIN1(n3513), .DIN2(g119) );
  hi1s1 U4458 ( .Q(n3513), .DIN(n3512) );
  nnd2s1 U4459 ( .Q(n3630), .DIN1(g1194), .DIN2(n3540) );
  hi1s1 U4460 ( .Q(n3540), .DIN(n3632) );
  nnd2s1 U4461 ( .Q(n3629), .DIN1(n3514), .DIN2(g123) );
  hi1s1 U4462 ( .Q(n3514), .DIN(n3511) );
  nnd2s1 U4463 ( .Q(n3627), .DIN1(g922), .DIN2(n3601) );
  hi1s1 U4464 ( .Q(n3601), .DIN(n3633) );
  nnd4s1 U4465 ( .Q(n3532), .DIN1(n3632), .DIN2(n3511), .DIN3(n3479), .DIN4(
        n3634) );
  and3s1 U4466 ( .Q(n3634), .DIN1(n3480), .DIN2(n3583), .DIN3(n3512) );
  nnd2s1 U4467 ( .Q(n3512), .DIN1(n3635), .DIN2(n2125) );
  nnd2s1 U4468 ( .Q(n3511), .DIN1(n3635), .DIN2(g42) );
  and4s1 U4469 ( .Q(n3635), .DIN1(n3636), .DIN2(g43), .DIN3(n2130), .DIN4(
        n2128) );
  hi1s1 U4470 ( .Q(n2130), .DIN(g44) );
  nnd2s1 U4471 ( .Q(n3632), .DIN1(n3637), .DIN2(n3638) );
  nnd4s1 U4472 ( .Q(n3616), .DIN1(n3639), .DIN2(n3640), .DIN3(n3641), .DIN4(
        n3642) );
  nor2s1 U4473 ( .Q(n3642), .DIN1(n3643), .DIN2(n3644) );
  nor2s1 U4474 ( .Q(n3644), .DIN1(n3547), .DIN2(\DFF_168/net455 ) );
  and2s1 U4475 ( .Q(n3643), .DIN1(g1744), .DIN2(n3488) );
  nnd2s1 U4476 ( .Q(n3641), .DIN1(g1721), .DIN2(n3519) );
  nnd2s1 U4477 ( .Q(n3640), .DIN1(n3492), .DIN2(g263) );
  nnd2s1 U4478 ( .Q(n3639), .DIN1(n3487), .DIN2(g287) );
  hi1s1 U4479 ( .Q(n3487), .DIN(n3645) );
  nnd4s1 U4480 ( .Q(n3615), .DIN1(n3646), .DIN2(n3647), .DIN3(n3648), .DIN4(
        n3649) );
  and3s1 U4481 ( .Q(n3649), .DIN1(n3650), .DIN2(n3651), .DIN3(n3652) );
  nnd2s1 U4482 ( .Q(n3652), .DIN1(n3474), .DIN2(g1567) );
  nnd2s1 U4483 ( .Q(n3651), .DIN1(g898), .DIN2(n3473) );
  nnd2s1 U4484 ( .Q(n3650), .DIN1(n3554), .DIN2(g1336) );
  nnd2s1 U4485 ( .Q(n3648), .DIN1(n3494), .DIN2(g1549) );
  hi1s1 U4486 ( .Q(n3494), .DIN(n3653) );
  nnd2s1 U4487 ( .Q(n3647), .DIN1(n3472), .DIN2(g1592) );
  hi1s1 U4488 ( .Q(n3472), .DIN(n3654) );
  nnd2s1 U4489 ( .Q(n3646), .DIN1(n3493), .DIN2(g1524) );
  nnd2s1 U4490 ( .Q(g10339), .DIN1(n3437), .DIN2(n3310) );
  nor4s1 U4491 ( .Q(n3310), .DIN1(n3655), .DIN2(n3656), .DIN3(n3657), .DIN4(
        n3658) );
  nnd4s1 U4492 ( .Q(n3658), .DIN1(n3659), .DIN2(n3660), .DIN3(n3661), .DIN4(
        n3662) );
  nor2s1 U4493 ( .Q(n3662), .DIN1(n3663), .DIN2(n3664) );
  and2s1 U4494 ( .Q(n3664), .DIN1(n3554), .DIN2(g1311) );
  nor2s1 U4495 ( .Q(n3663), .DIN1(n3547), .DIN2(\DFF_319/net606 ) );
  nnd2s1 U4496 ( .Q(n3661), .DIN1(n3519), .DIN2(g1741) );
  nnd4s1 U4497 ( .Q(n3660), .DIN1(n3665), .DIN2(n3480), .DIN3(n3666), .DIN4(
        n3667) );
  nor2s1 U4498 ( .Q(n3666), .DIN1(n3554), .DIN2(n3519) );
  nnd4s1 U4499 ( .Q(n3480), .DIN1(n3637), .DIN2(n3668), .DIN3(g46), .DIN4(g47)
         );
  nnd2s1 U4500 ( .Q(n3659), .DIN1(g1191), .DIN2(n3482) );
  nnd3s1 U4501 ( .Q(n3657), .DIN1(n3669), .DIN2(n3670), .DIN3(n3671) );
  nnd2s1 U4502 ( .Q(n3671), .DIN1(n3474), .DIN2(g1589) );
  nnd2s1 U4503 ( .Q(n3670), .DIN1(g947), .DIN2(n3530) );
  nnd2s1 U4504 ( .Q(n3669), .DIN1(g919), .DIN2(n3473) );
  and2s1 U4505 ( .Q(n3656), .DIN1(g284), .DIN2(n3492) );
  and2s1 U4506 ( .Q(n3655), .DIN1(g1546), .DIN2(n3493) );
  nnd2s1 U4507 ( .Q(g10336), .DIN1(n3437), .DIN2(n3293) );
  hi1s1 U4508 ( .Q(n3293), .DIN(g10774) );
  or3s1 U4509 ( .Q(g10774), .DIN1(n3672), .DIN2(n3673), .DIN3(n3674) );
  nnd4s1 U4510 ( .Q(n3674), .DIN1(n3675), .DIN2(n3676), .DIN3(n3677), .DIN4(
        n3678) );
  and3s1 U4511 ( .Q(n3678), .DIN1(n3679), .DIN2(n3680), .DIN3(n3681) );
  nnd2s1 U4512 ( .Q(n3681), .DIN1(n3474), .DIN2(g1586) );
  and2s1 U4513 ( .Q(n3474), .DIN1(n3636), .DIN2(n3682) );
  nnd2s1 U4514 ( .Q(n3680), .DIN1(g944), .DIN2(n3530) );
  hi1s1 U4515 ( .Q(n3530), .DIN(n3683) );
  nnd2s1 U4516 ( .Q(n3679), .DIN1(g916), .DIN2(n3473) );
  hi1s1 U4517 ( .Q(n3473), .DIN(n3684) );
  nnd2s1 U4518 ( .Q(n3677), .DIN1(g968), .DIN2(n3483) );
  hi1s1 U4519 ( .Q(n3483), .DIN(n3685) );
  nnd2s1 U4520 ( .Q(n3676), .DIN1(g1333), .DIN2(n3481) );
  hi1s1 U4521 ( .Q(n3481), .DIN(n3686) );
  nnd2s1 U4522 ( .Q(n3675), .DIN1(g1188), .DIN2(n3482) );
  nnd4s1 U4523 ( .Q(n3673), .DIN1(n3687), .DIN2(n3688), .DIN3(n3689), .DIN4(
        n3690) );
  nnd2s1 U4524 ( .Q(n3690), .DIN1(n3479), .DIN2(n3583) );
  and4s1 U4525 ( .Q(n3479), .DIN1(n3665), .DIN2(n3686), .DIN3(n3691), .DIN4(
        n3692) );
  nor2s1 U4526 ( .Q(n3691), .DIN1(n3482), .DIN2(n3488) );
  hi1s1 U4527 ( .Q(n3482), .DIN(n3667) );
  nnd2s1 U4528 ( .Q(n3667), .DIN1(n3693), .DIN2(n3638) );
  nnd2s1 U4529 ( .Q(n3686), .DIN1(n3638), .DIN2(n3694) );
  nor4s1 U4530 ( .Q(n3665), .DIN1(n3695), .DIN2(n3696), .DIN3(n3697), .DIN4(
        n3698) );
  nnd4s1 U4531 ( .Q(n3698), .DIN1(n3684), .DIN2(n3654), .DIN3(n3683), .DIN4(
        n3699) );
  and3s1 U4532 ( .Q(n3699), .DIN1(n3626), .DIN2(n3594), .DIN3(n3633) );
  nnd2s1 U4533 ( .Q(n3633), .DIN1(n3637), .DIN2(n3700) );
  nnd4s1 U4534 ( .Q(n3594), .DIN1(n3700), .DIN2(g44), .DIN3(g45), .DIN4(n3294)
         );
  nnd4s1 U4535 ( .Q(n3626), .DIN1(n3700), .DIN2(g43), .DIN3(n3701), .DIN4(g42)
         );
  nnd2s1 U4536 ( .Q(n3683), .DIN1(n3682), .DIN2(n3700) );
  nnd2s1 U4537 ( .Q(n3654), .DIN1(n3636), .DIN2(n3694) );
  nnd2s1 U4538 ( .Q(n3684), .DIN1(n3700), .DIN2(n3693) );
  nnd3s1 U4539 ( .Q(n3697), .DIN1(n3702), .DIN2(n3685), .DIN3(n3547) );
  nnd2s1 U4540 ( .Q(n3685), .DIN1(n3700), .DIN2(n3694) );
  and3s1 U4541 ( .Q(n3694), .DIN1(n2125), .DIN2(n2126), .DIN3(n3701) );
  and3s1 U4542 ( .Q(n3700), .DIN1(g46), .DIN2(n2124), .DIN3(n3668) );
  nnd2s1 U4543 ( .Q(n3702), .DIN1(n3636), .DIN2(n3682) );
  nnd2s1 U4544 ( .Q(n3689), .DIN1(g1308), .DIN2(n3554) );
  hi1s1 U4545 ( .Q(n3554), .DIN(n3583) );
  nnd2s1 U4546 ( .Q(n3583), .DIN1(n3682), .DIN2(n3638) );
  and2s1 U4547 ( .Q(n3682), .DIN1(n3701), .DIN2(n3294) );
  nor2s1 U4548 ( .Q(n3701), .DIN1(n2128), .DIN2(g44) );
  nnd2s1 U4549 ( .Q(n3688), .DIN1(n3488), .DIN2(g1762) );
  and2s1 U4550 ( .Q(n3488), .DIN1(n3703), .DIN2(n2125) );
  nnd2s1 U4551 ( .Q(n3687), .DIN1(g39), .DIN2(n3442) );
  nnd3s1 U4552 ( .Q(n3672), .DIN1(n3704), .DIN2(n3705), .DIN3(n3706) );
  nnd2s1 U4553 ( .Q(n3706), .DIN1(n3519), .DIN2(g1738) );
  hi1s1 U4554 ( .Q(n3519), .DIN(n3692) );
  nnd2s1 U4555 ( .Q(n3692), .DIN1(n3703), .DIN2(g42) );
  and4s1 U4556 ( .Q(n3703), .DIN1(g44), .DIN2(g43), .DIN3(n3638), .DIN4(g45)
         );
  and3s1 U4557 ( .Q(n3638), .DIN1(g47), .DIN2(n2121), .DIN3(n3668) );
  nnd2s1 U4558 ( .Q(n3705), .DIN1(n3493), .DIN2(g1543) );
  and2s1 U4559 ( .Q(n3493), .DIN1(n3695), .DIN2(n3653) );
  nnd2s1 U4560 ( .Q(n3695), .DIN1(n3653), .DIN2(n3707) );
  nnd2s1 U4561 ( .Q(n3707), .DIN1(n3636), .DIN2(n3693) );
  and4s1 U4562 ( .Q(n3693), .DIN1(g44), .DIN2(g43), .DIN3(g42), .DIN4(n2128)
         );
  nnd2s1 U4563 ( .Q(n3653), .DIN1(n3637), .DIN2(n3636) );
  and2s1 U4564 ( .Q(n3637), .DIN1(n3708), .DIN2(g43) );
  nnd2s1 U4565 ( .Q(n3704), .DIN1(n3492), .DIN2(g281) );
  and2s1 U4566 ( .Q(n3492), .DIN1(n3696), .DIN2(n3645) );
  nnd2s1 U4567 ( .Q(n3696), .DIN1(n3645), .DIN2(n3709) );
  nnd4s1 U4568 ( .Q(n3709), .DIN1(n3636), .DIN2(g44), .DIN3(n3294), .DIN4(
        n2128) );
  nor2s1 U4569 ( .Q(n3294), .DIN1(n2125), .DIN2(g43) );
  nnd3s1 U4570 ( .Q(n3645), .DIN1(n3636), .DIN2(n2126), .DIN3(n3708) );
  and3s1 U4571 ( .Q(n3708), .DIN1(n2125), .DIN2(n2128), .DIN3(g44) );
  hi1s1 U4572 ( .Q(n2128), .DIN(g45) );
  hi1s1 U4573 ( .Q(n2125), .DIN(g42) );
  hi1s1 U4574 ( .Q(n2126), .DIN(g43) );
  and3s1 U4575 ( .Q(n3636), .DIN1(n2121), .DIN2(n2124), .DIN3(n3668) );
  and2s1 U4576 ( .Q(n3668), .DIN1(n3710), .DIN2(n2081) );
  nnd2s1 U4577 ( .Q(n2081), .DIN1(n3711), .DIN2(n3712) );
  or3s1 U4578 ( .Q(n3712), .DIN1(g41), .DIN2(g48), .DIN3(g30) );
  nnd2s1 U4579 ( .Q(n3711), .DIN1(n3547), .DIN2(n3710) );
  nor2s1 U4580 ( .Q(n3710), .DIN1(n2129), .DIN2(g41) );
  hi1s1 U4581 ( .Q(n2124), .DIN(g47) );
  hi1s1 U4582 ( .Q(n2121), .DIN(g46) );
  nor2s1 U4583 ( .Q(n3437), .DIN1(n3442), .DIN2(g30) );
  hi1s1 U4584 ( .Q(n3442), .DIN(n3547) );
  nor2s1 U4585 ( .Q(n3547), .DIN1(n2129), .DIN2(g31) );
  hi1s1 U4586 ( .Q(n2129), .DIN(g48) );
  dffs1 \DFF_533/Q_reg  ( .QN(n2034), .Q(g8816), .CLK(CK), .DIN(g7784) );
  dffs1 \DFF_532/Q_reg  ( .Q(g1878), .CLK(CK), .DIN(g8695) );
  dffs1 \DFF_531/Q_reg  ( .Q(g12), .CLK(CK), .DIN(g7337) );
  dffs1 \DFF_530/Q_reg  ( .Q(g1724), .CLK(CK), .DIN(g10879) );
  dffs1 \DFF_529/Q_reg  ( .Q(g511), .CLK(CK), .DIN(g11336) );
  dffs1 \DFF_528/Q_reg  ( .Q(g1), .CLK(CK), .DIN(g8078) );
  dffs1 \DFF_526/Q_reg  ( .Q(g1360), .CLK(CK), .DIN(g9824) );
  dffs1 \DFF_525/Q_reg  ( .QN(n1966), .CLK(CK), .DIN(g6302) );
  dffs1 \DFF_524/Q_reg  ( .Q(g569), .CLK(CK), .DIN(g10876) );
  dffs1 \DFF_523/Q_reg  ( .Q(g1776), .CLK(CK), .DIN(g7812) );
  dffs1 \DFF_522/Q_reg  ( .Q(g534), .CLK(CK), .DIN(g11327) );
  dffs1 \DFF_521/Q_reg  ( .Q(g691), .CLK(CK), .DIN(g8430) );
  dffs1 \DFF_520/Q_reg  ( .Q(g1567), .CLK(CK), .DIN(g7352) );
  dffs1 \DFF_519/Q_reg  ( .Q(g1494), .CLK(CK), .DIN(g8446) );
  dffs1 \DFF_518/Q_reg  ( .Q(g643), .CLK(CK), .DIN(g8064) );
  dffs1 \DFF_517/Q_reg  ( .QN(n1934), .CLK(CK), .DIN(g6313) );
  dffs1 \DFF_516/Q_reg  ( .Q(g1621), .CLK(CK), .DIN(g8869) );
  dffs1 \DFF_515/Q_reg  ( .Q(g995), .CLK(CK), .DIN(g7801) );
  dffs1 \DFF_514/Q_reg  ( .Q(g1555), .CLK(CK), .DIN(g7348) );
  dffs1 \DFF_513/Q_reg  ( .QN(n2019), .Q(g8813), .CLK(CK), .DIN(g7781) );
  dffs1 \DFF_512/Q_reg  ( .QN(n2033), .Q(g435), .CLK(CK), .DIN(g11261) );
  dffs1 \DFF_511/Q_reg  ( .Q(g299), .CLK(CK), .DIN(g7772) );
  dffs1 \DFF_510/Q_reg  ( .Q(g1235), .CLK(CK), .DIN(g7296) );
  dffs1 \DFF_509/Q_reg  ( .Q(g1618), .CLK(CK), .DIN(g11611) );
  dffs1 \DFF_508/Q_reg  ( .QN(n1960), .Q(g127), .CLK(CK), .DIN(g8421) );
  dffs1 \DFF_507/Q_reg  ( .QN(n1943), .CLK(CK), .DIN(g11181) );
  dffs1 \DFF_506/Q_reg  ( .Q(g1351), .CLK(CK), .DIN(g11657) );
  dffs1 \DFF_505/Q_reg  ( .Q(g1528), .CLK(CK), .DIN(g7339) );
  dffs1 \DFF_504/Q_reg  ( .Q(g1666), .CLK(CK), .DIN(g11035) );
  dffs1 \DFF_503/Q_reg  ( .Q(g1440), .CLK(CK), .DIN(g8988) );
  dffs1 \DFF_502/Q_reg  ( .Q(g585), .CLK(CK), .DIN(g6293) );
  dffs1 \DFF_501/Q_reg  ( .Q(g1750), .CLK(CK), .DIN(g5665) );
  dffs1 \DFF_500/Q_reg  ( .Q(g5645), .CLK(CK), .DIN(g7752) );
  dffs1 \DFF_499/Q_reg  ( .Q(g339), .CLK(CK), .DIN(g11505) );
  dffs1 \DFF_498/Q_reg  ( .Q(g1300), .CLK(CK), .DIN(g7291) );
  dffs1 \DFF_497/Q_reg  ( .Q(g991), .CLK(CK), .DIN(g7802) );
  dffs1 \DFF_496/Q_reg  ( .QN(n2038), .Q(g8817), .CLK(CK), .DIN(g7774) );
  dffs1 \DFF_495/Q_reg  ( .Q(g1630), .CLK(CK), .DIN(g8872) );
  dffs1 \DFF_494/Q_reg  ( .Q(g1515), .CLK(CK), .DIN(g7333) );
  dffs1 \DFF_493/Q_reg  ( .Q(g1905), .CLK(CK), .DIN(g8283) );
  dffs1 \DFF_492/Q_reg  ( .QN(n2054), .Q(g431), .CLK(CK), .DIN(g11262) );
  dffs1 \DFF_491/Q_reg  ( .Q(g411), .CLK(CK), .DIN(g11268) );
  dffs1 \DFF_490/Q_reg  ( .QN(n1959), .Q(g162), .CLK(CK), .DIN(g8424) );
  dffs1 \DFF_489/Q_reg  ( .QN(\DFF_489/net776 ), .CLK(CK), .DIN(g5672) );
  dffs1 \DFF_488/Q_reg  ( .Q(g673), .CLK(CK), .DIN(g8428) );
  dffs1 \DFF_487/Q_reg  ( .QN(n2004), .CLK(CK), .DIN(g7314) );
  dffs1 \DFF_486/Q_reg  ( .QN(n2031), .Q(g1284), .CLK(CK), .DIN(g7294) );
  dffs1 \DFF_485/Q_reg  ( .Q(g266), .CLK(CK), .DIN(g7761) );
  dffs1 \DFF_484/Q_reg  ( .QN(n1965), .CLK(CK), .DIN(g6825) );
  dffs1 \DFF_483/Q_reg  ( .Q(g382), .CLK(CK), .DIN(g11442) );
  dffs1 \DFF_482/Q_reg  ( .Q(g1615), .CLK(CK), .DIN(g8868) );
  dffs1 \DFF_481/Q_reg  ( .Q(g1311), .CLK(CK), .DIN(g11628) );
  dffs1 \DFF_480/Q_reg  ( .Q(g1275), .CLK(CK), .DIN(g11443) );
  dffs1 \DFF_479/Q_reg  ( .QN(n2035), .Q(g8814), .CLK(CK), .DIN(g7782) );
  dffs1 \DFF_478/Q_reg  ( .Q(g321), .CLK(CK), .DIN(g5647) );
  dffs1 \DFF_477/Q_reg  ( .Q(g1607), .CLK(CK), .DIN(g7365) );
  dffs1 \DFF_476/Q_reg  ( .Q(g581), .CLK(CK), .DIN(g6295) );
  dffs1 \DFF_475/Q_reg  ( .QN(n2032), .Q(g525), .CLK(CK), .DIN(g11329) );
  dffs1 \DFF_474/Q_reg  ( .QN(n1961), .Q(g135), .CLK(CK), .DIN(g8419) );
  dffs1 \DFF_473/Q_reg  ( .QN(n2042), .CLK(CK), .DIN(g7321) );
  dffs1 \DFF_472/Q_reg  ( .QN(n1967), .CLK(CK), .DIN(g11184) );
  dffs1 \DFF_471/Q_reg  ( .Q(g1710), .CLK(CK), .DIN(g4901) );
  dffs1 \DFF_470/Q_reg  ( .Q(g1341), .CLK(CK), .DIN(g11655) );
  dffs1 \DFF_468/Q_reg  ( .QN(n1944), .Q(g1141), .CLK(CK), .DIN(g6311) );
  dffs1 \DFF_467/Q_reg  ( .Q(g324), .CLK(CK), .DIN(g5648) );
  dffs1 \DFF_466/Q_reg  ( .Q(g1586), .CLK(CK), .DIN(g7358) );
  dffs1 \DFF_465/Q_reg  ( .Q(g1687), .CLK(CK), .DIN(g11042) );
  dffs1 \DFF_464/Q_reg  ( .Q(g584), .CLK(CK), .DIN(g6292) );
  dffs1 \DFF_463/Q_reg  ( .Q(g1552), .CLK(CK), .DIN(g7347) );
  dffs1 \DFF_462/Q_reg  ( .Q(g755), .CLK(CK), .DIN(g6338) );
  dffs1 \DFF_461/Q_reg  ( .QN(n1957), .Q(g1909), .CLK(CK), .DIN(g9352) );
  dffs1 \DFF_460/Q_reg  ( .Q(g546), .CLK(CK), .DIN(g11043) );
  dffs1 \DFF_459/Q_reg  ( .Q(g506), .CLK(CK), .DIN(g11335) );
  dffs1 \DFF_458/Q_reg  ( .Q(g1321), .CLK(CK), .DIN(g11631) );
  dffs1 \DFF_457/Q_reg  ( .QN(n2015), .Q(g1121), .CLK(CK), .DIN(g6306) );
  dffs1 \DFF_456/Q_reg  ( .Q(g1598), .CLK(CK), .DIN(g7362) );
  dffs1 \DFF_455/Q_reg  ( .QN(n1948), .Q(g1834), .CLK(CK), .DIN(g9895) );
  dffs1 \DFF_454/Q_reg  ( .Q(g947), .CLK(CK), .DIN(g11399) );
  dffs1 \DFF_453/Q_reg  ( .Q(g1549), .CLK(CK), .DIN(g7346) );
  dffs1 \DFF_452/Q_reg  ( .QN(\DFF_452/net739 ), .CLK(CK), .DIN(g7320) );
  dffs1 \DFF_451/Q_reg  ( .Q(g582), .CLK(CK), .DIN(g6296) );
  dffs1 \DFF_450/Q_reg  ( .QN(n1968), .Q(g677), .CLK(CK), .DIN(g9341) );
  dffs1 \DFF_449/Q_reg  ( .QN(n1956), .Q(g1872), .CLK(CK), .DIN(g9348) );
  dffs1 \DFF_448/Q_reg  ( .Q(g1318), .CLK(CK), .DIN(g11630) );
  dffs1 \DFF_447/Q_reg  ( .QN(n2053), .Q(g521), .CLK(CK), .DIN(g11330) );
  dffs1 \DFF_446/Q_reg  ( .Q(g5647), .CLK(CK), .DIN(g7754) );
  dffs1 \DFF_445/Q_reg  ( .Q(g7), .CLK(CK), .DIN(g2731) );
  dffs1 \DFF_444/Q_reg  ( .QN(n1996), .Q(g131), .CLK(CK), .DIN(g8420) );
  dffs1 \DFF_443/Q_reg  ( .Q(g5649), .CLK(CK), .DIN(g7756) );
  dffs1 \DFF_442/Q_reg  ( .Q(g1260), .CLK(CK), .DIN(g7301) );
  dffs1 \DFF_441/Q_reg  ( .QN(\DFF_441/net728 ), .CLK(CK), .DIN(g874) );
  dffs1 \DFF_440/Q_reg  ( .Q(g348), .CLK(CK), .DIN(g11506) );
  dffs1 \DFF_438/Q_reg  ( .QN(n1927), .CLK(CK), .DIN(g6300) );
  dffs1 \DFF_437/Q_reg  ( .Q(g1490), .CLK(CK), .DIN(g8445) );
  dffs1 \DFF_436/Q_reg  ( .QN(\DFF_436/net723 ), .CLK(CK), .DIN(g113) );
  dffs1 \DFF_435/Q_reg  ( .Q(g1512), .CLK(CK), .DIN(g8449) );
  dffs1 \DFF_434/Q_reg  ( .QN(n2055), .Q(g790), .CLK(CK), .DIN(g8567) );
  dffs1 \DFF_433/Q_reg  ( .Q(g845), .CLK(CK), .DIN(g4186) );
  dffs1 \DFF_432/Q_reg  ( .Q(g1330), .CLK(CK), .DIN(g11634) );
  dffs1 \DFF_431/Q_reg  ( .Q(g754), .CLK(CK), .DIN(g4895) );
  dffs1 \DFF_430/Q_reg  ( .Q(g481), .CLK(CK), .DIN(g11324) );
  dffs1 \DFF_429/Q_reg  ( .QN(n1990), .Q(g4183), .CLK(CK), .DIN(g6801) );
  dffs1 \DFF_428/Q_reg  ( .Q(g999), .CLK(CK), .DIN(g7804) );
  dffs1 \DFF_427/Q_reg  ( .Q(g727), .CLK(CK), .DIN(g8434) );
  dffs1 \DFF_426/Q_reg  ( .Q(g1537), .CLK(CK), .DIN(g7342) );
  dffs1 \DFF_425/Q_reg  ( .Q(g1595), .CLK(CK), .DIN(g7361) );
  dffs1 \DFF_424/Q_reg  ( .QN(n1931), .CLK(CK), .DIN(g6835) );
  dffs1 \DFF_423/Q_reg  ( .Q(g1654), .CLK(CK), .DIN(g10874) );
  dffs1 \DFF_421/Q_reg  ( .QN(n2006), .CLK(CK), .DIN(g11183) );
  dffs1 \DFF_420/Q_reg  ( .Q(g1811), .CLK(CK), .DIN(g11185) );
  dffs1 \DFF_419/Q_reg  ( .Q(g406), .CLK(CK), .DIN(g11267) );
  dffs1 \DFF_418/Q_reg  ( .Q(g1223), .CLK(CK), .DIN(g8277) );
  dffs1 \DFF_417/Q_reg  ( .QN(n1929), .Q(g1107), .CLK(CK), .DIN(g6816) );
  dffs1 \DFF_416/Q_reg  ( .QN(n1970), .Q(g1145), .CLK(CK), .DIN(g6312) );
  dffs1 \DFF_415/Q_reg  ( .Q(g1403), .CLK(CK), .DIN(g8991) );
  dffs1 \DFF_414/Q_reg  ( .Q(g1003), .CLK(CK), .DIN(g7803) );
  dffs1 \DFF_413/Q_reg  ( .Q(g1027), .CLK(CK), .DIN(g7798) );
  dffs1 \DFF_412/Q_reg  ( .Q(g841), .CLK(CK), .DIN(g4185) );
  dffs1 \DFF_411/Q_reg  ( .Q(g589), .CLK(CK), .DIN(g6297) );
  dffs1 \DFF_410/Q_reg  ( .Q(g1756), .CLK(CK), .DIN(g5667) );
  dffs1 \DFF_409/Q_reg  ( .Q(g378), .CLK(CK), .DIN(g11441) );
  dffs1 \DFF_408/Q_reg  ( .Q(g956), .CLK(CK), .DIN(g11402) );
  dffs1 \DFF_407/Q_reg  ( .QN(n2051), .Q(g762), .CLK(CK), .DIN(g6798) );
  dffs1 \DFF_406/Q_reg  ( .Q(g421), .CLK(CK), .DIN(g11270) );
  dffs1 \DFF_405/Q_reg  ( .Q(g853), .CLK(CK), .DIN(g4188) );
  dffs1 \DFF_404/Q_reg  ( .Q(g1636), .CLK(CK), .DIN(g8874) );
  dffs1 \DFF_403/Q_reg  ( .QN(n2026), .CLK(CK), .DIN(g8066) );
  dffs1 \DFF_402/Q_reg  ( .Q(g1083), .CLK(CK), .DIN(g6807) );
  dffs1 \DFF_401/Q_reg  ( .QN(n2052), .Q(g1280), .CLK(CK), .DIN(g7295) );
  dffs1 \DFF_400/Q_reg  ( .QN(n1995), .Q(g201), .CLK(CK), .DIN(g7304) );
  dffs1 \DFF_399/Q_reg  ( .QN(n2014), .Q(g1125), .CLK(CK), .DIN(g6307) );
  dffs1 \DFF_398/Q_reg  ( .Q(g875), .CLK(CK), .DIN(g9822) );
  dffs1 \DFF_397/Q_reg  ( .Q(g5643), .CLK(CK), .DIN(g7750) );
  dffs1 \DFF_396/Q_reg  ( .Q(g1386), .CLK(CK), .DIN(g7318) );
  dffs1 \DFF_395/Q_reg  ( .QN(n2039), .Q(g658), .CLK(CK), .DIN(g9339) );
  dffs1 \DFF_394/Q_reg  ( .Q(g391), .CLK(CK), .DIN(g11264) );
  dffs1 \DFF_393/Q_reg  ( .QN(n2050), .Q(g4186), .CLK(CK), .DIN(g7786) );
  dffs1 \DFF_392/Q_reg  ( .Q(g1577), .CLK(CK), .DIN(g7355) );
  dffs1 \DFF_391/Q_reg  ( .Q(g1524), .CLK(CK), .DIN(g7338) );
  dffs1 \DFF_390/Q_reg  ( .Q(g275), .CLK(CK), .DIN(g7764) );
  dffs1 \DFF_389/Q_reg  ( .QN(n1999), .Q(g4184), .CLK(CK), .DIN(g6802) );
  dffs1 \DFF_388/Q_reg  ( .Q(g1747), .CLK(CK), .DIN(g5664) );
  dffs1 \DFF_387/Q_reg  ( .QN(n2049), .Q(g4188), .CLK(CK), .DIN(g8274) );
  dffs1 \DFF_386/Q_reg  ( .Q(g263), .CLK(CK), .DIN(g7760) );
  dffs1 \DFF_385/Q_reg  ( .QN(\DFF_385/net672 ), .CLK(CK), .DIN(g7366) );
  dffs1 \DFF_384/Q_reg  ( .QN(\DFF_384/net671 ), .CLK(CK), .DIN(g10868) );
  dffs1 \DFF_383/Q_reg  ( .QN(n2016), .Q(g1149), .CLK(CK), .DIN(g6305) );
  dffs1 \DFF_382/Q_reg  ( .QN(n1938), .Q(g139), .CLK(CK), .DIN(g8418) );
  dffs1 \DFF_381/Q_reg  ( .QN(n1936), .Q(g668), .CLK(CK), .DIN(g9340) );
  dffs1 \DFF_380/Q_reg  ( .QN(n2017), .Q(g119), .CLK(CK), .DIN(g7745) );
  dffs1 \DFF_379/Q_reg  ( .Q(g476), .CLK(CK), .DIN(g11338) );
  dffs1 \DFF_378/Q_reg  ( .Q(g440), .CLK(CK), .DIN(g11260) );
  dffs1 \DFF_377/Q_reg  ( .Q(g578), .CLK(CK), .DIN(g6292) );
  dffs1 \DFF_376/Q_reg  ( .Q(g1068), .CLK(CK), .DIN(g6803) );
  dffs1 \DFF_374/Q_reg  ( .Q(g1624), .CLK(CK), .DIN(g8870) );
  dffs1 \DFF_373/Q_reg  ( .Q(g1932), .CLK(CK), .DIN(g8286) );
  dffs1 \DFF_372/Q_reg  ( .Q(g1703), .CLK(CK), .DIN(g6843) );
  dffs1 \DFF_371/Q_reg  ( .Q(g1592), .CLK(CK), .DIN(g7360) );
  dffs1 \DFF_370/Q_reg  ( .Q(g1727), .CLK(CK), .DIN(g10880) );
  dffs1 \DFF_369/Q_reg  ( .QN(n1980), .Q(g1828), .CLK(CK), .DIN(g9827) );
  dffs1 \DFF_368/Q_reg  ( .Q(g448), .CLK(CK), .DIN(g11258) );
  dffs1 \DFF_367/Q_reg  ( .Q(g857), .CLK(CK), .DIN(g4189) );
  dffs1 \DFF_366/Q_reg  ( .QN(n1945), .Q(g1129), .CLK(CK), .DIN(g6308) );
  dffs1 \DFF_365/Q_reg  ( .Q(g950), .CLK(CK), .DIN(g11400) );
  dffs1 \DFF_364/Q_reg  ( .Q(g182), .CLK(CK), .DIN(g7749) );
  dffs1 \DFF_363/Q_reg  ( .QN(n2022), .Q(g8819), .CLK(CK), .DIN(g7776) );
  dffs1 \DFF_362/Q_reg  ( .QN(n1978), .Q(g605), .CLK(CK), .DIN(g9820) );
  dffs1 \DFF_361/Q_reg  ( .Q(g1218), .CLK(CK), .DIN(g8276) );
  dffs1 \DFF_360/Q_reg  ( .Q(g2613), .CLK(CK), .DIN(g8781) );
  dffs1 \DFF_359/Q_reg  ( .QN(n2009), .Q(g731), .CLK(CK), .DIN(g9347) );
  dffs1 \DFF_358/Q_reg  ( .QN(n1951), .Q(g591), .CLK(CK), .DIN(g9818) );
  dffs1 \DFF_357/Q_reg  ( .Q(g874), .CLK(CK), .DIN(g9821) );
  dffs1 \DFF_356/Q_reg  ( .Q(g5646), .CLK(CK), .DIN(g7753) );
  dffs1 \DFF_355/Q_reg  ( .Q(g1255), .CLK(CK), .DIN(g7300) );
  dffs1 \DFF_354/Q_reg  ( .QN(n2010), .Q(g1891), .CLK(CK), .DIN(g9350) );
  dffs1 \DFF_353/Q_reg  ( .QN(n2013), .Q(g1137), .CLK(CK), .DIN(g6310) );
  dffs1 \DFF_352/Q_reg  ( .QN(n1998), .CLK(CK), .DIN(g5673) );
  dffs1 \DFF_351/Q_reg  ( .Q(g968), .CLK(CK), .DIN(g11406) );
  dffs1 \DFF_350/Q_reg  ( .Q(g37), .CLK(CK), .DIN(g10871) );
  dffs1 \DFF_349/Q_reg  ( .Q(g1887), .CLK(CK), .DIN(g8281) );
  dffs1 \DFF_347/Q_reg  ( .Q(g4190), .CLK(CK), .DIN(g8568) );
  dffs1 \DFF_346/Q_reg  ( .Q(g1806), .CLK(CK), .DIN(g8573) );
  dffs1 \DFF_345/Q_reg  ( .Q(g272), .CLK(CK), .DIN(g7763) );
  dffs1 \DFF_344/Q_reg  ( .Q(g1336), .CLK(CK), .DIN(g11654) );
  dffs1 \DFF_343/Q_reg  ( .Q(g849), .CLK(CK), .DIN(g4187) );
  dffs1 \DFF_342/Q_reg  ( .Q(g1314), .CLK(CK), .DIN(g11629) );
  dffs1 \DFF_340/Q_reg  ( .QN(n2046), .Q(g936), .CLK(CK), .DIN(g8571) );
  dffs1 \DFF_339/Q_reg  ( .Q(g1923), .CLK(CK), .DIN(g8285) );
  dffs1 \DFF_338/Q_reg  ( .Q(g833), .CLK(CK), .DIN(g4183) );
  dffs1 \DFF_337/Q_reg  ( .QN(n1926), .Q(g148), .CLK(CK), .DIN(g8427) );
  dffs1 \DFF_336/Q_reg  ( .QN(\DFF_336/net623 ), .CLK(CK), .DIN(g7287) );
  dffs1 \DFF_335/Q_reg  ( .QN(n2011), .Q(g108), .CLK(CK), .DIN(g11593) );
  dffs1 \DFF_334/Q_reg  ( .Q(g1245), .CLK(CK), .DIN(g7298) );
  dffs1 \DFF_333/Q_reg  ( .QN(n1932), .Q(g1900), .CLK(CK), .DIN(g9351) );
  dffs1 \DFF_332/Q_reg  ( .QN(n1984), .Q(g1781), .CLK(CK), .DIN(g7813) );
  dffs1 \DFF_331/Q_reg  ( .QN(n1962), .Q(g213), .CLK(CK), .DIN(g7313) );
  dffs1 \DFF_330/Q_reg  ( .QN(\DFF_330/net617 ), .CLK(CK), .DIN(g5670) );
  dffs1 \DFF_329/Q_reg  ( .Q(g491), .CLK(CK), .DIN(g11332) );
  dffs1 \DFF_328/Q_reg  ( .Q(g3069), .CLK(CK), .DIN(g4898) );
  dffs1 \DFF_327/Q_reg  ( .QN(n1941), .CLK(CK), .DIN(g7312) );
  dffs1 \DFF_326/Q_reg  ( .Q(g1540), .CLK(CK), .DIN(g7343) );
  dffs1 \DFF_325/Q_reg  ( .Q(g1324), .CLK(CK), .DIN(g11632) );
  dffs1 \DFF_324/Q_reg  ( .QN(n1952), .Q(g1796), .CLK(CK), .DIN(g8280) );
  dffs1 \DFF_323/Q_reg  ( .Q(g1610), .CLK(CK), .DIN(g6845) );
  dffs1 \DFF_322/Q_reg  ( .Q(g1270), .CLK(CK), .DIN(g7303) );
  dffs1 \DFF_321/Q_reg  ( .Q(g1733), .CLK(CK), .DIN(g10882) );
  dffs1 \DFF_320/Q_reg  ( .Q(g1765), .CLK(CK), .DIN(g3329) );
  dffs1 \DFF_319/Q_reg  ( .QN(\DFF_319/net606 ), .CLK(CK), .DIN(g10775) );
  dffs1 \DFF_318/Q_reg  ( .Q(g2044), .CLK(CK), .DIN(g6339) );
  dffs1 \DFF_317/Q_reg  ( .Q(g953), .CLK(CK), .DIN(g11401) );
  dffs1 \DFF_316/Q_reg  ( .QN(n1933), .Q(g686), .CLK(CK), .DIN(g9342) );
  dffs1 \DFF_315/Q_reg  ( .Q(g1520), .CLK(CK), .DIN(g7334) );
  dffs1 \DFF_314/Q_reg  ( .Q(g170), .CLK(CK), .DIN(g8422) );
  dffs1 \DFF_313/Q_reg  ( .Q(g1941), .CLK(CK), .DIN(g8287) );
  dffs1 \DFF_312/Q_reg  ( .Q(g944), .CLK(CK), .DIN(g11398) );
  dffs1 \DFF_311/Q_reg  ( .Q(g2731), .CLK(CK), .DIN(g11408) );
  dffs1 \DFF_310/Q_reg  ( .QN(n1985), .Q(g599), .CLK(CK), .DIN(g9819) );
  dffs1 \DFF_309/Q_reg  ( .Q(g837), .CLK(CK), .DIN(g4184) );
  dffs1 \DFF_308/Q_reg  ( .Q(g366), .CLK(CK), .DIN(g11512) );
  dffs1 \DFF_307/Q_reg  ( .Q(g178), .CLK(CK), .DIN(g7748) );
  dffs1 \DFF_306/Q_reg  ( .Q(g1462), .CLK(CK), .DIN(g8438) );
  dffs1 \DFF_304/Q_reg  ( .Q(g2639), .CLK(CK), .DIN(g2638) );
  dffs1 \DFF_303/Q_reg  ( .QN(n1939), .Q(g237), .CLK(CK), .DIN(g7306) );
  dffs1 \DFF_302/Q_reg  ( .QN(n1953), .Q(g1822), .CLK(CK), .DIN(g9826) );
  dffs1 \DFF_301/Q_reg  ( .QN(n2056), .Q(g782), .CLK(CK), .DIN(g8273) );
  dffs1 \DFF_300/Q_reg  ( .QN(n2028), .Q(g1918), .CLK(CK), .DIN(g9353) );
  dffs1 \DFF_299/Q_reg  ( .Q(g1212), .CLK(CK), .DIN(g1217) );
  dffs1 \DFF_297/Q_reg  ( .QN(n1986), .Q(g1814), .CLK(CK), .DIN(g9825) );
  dffs1 \DFF_296/Q_reg  ( .QN(n1925), .Q(g143), .CLK(CK), .DIN(g7746) );
  dffs1 \DFF_295/Q_reg  ( .Q(g1955), .CLK(CK), .DIN(g6338) );
  dffs1 \DFF_294/Q_reg  ( .Q(g971), .CLK(CK), .DIN(g11470) );
  dffs1 \DFF_293/Q_reg  ( .Q(g986), .CLK(CK), .DIN(g11473) );
  dffs1 \DFF_292/Q_reg  ( .Q(g1071), .CLK(CK), .DIN(g6804) );
  dffs1 \DFF_291/Q_reg  ( .Q(g2986), .CLK(CK), .DIN(g4897) );
  dffs1 \DFF_290/Q_reg  ( .Q(g1089), .CLK(CK), .DIN(g6809) );
  dffs1 \DFF_289/Q_reg  ( .QN(n2024), .CLK(CK), .DIN(g7809) );
  dffs1 \DFF_288/Q_reg  ( .Q(g566), .CLK(CK), .DIN(g11051) );
  dffs1 \DFF_287/Q_reg  ( .QN(n2036), .Q(g8812), .CLK(CK), .DIN(g7780) );
  dffs1 \DFF_286/Q_reg  ( .QN(n1994), .Q(g722), .CLK(CK), .DIN(g9346) );
  dffs1 \DFF_285/Q_reg  ( .Q(g1657), .CLK(CK), .DIN(g10875) );
  dffs1 \DFF_284/Q_reg  ( .QN(n1946), .Q(g192), .CLK(CK), .DIN(g6837) );
  dffs1 \DFF_283/Q_reg  ( .Q(g360), .CLK(CK), .DIN(g11510) );
  dffs1 \DFF_282/Q_reg  ( .Q(g1762), .CLK(CK), .DIN(g5669) );
  dffs1 \DFF_281/Q_reg  ( .Q(g700), .CLK(CK), .DIN(g8431) );
  dffs1 \DFF_280/Q_reg  ( .Q(g1663), .CLK(CK), .DIN(g11034) );
  dffs1 \DFF_279/Q_reg  ( .Q(g296), .CLK(CK), .DIN(g7771) );
  dffs1 \DFF_278/Q_reg  ( .QN(n1949), .Q(g1110), .CLK(CK), .DIN(g6817) );
  dffs1 \DFF_277/Q_reg  ( .Q(g1482), .CLK(CK), .DIN(g8443) );
  dffs1 \DFF_276/Q_reg  ( .QN(n2074), .Q(g1690), .CLK(CK), .DIN(g6844) );
  dffs1 \DFF_275/Q_reg  ( .QN(\DFF_275/net562 ), .CLK(CK), .DIN(g4217) );
  dffs1 \DFF_273/Q_reg  ( .Q(g1478), .CLK(CK), .DIN(g8442) );
  dffs1 \DFF_272/Q_reg  ( .Q(g1738), .CLK(CK), .DIN(g5661) );
  dffs1 \DFF_271/Q_reg  ( .QN(n2008), .Q(g1945), .CLK(CK), .DIN(g9356) );
  dffs1 \DFF_270/Q_reg  ( .QN(\DFF_270/net557 ), .Q(g5644), .CLK(CK), .DIN(
        g7751) );
  dffs1 \DFF_269/Q_reg  ( .Q(g865), .CLK(CK), .DIN(g8275) );
  dffs1 \DFF_268/Q_reg  ( .Q(g1771), .CLK(CK), .DIN(g7811) );
  dffs1 \DFF_267/Q_reg  ( .Q(g8), .CLK(CK), .DIN(g2613) );
  dffs1 \DFF_266/Q_reg  ( .Q(g345), .CLK(CK), .DIN(g11642) );
  dffs1 \DFF_265/Q_reg  ( .Q(g305), .CLK(CK), .DIN(g5643) );
  dffs1 \DFF_264/Q_reg  ( .QN(n2073), .Q(g456), .CLK(CK), .DIN(g11466) );
  dffs1 \DFF_263/Q_reg  ( .Q(g336), .CLK(CK), .DIN(g11653) );
  dffs1 \DFF_262/Q_reg  ( .Q(g17), .CLK(CK), .DIN(g4894) );
  dffs1 \DFF_261/Q_reg  ( .QN(n1982), .Q(g617), .CLK(CK), .DIN(g8780) );
  dffs1 \DFF_260/Q_reg  ( .Q(g560), .CLK(CK), .DIN(g11049) );
  dffs1 \DFF_259/Q_reg  ( .Q(g287), .CLK(CK), .DIN(g7768) );
  dffs1 \DFF_258/Q_reg  ( .Q(g1546), .CLK(CK), .DIN(g7345) );
  dffs1 \DFF_256/Q_reg  ( .Q(g1561), .CLK(CK), .DIN(g7350) );
  dffs1 \DFF_255/Q_reg  ( .QN(n1977), .Q(g466), .CLK(CK), .DIN(g11468) );
  dffs1 \DFF_254/Q_reg  ( .Q(g1583), .CLK(CK), .DIN(g7357) );
  dffs1 \DFF_253/Q_reg  ( .Q(g770), .CLK(CK), .DIN(g7288) );
  dffs1 \DFF_252/Q_reg  ( .Q(g1850), .CLK(CK), .DIN(g5671) );
  dffs1 \DFF_251/Q_reg  ( .Q(g290), .CLK(CK), .DIN(g7769) );
  dffs1 \DFF_250/Q_reg  ( .Q(g1292), .CLK(CK), .DIN(g7293) );
  dffs1 \DFF_249/Q_reg  ( .Q(g1627), .CLK(CK), .DIN(g8871) );
  dffs1 \DFF_248/Q_reg  ( .Q(g861), .CLK(CK), .DIN(g4190) );
  dffs1 \DFF_247/Q_reg  ( .Q(g778), .CLK(CK), .DIN(g8076) );
  dffs1 \DFF_246/Q_reg  ( .Q(g5652), .CLK(CK), .DIN(g7759) );
  dffs1 \DFF_245/Q_reg  ( .Q(g516), .CLK(CK), .DIN(g11337) );
  dffs1 \DFF_244/Q_reg  ( .Q(g5650), .CLK(CK), .DIN(g7757) );
  dffs1 \DFF_243/Q_reg  ( .QN(n2047), .Q(g928), .CLK(CK), .DIN(g8569) );
  dffs1 \DFF_242/Q_reg  ( .QN(\DFF_242/net529 ), .CLK(CK), .DIN(g10869) );
  dffs1 \DFF_241/Q_reg  ( .Q(g1357), .CLK(CK), .DIN(g6330) );
  dffs1 \DFF_240/Q_reg  ( .QN(n2005), .CLK(CK), .DIN(g6303) );
  dffs1 \DFF_239/Q_reg  ( .Q(g330), .CLK(CK), .DIN(g5650) );
  dffs1 \DFF_238/Q_reg  ( .Q(g363), .CLK(CK), .DIN(g11511) );
  dffs1 \DFF_237/Q_reg  ( .QN(n2012), .Q(g1453), .CLK(CK), .DIN(g7326) );
  dffs1 \DFF_235/Q_reg  ( .Q(g1432), .CLK(CK), .DIN(g8990) );
  dffs1 \DFF_234/Q_reg  ( .Q(g1032), .CLK(CK), .DIN(g7800) );
  dffs1 \DFF_233/Q_reg  ( .QN(g6919), .CLK(CK), .DIN(g2044) );
  dffs1 \DFF_232/Q_reg  ( .QN(n1942), .CLK(CK), .DIN(g6301) );
  dffs1 \DFF_231/Q_reg  ( .Q(g1250), .CLK(CK), .DIN(g7299) );
  dffs1 \DFF_230/Q_reg  ( .Q(g342), .CLK(CK), .DIN(g11513) );
  dffs1 \DFF_229/Q_reg  ( .Q(g302), .CLK(CK), .DIN(g7773) );
  dffs1 \DFF_228/Q_reg  ( .QN(\DFF_228/net515 ), .CLK(CK), .DIN(g10870) );
  dffs1 \DFF_227/Q_reg  ( .Q(g4182), .CLK(CK), .DIN(g6800) );
  dffs1 \DFF_226/Q_reg  ( .Q(g1356), .CLK(CK), .DIN(g6818) );
  dffs1 \DFF_225/Q_reg  ( .Q(g318), .CLK(CK), .DIN(g5646) );
  dffs1 \DFF_224/Q_reg  ( .QN(n2018), .Q(g8815), .CLK(CK), .DIN(g7783) );
  dffs1 \DFF_223/Q_reg  ( .QN(n1983), .Q(g1840), .CLK(CK), .DIN(g8694) );
  dffs1 \DFF_222/Q_reg  ( .Q(g5651), .CLK(CK), .DIN(g7758) );
  dffs1 \DFF_221/Q_reg  ( .Q(g501), .CLK(CK), .DIN(g11334) );
  dffs1 \DFF_220/Q_reg  ( .Q(g166), .CLK(CK), .DIN(g7747) );
  dffs1 \DFF_218/Q_reg  ( .Q(g1601), .CLK(CK), .DIN(g7363) );
  dffs1 \DFF_217/Q_reg  ( .Q(g386), .CLK(CK), .DIN(g11263) );
  dffs1 \DFF_216/Q_reg  ( .Q(g357), .CLK(CK), .DIN(g11509) );
  dffs1 \DFF_215/Q_reg  ( .Q(g1317), .CLK(CK), .DIN(g1356) );
  dffs1 \DFF_214/Q_reg  ( .QN(n1969), .Q(g1117), .CLK(CK), .DIN(g6299) );
  dffs1 \DFF_213/Q_reg  ( .QN(n2037), .Q(g8810), .CLK(CK), .DIN(g7778) );
  dffs1 \DFF_212/Q_reg  ( .QN(n1993), .Q(g1936), .CLK(CK), .DIN(g9355) );
  dffs1 \DFF_211/Q_reg  ( .Q(g575), .CLK(CK), .DIN(g11052) );
  dffs1 \DFF_210/Q_reg  ( .Q(g530), .CLK(CK), .DIN(g11328) );
  dffs1 \DFF_209/Q_reg  ( .Q(g1914), .CLK(CK), .DIN(g8284) );
  dffs1 \DFF_208/Q_reg  ( .Q(g563), .CLK(CK), .DIN(g11050) );
  dffs1 \DFF_207/Q_reg  ( .Q(g374), .CLK(CK), .DIN(g11440) );
  dffs1 \DFF_206/Q_reg  ( .Q(g1681), .CLK(CK), .DIN(g11040) );
  dffs1 \DFF_205/Q_reg  ( .Q(g542), .CLK(CK), .DIN(g11325) );
  dffs1 \DFF_204/Q_reg  ( .Q(g416), .CLK(CK), .DIN(g11269) );
  dffs1 \DFF_203/Q_reg  ( .Q(g538), .CLK(CK), .DIN(g11326) );
  dffs1 \DFF_202/Q_reg  ( .Q(g1240), .CLK(CK), .DIN(g7297) );
  dffs1 \DFF_201/Q_reg  ( .Q(g1508), .CLK(CK), .DIN(g7329) );
  dffs1 \DFF_200/Q_reg  ( .Q(g1753), .CLK(CK), .DIN(g5666) );
  dffs1 \DFF_199/Q_reg  ( .Q(g1633), .CLK(CK), .DIN(g8873) );
  dffs1 \DFF_198/Q_reg  ( .QN(n2000), .Q(g1346), .CLK(CK), .DIN(g11656) );
  dffs1 \DFF_197/Q_reg  ( .Q(g293), .CLK(CK), .DIN(g7770) );
  dffs1 \DFF_196/Q_reg  ( .Q(g654), .CLK(CK), .DIN(g8067) );
  dffs1 \DFF_195/Q_reg  ( .Q(g1327), .CLK(CK), .DIN(g11633) );
  dffs1 \DFF_194/Q_reg  ( .QN(\DFF_194/net481 ), .CLK(CK), .DIN(g3069) );
  dffs1 \DFF_193/Q_reg  ( .Q(g5648), .CLK(CK), .DIN(g7755) );
  dffs1 \DFF_192/Q_reg  ( .Q(g1023), .CLK(CK), .DIN(g7799) );
  dffs1 \DFF_191/Q_reg  ( .QN(n1997), .CLK(CK), .DIN(g5657) );
  dffs1 \DFF_190/Q_reg  ( .QN(n1992), .Q(g158), .CLK(CK), .DIN(g8425) );
  dffs1 \DFF_189/Q_reg  ( .QN(n1964), .CLK(CK), .DIN(g7316) );
  dffs1 \DFF_188/Q_reg  ( .Q(g869), .CLK(CK), .DIN(g875) );
  dffs1 \DFF_187/Q_reg  ( .Q(g586), .CLK(CK), .DIN(g6294) );
  dffs1 \DFF_186/Q_reg  ( .Q(g557), .CLK(CK), .DIN(g11048) );
  dffs1 \DFF_185/Q_reg  ( .QN(n1947), .Q(g231), .CLK(CK), .DIN(g7319) );
  dffs1 \DFF_184/Q_reg  ( .Q(g4187), .CLK(CK), .DIN(g8077) );
  dffs1 \DFF_183/Q_reg  ( .Q(g309), .CLK(CK), .DIN(g5652) );
  dffs1 \DFF_182/Q_reg  ( .QN(n1973), .CLK(CK), .DIN(g7324) );
  dffs1 \DFF_181/Q_reg  ( .Q(g965), .CLK(CK), .DIN(g11405) );
  dffs1 \DFF_180/Q_reg  ( .Q(g664), .CLK(CK), .DIN(g8782) );
  dffs1 \DFF_179/Q_reg  ( .Q(g9), .CLK(CK), .DIN(g7336) );
  dffs1 \DFF_178/Q_reg  ( .QN(n1989), .Q(g1857), .CLK(CK), .DIN(g11409) );
  dffs1 \DFF_177/Q_reg  ( .Q(g401), .CLK(CK), .DIN(g11266) );
  dffs1 \DFF_176/Q_reg  ( .Q(g269), .CLK(CK), .DIN(g7762) );
  dffs1 \DFF_175/Q_reg  ( .Q(g333), .CLK(CK), .DIN(g5651) );
  dffs1 \DFF_174/Q_reg  ( .QN(n2061), .Q(g5653), .CLK(CK), .DIN(g6336) );
  dffs1 \DFF_173/Q_reg  ( .Q(g1080), .CLK(CK), .DIN(g6806) );
  dffs1 \DFF_172/Q_reg  ( .Q(g1474), .CLK(CK), .DIN(g8441) );
  dffs1 \DFF_171/Q_reg  ( .Q(g444), .CLK(CK), .DIN(g11259) );
  dffs1 \DFF_170/Q_reg  ( .Q(g1074), .CLK(CK), .DIN(g6813) );
  dffs1 \DFF_169/Q_reg  ( .Q(g1411), .CLK(CK), .DIN(g7331) );
  dffs1 \DFF_168/Q_reg  ( .QN(\DFF_168/net455 ), .CLK(CK), .DIN(g10867) );
  dffs1 \DFF_167/Q_reg  ( .Q(g1011), .CLK(CK), .DIN(g7805) );
  dffs1 \DFF_166/Q_reg  ( .Q(g572), .CLK(CK), .DIN(g10877) );
  dffs1 \DFF_165/Q_reg  ( .QN(n1991), .Q(g1458), .CLK(CK), .DIN(g7327) );
  dffs1 \DFF_164/Q_reg  ( .Q(g1531), .CLK(CK), .DIN(g7340) );
  dffs1 \DFF_163/Q_reg  ( .QN(n1940), .CLK(CK), .DIN(g7308) );
  dffs1 \DFF_162/Q_reg  ( .Q(g1669), .CLK(CK), .DIN(g11036) );
  dffs1 \DFF_161/Q_reg  ( .Q(g105), .CLK(CK), .DIN(g11180) );
  dffs1 \DFF_159/Q_reg  ( .Q(g549), .CLK(CK), .DIN(g11044) );
  dffs1 \DFF_158/Q_reg  ( .QN(n1974), .Q(g1101), .CLK(CK), .DIN(g6814) );
  dffs1 \DFF_157/Q_reg  ( .QN(\DFF_157/net444 ), .CLK(CK), .DIN(g5656) );
  dffs1 \DFF_156/Q_reg  ( .Q(g2638), .CLK(CK), .DIN(g755) );
  dffs1 \DFF_155/Q_reg  ( .Q(g1950), .CLK(CK), .DIN(g8288) );
  dffs1 \DFF_154/Q_reg  ( .Q(g580), .CLK(CK), .DIN(g6294) );
  dffs1 \DFF_153/Q_reg  ( .Q(g1397), .CLK(CK), .DIN(g7322) );
  dffs1 \DFF_152/Q_reg  ( .QN(n1950), .Q(g471), .CLK(CK), .DIN(g11469) );
  dffs1 \DFF_151/Q_reg  ( .Q(g486), .CLK(CK), .DIN(g11331) );
  dffs1 \DFF_150/Q_reg  ( .Q(g588), .CLK(CK), .DIN(g6296) );
  dffs1 \DFF_149/Q_reg  ( .QN(n2058), .Q(g766), .CLK(CK), .DIN(g6799) );
  dffs1 \DFF_148/Q_reg  ( .Q(g962), .CLK(CK), .DIN(g11404) );
  dffs1 \DFF_147/Q_reg  ( .QN(n1937), .Q(g153), .CLK(CK), .DIN(g8426) );
  dffs1 \DFF_146/Q_reg  ( .Q(g1333), .CLK(CK), .DIN(g11635) );
  dffs1 \DFF_145/Q_reg  ( .QN(n1971), .Q(g1133), .CLK(CK), .DIN(g6309) );
  dffs1 \DFF_143/Q_reg  ( .Q(g1448), .CLK(CK), .DIN(g11594) );
  dffs1 \DFF_142/Q_reg  ( .Q(g1365), .CLK(CK), .DIN(g7307) );
  dffs1 \DFF_141/Q_reg  ( .Q(g1861), .CLK(CK), .DIN(g7815) );
  dffs1 \DFF_140/Q_reg  ( .Q(g1571), .CLK(CK), .DIN(g7353) );
  dffs1 \DFF_139/Q_reg  ( .Q(g1466), .CLK(CK), .DIN(g8439) );
  dffs1 \DFF_138/Q_reg  ( .Q(g1589), .CLK(CK), .DIN(g7359) );
  dffs1 \DFF_137/Q_reg  ( .Q(g1217), .CLK(CK), .DIN(g9823) );
  dffs1 \DFF_136/Q_reg  ( .QN(\DFF_136/net423 ), .CLK(CK), .DIN(g5654) );
  dffs1 \DFF_135/Q_reg  ( .QN(n1975), .Q(g611), .CLK(CK), .DIN(g9930) );
  dffs1 \DFF_134/Q_reg  ( .Q(g1308), .CLK(CK), .DIN(g11627) );
  dffs1 \DFF_133/Q_reg  ( .Q(g281), .CLK(CK), .DIN(g7766) );
  dffs1 \DFF_132/Q_reg  ( .QN(n2040), .Q(g225), .CLK(CK), .DIN(g7309) );
  dffs1 \DFF_131/Q_reg  ( .Q(g1741), .CLK(CK), .DIN(g5662) );
  dffs1 \DFF_130/Q_reg  ( .Q(g1564), .CLK(CK), .DIN(g7351) );
  dffs1 \DFF_129/Q_reg  ( .Q(g579), .CLK(CK), .DIN(g6293) );
  dffs1 \DFF_128/Q_reg  ( .Q(g1428), .CLK(CK), .DIN(g8992) );
  dffs1 \DFF_127/Q_reg  ( .Q(g4185), .CLK(CK), .DIN(g7289) );
  dffs1 \DFF_126/Q_reg  ( .QN(\DFF_126/net413 ), .CLK(CK), .DIN(g1360) );
  dffs1 \DFF_125/Q_reg  ( .QN(n1972), .Q(g219), .CLK(CK), .DIN(g7310) );
  dffs1 \DFF_124/Q_reg  ( .Q(g426), .CLK(CK), .DIN(g11256) );
  dffs1 \DFF_123/Q_reg  ( .Q(g284), .CLK(CK), .DIN(g7767) );
  dffs1 \DFF_122/Q_reg  ( .Q(g16), .CLK(CK), .DIN(g4906) );
  dffs1 \DFF_121/Q_reg  ( .QN(\DFF_121/net408 ), .CLK(CK), .DIN(g2986) );
  dffs1 \DFF_120/Q_reg  ( .Q(g1721), .CLK(CK), .DIN(g10878) );
  dffs1 \DFF_119/Q_reg  ( .Q(g1227), .CLK(CK), .DIN(g8278) );
  dffs1 \DFF_118/Q_reg  ( .Q(g1415), .CLK(CK), .DIN(g7335) );
  dffs1 \DFF_117/Q_reg  ( .Q(g632), .CLK(CK), .DIN(g5655) );
  dffs1 \DFF_116/Q_reg  ( .Q(g38), .CLK(CK), .DIN(g10872) );
  dffs1 \DFF_115/Q_reg  ( .Q(g1015), .CLK(CK), .DIN(g7808) );
  dffs1 \DFF_114/Q_reg  ( .Q(g396), .CLK(CK), .DIN(g11265) );
  dffs1 \DFF_113/Q_reg  ( .QN(n1979), .Q(g1718), .CLK(CK), .DIN(g6337) );
  dffs1 \DFF_112/Q_reg  ( .Q(g758), .CLK(CK), .DIN(g6797) );
  dffs1 \DFF_111/Q_reg  ( .Q(g1868), .CLK(CK), .DIN(g7817) );
  dffs1 \DFF_109/Q_reg  ( .Q(g1407), .CLK(CK), .DIN(g8993) );
  dffs1 \DFF_108/Q_reg  ( .Q(g1007), .CLK(CK), .DIN(g7806) );
  dffs1 \DFF_106/Q_reg  ( .Q(g959), .CLK(CK), .DIN(g11403) );
  dffs1 \DFF_105/Q_reg  ( .QN(n2041), .Q(g186), .CLK(CK), .DIN(g7317) );
  dffs1 \DFF_104/Q_reg  ( .Q(g1801), .CLK(CK), .DIN(g8450) );
  dffs1 \DFF_103/Q_reg  ( .Q(g1766), .CLK(CK), .DIN(g7810) );
  dffs1 \DFF_102/Q_reg  ( .Q(g174), .CLK(CK), .DIN(g8423) );
  dffs1 \DFF_101/Q_reg  ( .Q(g1678), .CLK(CK), .DIN(g11039) );
  dffs1 \DFF_100/Q_reg  ( .Q(g583), .CLK(CK), .DIN(g6297) );
  dffs1 \DFF_99/Q_reg  ( .QN(n2043), .Q(g4189), .CLK(CK), .DIN(g8437) );
  dffs1 \DFF_98/Q_reg  ( .Q(g1470), .CLK(CK), .DIN(g8440) );
  dffs1 \DFF_97/Q_reg  ( .Q(g1504), .CLK(CK), .DIN(g7328) );
  dffs1 \DFF_96/Q_reg  ( .Q(g1730), .CLK(CK), .DIN(g10881) );
  dffs1 \DFF_95/Q_reg  ( .Q(g1486), .CLK(CK), .DIN(g8444) );
  dffs1 \DFF_94/Q_reg  ( .Q(g1086), .CLK(CK), .DIN(g6808) );
  dffs1 \DFF_93/Q_reg  ( .QN(\DFF_93/net380 ), .CLK(CK), .DIN(g3007) );
  dffs1 \DFF_92/Q_reg  ( .QN(n2030), .CLK(CK), .DIN(g11397) );
  dffs1 \DFF_91/Q_reg  ( .QN(n2020), .Q(g8811), .CLK(CK), .DIN(g7779) );
  dffs1 \DFF_90/Q_reg  ( .Q(g1419), .CLK(CK), .DIN(g7332) );
  dffs1 \DFF_89/Q_reg  ( .Q(g745), .CLK(CK), .DIN(g2639) );
  dffs1 \DFF_88/Q_reg  ( .Q(g1362), .CLK(CK), .DIN(g7305) );
  dffs1 \DFF_87/Q_reg  ( .Q(g1019), .CLK(CK), .DIN(g7807) );
  dffs1 \DFF_86/Q_reg  ( .Q(g736), .CLK(CK), .DIN(g8435) );
  dffs1 \DFF_85/Q_reg  ( .Q(g1896), .CLK(CK), .DIN(g8282) );
  dffs1 \DFF_83/Q_reg  ( .QN(n2007), .Q(g932), .CLK(CK), .DIN(g8570) );
  dffs1 \DFF_82/Q_reg  ( .Q(g1098), .CLK(CK), .DIN(g6812) );
  dffs1 \DFF_81/Q_reg  ( .Q(g1604), .CLK(CK), .DIN(g7364) );
  dffs1 \DFF_80/Q_reg  ( .Q(g1957), .CLK(CK), .DIN(g1956) );
  dffs1 \DFF_79/Q_reg  ( .Q(g351), .CLK(CK), .DIN(g11507) );
  dffs1 \DFF_78/Q_reg  ( .Q(g1759), .CLK(CK), .DIN(g5668) );
  dffs1 \DFF_77/Q_reg  ( .Q(g1707), .CLK(CK), .DIN(g4907) );
  dffs1 \DFF_76/Q_reg  ( .QN(n1963), .Q(g248), .CLK(CK), .DIN(g7323) );
  dffs1 \DFF_75/Q_reg  ( .QN(n2025), .Q(g1791), .CLK(CK), .DIN(g8080) );
  dffs1 \DFF_74/Q_reg  ( .Q(g1639), .CLK(CK), .DIN(g8448) );
  dffs1 \DFF_73/Q_reg  ( .Q(g1684), .CLK(CK), .DIN(g11041) );
  dffs1 \DFF_72/Q_reg  ( .QN(n1981), .Q(g639), .CLK(CK), .DIN(g8063) );
  dffs1 \DFF_71/Q_reg  ( .Q(g113), .CLK(CK), .DIN(g7285) );
  dffs1 \DFF_70/Q_reg  ( .Q(g354), .CLK(CK), .DIN(g11508) );
  dffs1 \DFF_69/Q_reg  ( .Q(g1675), .CLK(CK), .DIN(g11038) );
  dffs1 \DFF_68/Q_reg  ( .Q(g1956), .CLK(CK), .DIN(g1955) );
  dffs1 \DFF_67/Q_reg  ( .QN(n2003), .CLK(CK), .DIN(g7311) );
  dffs1 \DFF_66/Q_reg  ( .Q(g1389), .CLK(CK), .DIN(g6836) );
  dffs1 \DFF_65/Q_reg  ( .Q(g327), .CLK(CK), .DIN(g5649) );
  dffs1 \DFF_64/Q_reg  ( .Q(g646), .CLK(CK), .DIN(g8065) );
  dffs1 \DFF_63/Q_reg  ( .QN(n2021), .Q(g8806), .CLK(CK), .DIN(g7777) );
  dffs1 \DFF_62/Q_reg  ( .Q(g587), .CLK(CK), .DIN(g6295) );
  dffs1 \DFF_61/Q_reg  ( .Q(g1296), .CLK(CK), .DIN(g7292) );
  dffs1 \DFF_60/Q_reg  ( .Q(g682), .CLK(CK), .DIN(g8429) );
  dffs1 \DFF_59/Q_reg  ( .Q(g1786), .CLK(CK), .DIN(g7814) );
  dffs1 \DFF_58/Q_reg  ( .Q(g1265), .CLK(CK), .DIN(g7302) );
  dffs1 \DFF_57/Q_reg  ( .QN(n2029), .Q(g704), .CLK(CK), .DIN(g9344) );
  dffs1 \DFF_56/Q_reg  ( .Q(g1095), .CLK(CK), .DIN(g6811) );
  dffs1 \DFF_55/Q_reg  ( .Q(g829), .CLK(CK), .DIN(g4182) );
  dffs1 \DFF_54/Q_reg  ( .Q(g590), .CLK(CK), .DIN(n2062) );
  dffs1 \DFF_53/Q_reg  ( .Q(g3007), .CLK(CK), .DIN(g4896) );
  dffs1 \DFF_52/Q_reg  ( .Q(g981), .CLK(CK), .DIN(g11472) );
  dffs1 \DFF_51/Q_reg  ( .Q(g496), .CLK(CK), .DIN(g11333) );
  dffs1 \DFF_50/Q_reg  ( .Q(g554), .CLK(CK), .DIN(g11047) );
  dffs1 \DFF_49/Q_reg  ( .QN(n2023), .Q(g8818), .CLK(CK), .DIN(g7775) );
  dffs1 \DFF_48/Q_reg  ( .Q(g718), .CLK(CK), .DIN(g8433) );
  dffs1 \DFF_47/Q_reg  ( .Q(g1436), .CLK(CK), .DIN(g8989) );
  dffs1 \DFF_46/Q_reg  ( .Q(g278), .CLK(CK), .DIN(g7765) );
  dffs1 \DFF_45/Q_reg  ( .Q(g1660), .CLK(CK), .DIN(g11033) );
  dffs1 \DFF_44/Q_reg  ( .QN(n1954), .Q(g1927), .CLK(CK), .DIN(g9354) );
  dffs1 \DFF_43/Q_reg  ( .QN(n1987), .Q(g622), .CLK(CK), .DIN(g9338) );
  dffs1 \DFF_42/Q_reg  ( .Q(g1534), .CLK(CK), .DIN(g7341) );
  dffs1 \DFF_41/Q_reg  ( .Q(g315), .CLK(CK), .DIN(g5645) );
  dffs1 \DFF_39/Q_reg  ( .Q(g1543), .CLK(CK), .DIN(g7344) );
  dffs1 \DFF_38/Q_reg  ( .Q(g786), .CLK(CK), .DIN(g8436) );
  dffs1 \DFF_37/Q_reg  ( .Q(g757), .CLK(CK), .DIN(g11179) );
  dffs1 \DFF_36/Q_reg  ( .Q(g1444), .CLK(CK), .DIN(g8987) );
  dffs1 \DFF_34/Q_reg  ( .Q(g1499), .CLK(CK), .DIN(g8447) );
  dffs1 \DFF_33/Q_reg  ( .QN(n2002), .Q(g243), .CLK(CK), .DIN(g7325) );
  dffs1 \DFF_32/Q_reg  ( .Q(g1304), .CLK(CK), .DIN(g7290) );
  dffs1 \DFF_31/Q_reg  ( .QN(n1976), .Q(g1104), .CLK(CK), .DIN(g6815) );
  dffs1 \DFF_30/Q_reg  ( .QN(n2057), .Q(g774), .CLK(CK), .DIN(g7785) );
  dffs1 \DFF_29/Q_reg  ( .Q(g4), .CLK(CK), .DIN(g8079) );
  dffs1 \DFF_28/Q_reg  ( .QN(n2048), .Q(g1231), .CLK(CK), .DIN(g8279) );
  dffs1 \DFF_27/Q_reg  ( .Q(g1077), .CLK(CK), .DIN(g6805) );
  dffs1 \DFF_26/Q_reg  ( .Q(g1672), .CLK(CK), .DIN(g11037) );
  dffs1 \DFF_25/Q_reg  ( .Q(g1737), .CLK(CK), .DIN(g1736) );
  dffs1 \DFF_24/Q_reg  ( .Q(g1424), .CLK(CK), .DIN(g7330) );
  dffs1 \DFF_23/Q_reg  ( .QN(n1928), .CLK(CK), .DIN(g11182) );
  dffs1 \DFF_22/Q_reg  ( .Q(g39), .CLK(CK), .DIN(g10774) );
  dffs1 \DFF_21/Q_reg  ( .Q(g1736), .CLK(CK), .DIN(g6846) );
  dffs1 \DFF_20/Q_reg  ( .Q(g1580), .CLK(CK), .DIN(g7356) );
  dffs1 \DFF_19/Q_reg  ( .Q(g369), .CLK(CK), .DIN(g11439) );
  dffs1 \DFF_18/Q_reg  ( .QN(n2027), .CLK(CK), .DIN(g7816) );
  dffs1 \DFF_17/Q_reg  ( .Q(g1574), .CLK(CK), .DIN(g7354) );
  dffs1 \DFF_16/Q_reg  ( .Q(g1092), .CLK(CK), .DIN(g6810) );
  dffs1 \DFF_15/Q_reg  ( .Q(g709), .CLK(CK), .DIN(g8432) );
  dffs1 \DFF_14/Q_reg  ( .QN(n2044), .Q(g976), .CLK(CK), .DIN(g11471) );
  dffs1 \DFF_13/Q_reg  ( .QN(n2045), .Q(g940), .CLK(CK), .DIN(g8572) );
  dffs1 \DFF_12/Q_reg  ( .QN(n1930), .Q(g461), .CLK(CK), .DIN(g11467) );
  dffs1 \DFF_11/Q_reg  ( .QN(n1958), .Q(g695), .CLK(CK), .DIN(g9343) );
  dffs1 \DFF_10/Q_reg  ( .Q(g1558), .CLK(CK), .DIN(g7349) );
  dffs1 \DFF_9/Q_reg  ( .Q(g1744), .CLK(CK), .DIN(g5663) );
  dffs1 \DFF_7/Q_reg  ( .QN(n1988), .Q(g1153), .CLK(CK), .DIN(g6304) );
  dffs1 \DFF_6/Q_reg  ( .QN(n1955), .Q(g713), .CLK(CK), .DIN(g9345) );
  dffs1 \DFF_5/Q_reg  ( .QN(n2001), .Q(g207), .CLK(CK), .DIN(g7315) );
  dffs1 \DFF_4/Q_reg  ( .Q(g123), .CLK(CK), .DIN(g8272) );
  dffs1 \DFF_3/Q_reg  ( .Q(g452), .CLK(CK), .DIN(g11257) );
  dffs1 \DFF_2/Q_reg  ( .Q(g312), .CLK(CK), .DIN(g5644) );
  dffs1 \DFF_1/Q_reg  ( .QN(n1935), .Q(g1882), .CLK(CK), .DIN(g9349) );
  dffs1 \DFF_0/Q_reg  ( .Q(g1289), .CLK(CK), .DIN(g5660) );
endmodule

