module c880 (N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880);

input N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268;

output N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880;

wire N269, N270, N273, N276, N279, N280, N284, N285, N286, N287, N290, N291, N292, N293, N294, N295, N296, N297, N298, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N316, N317, N318, N319, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N360, N363, N366, N369, N375, N376, N379, N382, N385, N392, N393, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N424, N425, N426, N427, N432, N437, N442, N443, N444, N445, N451, N460, N463, N466, N475, N476, N477, N478, N479, N480, N481, N482, N483, N488, N489, N490, N491, N492, N495, N498, N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N533, N536, N537, N538, N539, N540, N541, N542, N543, N544, N547, N550, N551, N552, N553, N557, N561, N565, N569, N573, N577, N581, N585, N586, N587, N588, N589, N590, N593, N596, N597, N600, N605, N606, N609, N615, N616, N619, N624, N625, N628, N631, N632, N635, N640, N641, N644, N650, N651, N654, N659, N660, N661, N662, N665, N669, N670, N673, N677, N678, N682, N686, N687, N692, N696, N697, N700, N704, N705, N708, N712, N713, N717, N721, N722, N727, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763, N764, N765, N766, N769, N770, N771, N772, N773, N777, N778, N781, N782, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796, N802, N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N819, N822, N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862, N867, N868, N869, N870, N871, N872, N873, N875, N876, N877;

nnd4s1 U1 (.Q(N269), .DIN1(N1), .DIN2(N8), .DIN3(N13), .DIN4(N17));
nnd4s1 U2 (.Q(N270), .DIN1(N1), .DIN2(N26), .DIN3(N13), .DIN4(N17));
and3s1 U3 (.Q(N273), .DIN1(N29), .DIN2(N36), .DIN3(N42));
and3s1 U4 (.Q(N276), .DIN1(N1), .DIN2(N26), .DIN3(N51));
nnd4s1 U5 (.Q(N279), .DIN1(N1), .DIN2(N8), .DIN3(N51), .DIN4(N17));
nnd4s1 U6 (.Q(N280), .DIN1(N1), .DIN2(N8), .DIN3(N13), .DIN4(N55));
nnd4s1 U7 (.Q(N284), .DIN1(N59), .DIN2(N42), .DIN3(N68), .DIN4(N72));
nnd2s1 U8 (.Q(N285), .DIN1(N29), .DIN2(N68));
nnd3s1 U9 (.Q(N286), .DIN1(N59), .DIN2(N68), .DIN3(N74));
and3s1 U10 (.Q(N287), .DIN1(N29), .DIN2(N75), .DIN3(N80));
and3s1 U11 (.Q(N290), .DIN1(N29), .DIN2(N75), .DIN3(N42));
and3s1 U12 (.Q(N291), .DIN1(N29), .DIN2(N36), .DIN3(N80));
and3s1 U13 (.Q(N292), .DIN1(N29), .DIN2(N36), .DIN3(N42));
and3s1 U14 (.Q(N293), .DIN1(N59), .DIN2(N75), .DIN3(N80));
and3s1 U15 (.Q(N294), .DIN1(N59), .DIN2(N75), .DIN3(N42));
and3s1 U16 (.Q(N295), .DIN1(N59), .DIN2(N36), .DIN3(N80));
and3s1 U17 (.Q(N296), .DIN1(N59), .DIN2(N36), .DIN3(N42));
and2s1 U18 (.Q(N297), .DIN1(N85), .DIN2(N86));
or2s1 U19 (.Q(N298), .DIN1(N87), .DIN2(N88));
nnd2s1 U20 (.Q(N301), .DIN1(N91), .DIN2(N96));
or2s1 U21 (.Q(N302), .DIN1(N91), .DIN2(N96));
nnd2s1 U22 (.Q(N303), .DIN1(N101), .DIN2(N106));
or2s1 U23 (.Q(N304), .DIN1(N101), .DIN2(N106));
nnd2s1 U24 (.Q(N305), .DIN1(N111), .DIN2(N116));
or2s1 U25 (.Q(N306), .DIN1(N111), .DIN2(N116));
nnd2s1 U26 (.Q(N307), .DIN1(N121), .DIN2(N126));
or2s1 U27 (.Q(N308), .DIN1(N121), .DIN2(N126));
and2s1 U28 (.Q(N309), .DIN1(N8), .DIN2(N138));
hi1s1 U29 (.Q(N310), .DIN(N268));
and2s1 U30 (.Q(N316), .DIN1(N51), .DIN2(N138));
and2s1 U31 (.Q(N317), .DIN1(N17), .DIN2(N138));
and2s1 U32 (.Q(N318), .DIN1(N152), .DIN2(N138));
nnd2s1 U33 (.Q(N319), .DIN1(N59), .DIN2(N156));
nor2s1 U34 (.Q(N322), .DIN1(N17), .DIN2(N42));
and2s1 U35 (.Q(N323), .DIN1(N17), .DIN2(N42));
nnd2s1 U36 (.Q(N324), .DIN1(N159), .DIN2(N165));
or2s1 U37 (.Q(N325), .DIN1(N159), .DIN2(N165));
nnd2s1 U38 (.Q(N326), .DIN1(N171), .DIN2(N177));
or2s1 U39 (.Q(N327), .DIN1(N171), .DIN2(N177));
nnd2s1 U40 (.Q(N328), .DIN1(N183), .DIN2(N189));
or2s1 U41 (.Q(N329), .DIN1(N183), .DIN2(N189));
nnd2s1 U42 (.Q(N330), .DIN1(N195), .DIN2(N201));
or2s1 U43 (.Q(N331), .DIN1(N195), .DIN2(N201));
and2s1 U44 (.Q(N332), .DIN1(N210), .DIN2(N91));
and2s1 U45 (.Q(N333), .DIN1(N210), .DIN2(N96));
and2s1 U46 (.Q(N334), .DIN1(N210), .DIN2(N101));
and2s1 U47 (.Q(N335), .DIN1(N210), .DIN2(N106));
and2s1 U48 (.Q(N336), .DIN1(N210), .DIN2(N111));
and2s1 U49 (.Q(N337), .DIN1(N255), .DIN2(N259));
and2s1 U50 (.Q(N338), .DIN1(N210), .DIN2(N116));
and2s1 U51 (.Q(N339), .DIN1(N255), .DIN2(N260));
and2s1 U52 (.Q(N340), .DIN1(N210), .DIN2(N121));
and2s1 U53 (.Q(N341), .DIN1(N255), .DIN2(N267));
hi1s1 U54 (.Q(N342), .DIN(N269));
hi1s1 U55 (.Q(N343), .DIN(N273));
or2s1 U56 (.Q(N344), .DIN1(N270), .DIN2(N273));
hi1s1 U57 (.Q(N345), .DIN(N276));
hi1s1 U58 (.Q(N346), .DIN(N276));
hi1s1 U59 (.Q(N347), .DIN(N279));
nor2s1 U60 (.Q(N348), .DIN1(N280), .DIN2(N284));
or2s1 U61 (.Q(N349), .DIN1(N280), .DIN2(N285));
or2s1 U62 (.Q(N350), .DIN1(N280), .DIN2(N286));
hi1s1 U63 (.Q(N351), .DIN(N293));
hi1s1 U64 (.Q(N352), .DIN(N294));
hi1s1 U65 (.Q(N353), .DIN(N295));
hi1s1 U66 (.Q(N354), .DIN(N296));
nnd2s1 U67 (.Q(N355), .DIN1(N89), .DIN2(N298));
and2s1 U68 (.Q(N356), .DIN1(N90), .DIN2(N298));
nnd2s1 U69 (.Q(N357), .DIN1(N301), .DIN2(N302));
nnd2s1 U70 (.Q(N360), .DIN1(N303), .DIN2(N304));
nnd2s1 U71 (.Q(N363), .DIN1(N305), .DIN2(N306));
nnd2s1 U72 (.Q(N366), .DIN1(N307), .DIN2(N308));
hi1s1 U73 (.Q(N369), .DIN(N310));
nor2s1 U74 (.Q(N375), .DIN1(N322), .DIN2(N323));
nnd2s1 U75 (.Q(N376), .DIN1(N324), .DIN2(N325));
nnd2s1 U76 (.Q(N379), .DIN1(N326), .DIN2(N327));
nnd2s1 U77 (.Q(N382), .DIN1(N328), .DIN2(N329));
nnd2s1 U78 (.Q(N385), .DIN1(N330), .DIN2(N331));
nb1s1 U79 (.Q(N388), .DIN(N290));
nb1s1 U80 (.Q(N389), .DIN(N291));
nb1s1 U81 (.Q(N390), .DIN(N292));
nb1s1 U82 (.Q(N391), .DIN(N297));
or2s1 U83 (.Q(N392), .DIN1(N270), .DIN2(N343));
hi1s1 U84 (.Q(N393), .DIN(N345));
hi1s1 U85 (.Q(N399), .DIN(N346));
and2s1 U86 (.Q(N400), .DIN1(N348), .DIN2(N73));
hi1s1 U87 (.Q(N401), .DIN(N349));
hi1s1 U88 (.Q(N402), .DIN(N350));
hi1s1 U89 (.Q(N403), .DIN(N355));
hi1s1 U90 (.Q(N404), .DIN(N357));
hi1s1 U91 (.Q(N405), .DIN(N360));
and2s1 U92 (.Q(N406), .DIN1(N357), .DIN2(N360));
hi1s1 U93 (.Q(N407), .DIN(N363));
hi1s1 U94 (.Q(N408), .DIN(N366));
and2s1 U95 (.Q(N409), .DIN1(N363), .DIN2(N366));
nnd2s1 U96 (.Q(N410), .DIN1(N347), .DIN2(N352));
hi1s1 U97 (.Q(N411), .DIN(N376));
hi1s1 U98 (.Q(N412), .DIN(N379));
and2s1 U99 (.Q(N413), .DIN1(N376), .DIN2(N379));
hi1s1 U100 (.Q(N414), .DIN(N382));
hi1s1 U101 (.Q(N415), .DIN(N385));
and2s1 U102 (.Q(N416), .DIN1(N382), .DIN2(N385));
and2s1 U103 (.Q(N417), .DIN1(N210), .DIN2(N369));
nb1s1 U104 (.Q(N418), .DIN(N342));
nb1s1 U105 (.Q(N419), .DIN(N344));
nb1s1 U106 (.Q(N420), .DIN(N351));
nb1s1 U107 (.Q(N421), .DIN(N353));
nb1s1 U108 (.Q(N422), .DIN(N354));
nb1s1 U109 (.Q(N423), .DIN(N356));
hi1s1 U110 (.Q(N424), .DIN(N400));
and2s1 U111 (.Q(N425), .DIN1(N404), .DIN2(N405));
and2s1 U112 (.Q(N426), .DIN1(N407), .DIN2(N408));
and3s1 U113 (.Q(N427), .DIN1(N319), .DIN2(N393), .DIN3(N55));
and3s1 U114 (.Q(N432), .DIN1(N393), .DIN2(N17), .DIN3(N287));
nnd3s1 U115 (.Q(N437), .DIN1(N393), .DIN2(N287), .DIN3(N55));
nnd4s1 U116 (.Q(N442), .DIN1(N375), .DIN2(N59), .DIN3(N156), .DIN4(N393));
nnd3s1 U117 (.Q(N443), .DIN1(N393), .DIN2(N319), .DIN3(N17));
and2s1 U118 (.Q(N444), .DIN1(N411), .DIN2(N412));
and2s1 U119 (.Q(N445), .DIN1(N414), .DIN2(N415));
nb1s1 U120 (.Q(N446), .DIN(N392));
nb1s1 U121 (.Q(N447), .DIN(N399));
nb1s1 U122 (.Q(N448), .DIN(N401));
nb1s1 U123 (.Q(N449), .DIN(N402));
nb1s1 U124 (.Q(N450), .DIN(N403));
hi1s1 U125 (.Q(N451), .DIN(N424));
nor2s1 U126 (.Q(N460), .DIN1(N406), .DIN2(N425));
nor2s1 U127 (.Q(N463), .DIN1(N409), .DIN2(N426));
nnd2s1 U128 (.Q(N466), .DIN1(N442), .DIN2(N410));
and2s1 U129 (.Q(N475), .DIN1(N143), .DIN2(N427));
and2s1 U130 (.Q(N476), .DIN1(N310), .DIN2(N432));
and2s1 U131 (.Q(N477), .DIN1(N146), .DIN2(N427));
and2s1 U132 (.Q(N478), .DIN1(N310), .DIN2(N432));
and2s1 U133 (.Q(N479), .DIN1(N149), .DIN2(N427));
and2s1 U134 (.Q(N480), .DIN1(N310), .DIN2(N432));
and2s1 U135 (.Q(N481), .DIN1(N153), .DIN2(N427));
and2s1 U136 (.Q(N482), .DIN1(N310), .DIN2(N432));
nnd2s1 U137 (.Q(N483), .DIN1(N443), .DIN2(N1));
or2s1 U138 (.Q(N488), .DIN1(N369), .DIN2(N437));
or2s1 U139 (.Q(N489), .DIN1(N369), .DIN2(N437));
or2s1 U140 (.Q(N490), .DIN1(N369), .DIN2(N437));
or2s1 U141 (.Q(N491), .DIN1(N369), .DIN2(N437));
nor2s1 U142 (.Q(N492), .DIN1(N413), .DIN2(N444));
nor2s1 U143 (.Q(N495), .DIN1(N416), .DIN2(N445));
nnd2s1 U144 (.Q(N498), .DIN1(N130), .DIN2(N460));
or2s1 U145 (.Q(N499), .DIN1(N130), .DIN2(N460));
nnd2s1 U146 (.Q(N500), .DIN1(N463), .DIN2(N135));
or2s1 U147 (.Q(N501), .DIN1(N463), .DIN2(N135));
and2s1 U148 (.Q(N502), .DIN1(N91), .DIN2(N466));
nor2s1 U149 (.Q(N503), .DIN1(N475), .DIN2(N476));
and2s1 U150 (.Q(N504), .DIN1(N96), .DIN2(N466));
nor2s1 U151 (.Q(N505), .DIN1(N477), .DIN2(N478));
and2s1 U152 (.Q(N506), .DIN1(N101), .DIN2(N466));
nor2s1 U153 (.Q(N507), .DIN1(N479), .DIN2(N480));
and2s1 U154 (.Q(N508), .DIN1(N106), .DIN2(N466));
nor2s1 U155 (.Q(N509), .DIN1(N481), .DIN2(N482));
and2s1 U156 (.Q(N510), .DIN1(N143), .DIN2(N483));
and2s1 U157 (.Q(N511), .DIN1(N111), .DIN2(N466));
and2s1 U158 (.Q(N512), .DIN1(N146), .DIN2(N483));
and2s1 U159 (.Q(N513), .DIN1(N116), .DIN2(N466));
and2s1 U160 (.Q(N514), .DIN1(N149), .DIN2(N483));
and2s1 U161 (.Q(N515), .DIN1(N121), .DIN2(N466));
and2s1 U162 (.Q(N516), .DIN1(N153), .DIN2(N483));
and2s1 U163 (.Q(N517), .DIN1(N126), .DIN2(N466));
nnd2s1 U164 (.Q(N518), .DIN1(N130), .DIN2(N492));
or2s1 U165 (.Q(N519), .DIN1(N130), .DIN2(N492));
nnd2s1 U166 (.Q(N520), .DIN1(N495), .DIN2(N207));
or2s1 U167 (.Q(N521), .DIN1(N495), .DIN2(N207));
and2s1 U168 (.Q(N522), .DIN1(N451), .DIN2(N159));
and2s1 U169 (.Q(N523), .DIN1(N451), .DIN2(N165));
and2s1 U170 (.Q(N524), .DIN1(N451), .DIN2(N171));
and2s1 U171 (.Q(N525), .DIN1(N451), .DIN2(N177));
and2s1 U172 (.Q(N526), .DIN1(N451), .DIN2(N183));
nnd2s1 U173 (.Q(N527), .DIN1(N451), .DIN2(N189));
nnd2s1 U174 (.Q(N528), .DIN1(N451), .DIN2(N195));
nnd2s1 U175 (.Q(N529), .DIN1(N451), .DIN2(N201));
nnd2s1 U176 (.Q(N530), .DIN1(N498), .DIN2(N499));
nnd2s1 U177 (.Q(N533), .DIN1(N500), .DIN2(N501));
nor2s1 U178 (.Q(N536), .DIN1(N309), .DIN2(N502));
nor2s1 U179 (.Q(N537), .DIN1(N316), .DIN2(N504));
nor2s1 U180 (.Q(N538), .DIN1(N317), .DIN2(N506));
nor2s1 U181 (.Q(N539), .DIN1(N318), .DIN2(N508));
nor2s1 U182 (.Q(N540), .DIN1(N510), .DIN2(N511));
nor2s1 U183 (.Q(N541), .DIN1(N512), .DIN2(N513));
nor2s1 U184 (.Q(N542), .DIN1(N514), .DIN2(N515));
nor2s1 U185 (.Q(N543), .DIN1(N516), .DIN2(N517));
nnd2s1 U186 (.Q(N544), .DIN1(N518), .DIN2(N519));
nnd2s1 U187 (.Q(N547), .DIN1(N520), .DIN2(N521));
hi1s1 U188 (.Q(N550), .DIN(N530));
hi1s1 U189 (.Q(N551), .DIN(N533));
and2s1 U190 (.Q(N552), .DIN1(N530), .DIN2(N533));
nnd2s1 U191 (.Q(N553), .DIN1(N536), .DIN2(N503));
nnd2s1 U192 (.Q(N557), .DIN1(N537), .DIN2(N505));
nnd2s1 U193 (.Q(N561), .DIN1(N538), .DIN2(N507));
nnd2s1 U194 (.Q(N565), .DIN1(N539), .DIN2(N509));
nnd2s1 U195 (.Q(N569), .DIN1(N488), .DIN2(N540));
nnd2s1 U196 (.Q(N573), .DIN1(N489), .DIN2(N541));
nnd2s1 U197 (.Q(N577), .DIN1(N490), .DIN2(N542));
nnd2s1 U198 (.Q(N581), .DIN1(N491), .DIN2(N543));
hi1s1 U199 (.Q(N585), .DIN(N544));
hi1s1 U200 (.Q(N586), .DIN(N547));
and2s1 U201 (.Q(N587), .DIN1(N544), .DIN2(N547));
and2s1 U202 (.Q(N588), .DIN1(N550), .DIN2(N551));
and2s1 U203 (.Q(N589), .DIN1(N585), .DIN2(N586));
nnd2s1 U204 (.Q(N590), .DIN1(N553), .DIN2(N159));
or2s1 U205 (.Q(N593), .DIN1(N553), .DIN2(N159));
and2s1 U206 (.Q(N596), .DIN1(N246), .DIN2(N553));
nnd2s1 U207 (.Q(N597), .DIN1(N557), .DIN2(N165));
or2s1 U208 (.Q(N600), .DIN1(N557), .DIN2(N165));
and2s1 U209 (.Q(N605), .DIN1(N246), .DIN2(N557));
nnd2s1 U210 (.Q(N606), .DIN1(N561), .DIN2(N171));
or2s1 U211 (.Q(N609), .DIN1(N561), .DIN2(N171));
and2s1 U212 (.Q(N615), .DIN1(N246), .DIN2(N561));
nnd2s1 U213 (.Q(N616), .DIN1(N565), .DIN2(N177));
or2s1 U214 (.Q(N619), .DIN1(N565), .DIN2(N177));
and2s1 U215 (.Q(N624), .DIN1(N246), .DIN2(N565));
nnd2s1 U216 (.Q(N625), .DIN1(N569), .DIN2(N183));
or2s1 U217 (.Q(N628), .DIN1(N569), .DIN2(N183));
and2s1 U218 (.Q(N631), .DIN1(N246), .DIN2(N569));
nnd2s1 U219 (.Q(N632), .DIN1(N573), .DIN2(N189));
or2s1 U220 (.Q(N635), .DIN1(N573), .DIN2(N189));
and2s1 U221 (.Q(N640), .DIN1(N246), .DIN2(N573));
nnd2s1 U222 (.Q(N641), .DIN1(N577), .DIN2(N195));
or2s1 U223 (.Q(N644), .DIN1(N577), .DIN2(N195));
and2s1 U224 (.Q(N650), .DIN1(N246), .DIN2(N577));
nnd2s1 U225 (.Q(N651), .DIN1(N581), .DIN2(N201));
or2s1 U226 (.Q(N654), .DIN1(N581), .DIN2(N201));
and2s1 U227 (.Q(N659), .DIN1(N246), .DIN2(N581));
nor2s1 U228 (.Q(N660), .DIN1(N552), .DIN2(N588));
nor2s1 U229 (.Q(N661), .DIN1(N587), .DIN2(N589));
hi1s1 U230 (.Q(N662), .DIN(N590));
and2s1 U231 (.Q(N665), .DIN1(N593), .DIN2(N590));
nor2s1 U232 (.Q(N669), .DIN1(N596), .DIN2(N522));
hi1s1 U233 (.Q(N670), .DIN(N597));
and2s1 U234 (.Q(N673), .DIN1(N600), .DIN2(N597));
nor2s1 U235 (.Q(N677), .DIN1(N605), .DIN2(N523));
hi1s1 U236 (.Q(N678), .DIN(N606));
and2s1 U237 (.Q(N682), .DIN1(N609), .DIN2(N606));
nor2s1 U238 (.Q(N686), .DIN1(N615), .DIN2(N524));
hi1s1 U239 (.Q(N687), .DIN(N616));
and2s1 U240 (.Q(N692), .DIN1(N619), .DIN2(N616));
nor2s1 U241 (.Q(N696), .DIN1(N624), .DIN2(N525));
hi1s1 U242 (.Q(N697), .DIN(N625));
and2s1 U243 (.Q(N700), .DIN1(N628), .DIN2(N625));
nor2s1 U244 (.Q(N704), .DIN1(N631), .DIN2(N526));
hi1s1 U245 (.Q(N705), .DIN(N632));
and2s1 U246 (.Q(N708), .DIN1(N635), .DIN2(N632));
nor2s1 U247 (.Q(N712), .DIN1(N337), .DIN2(N640));
hi1s1 U248 (.Q(N713), .DIN(N641));
and2s1 U249 (.Q(N717), .DIN1(N644), .DIN2(N641));
nor2s1 U250 (.Q(N721), .DIN1(N339), .DIN2(N650));
hi1s1 U251 (.Q(N722), .DIN(N651));
and2s1 U252 (.Q(N727), .DIN1(N654), .DIN2(N651));
nor2s1 U253 (.Q(N731), .DIN1(N341), .DIN2(N659));
nnd2s1 U254 (.Q(N732), .DIN1(N654), .DIN2(N261));
nnd3s1 U255 (.Q(N733), .DIN1(N644), .DIN2(N654), .DIN3(N261));
nnd4s1 U256 (.Q(N734), .DIN1(N635), .DIN2(N644), .DIN3(N654), .DIN4(N261));
hi1s1 U257 (.Q(N735), .DIN(N662));
and2s1 U258 (.Q(N736), .DIN1(N228), .DIN2(N665));
and2s1 U259 (.Q(N737), .DIN1(N237), .DIN2(N662));
hi1s1 U260 (.Q(N738), .DIN(N670));
and2s1 U261 (.Q(N739), .DIN1(N228), .DIN2(N673));
and2s1 U262 (.Q(N740), .DIN1(N237), .DIN2(N670));
hi1s1 U263 (.Q(N741), .DIN(N678));
and2s1 U264 (.Q(N742), .DIN1(N228), .DIN2(N682));
and2s1 U265 (.Q(N743), .DIN1(N237), .DIN2(N678));
hi1s1 U266 (.Q(N744), .DIN(N687));
and2s1 U267 (.Q(N745), .DIN1(N228), .DIN2(N692));
and2s1 U268 (.Q(N746), .DIN1(N237), .DIN2(N687));
hi1s1 U269 (.Q(N747), .DIN(N697));
and2s1 U270 (.Q(N748), .DIN1(N228), .DIN2(N700));
and2s1 U271 (.Q(N749), .DIN1(N237), .DIN2(N697));
hi1s1 U272 (.Q(N750), .DIN(N705));
and2s1 U273 (.Q(N751), .DIN1(N228), .DIN2(N708));
and2s1 U274 (.Q(N752), .DIN1(N237), .DIN2(N705));
hi1s1 U275 (.Q(N753), .DIN(N713));
and2s1 U276 (.Q(N754), .DIN1(N228), .DIN2(N717));
and2s1 U277 (.Q(N755), .DIN1(N237), .DIN2(N713));
hi1s1 U278 (.Q(N756), .DIN(N722));
nor2s1 U279 (.Q(N757), .DIN1(N727), .DIN2(N261));
and2s1 U280 (.Q(N758), .DIN1(N727), .DIN2(N261));
and2s1 U281 (.Q(N759), .DIN1(N228), .DIN2(N727));
and2s1 U282 (.Q(N760), .DIN1(N237), .DIN2(N722));
nnd2s1 U283 (.Q(N761), .DIN1(N644), .DIN2(N722));
nnd2s1 U284 (.Q(N762), .DIN1(N635), .DIN2(N713));
nnd3s1 U285 (.Q(N763), .DIN1(N635), .DIN2(N644), .DIN3(N722));
nnd2s1 U286 (.Q(N764), .DIN1(N609), .DIN2(N687));
nnd2s1 U287 (.Q(N765), .DIN1(N600), .DIN2(N678));
nnd3s1 U288 (.Q(N766), .DIN1(N600), .DIN2(N609), .DIN3(N687));
nb1s1 U289 (.Q(N767), .DIN(N660));
nb1s1 U290 (.Q(N768), .DIN(N661));
nor2s1 U291 (.Q(N769), .DIN1(N736), .DIN2(N737));
nor2s1 U292 (.Q(N770), .DIN1(N739), .DIN2(N740));
nor2s1 U293 (.Q(N771), .DIN1(N742), .DIN2(N743));
nor2s1 U294 (.Q(N772), .DIN1(N745), .DIN2(N746));
nnd4s1 U295 (.Q(N773), .DIN1(N750), .DIN2(N762), .DIN3(N763), .DIN4(N734));
nor2s1 U296 (.Q(N777), .DIN1(N748), .DIN2(N749));
nnd3s1 U297 (.Q(N778), .DIN1(N753), .DIN2(N761), .DIN3(N733));
nor2s1 U298 (.Q(N781), .DIN1(N751), .DIN2(N752));
nnd2s1 U299 (.Q(N782), .DIN1(N756), .DIN2(N732));
nor2s1 U300 (.Q(N785), .DIN1(N754), .DIN2(N755));
nor2s1 U301 (.Q(N786), .DIN1(N757), .DIN2(N758));
nor2s1 U302 (.Q(N787), .DIN1(N759), .DIN2(N760));
nor2s1 U303 (.Q(N788), .DIN1(N700), .DIN2(N773));
and2s1 U304 (.Q(N789), .DIN1(N700), .DIN2(N773));
nor2s1 U305 (.Q(N790), .DIN1(N708), .DIN2(N778));
and2s1 U306 (.Q(N791), .DIN1(N708), .DIN2(N778));
nor2s1 U307 (.Q(N792), .DIN1(N717), .DIN2(N782));
and2s1 U308 (.Q(N793), .DIN1(N717), .DIN2(N782));
and2s1 U309 (.Q(N794), .DIN1(N219), .DIN2(N786));
nnd2s1 U310 (.Q(N795), .DIN1(N628), .DIN2(N773));
nnd2s1 U311 (.Q(N796), .DIN1(N795), .DIN2(N747));
nor2s1 U312 (.Q(N802), .DIN1(N788), .DIN2(N789));
nor2s1 U313 (.Q(N803), .DIN1(N790), .DIN2(N791));
nor2s1 U314 (.Q(N804), .DIN1(N792), .DIN2(N793));
nor2s1 U315 (.Q(N805), .DIN1(N340), .DIN2(N794));
nor2s1 U316 (.Q(N806), .DIN1(N692), .DIN2(N796));
and2s1 U317 (.Q(N807), .DIN1(N692), .DIN2(N796));
and2s1 U318 (.Q(N808), .DIN1(N219), .DIN2(N802));
and2s1 U319 (.Q(N809), .DIN1(N219), .DIN2(N803));
and2s1 U320 (.Q(N810), .DIN1(N219), .DIN2(N804));
nnd4s1 U321 (.Q(N811), .DIN1(N805), .DIN2(N787), .DIN3(N731), .DIN4(N529));
nnd2s1 U322 (.Q(N812), .DIN1(N619), .DIN2(N796));
nnd3s1 U323 (.Q(N813), .DIN1(N609), .DIN2(N619), .DIN3(N796));
nnd4s1 U324 (.Q(N814), .DIN1(N600), .DIN2(N609), .DIN3(N619), .DIN4(N796));
nnd4s1 U325 (.Q(N815), .DIN1(N738), .DIN2(N765), .DIN3(N766), .DIN4(N814));
nnd3s1 U326 (.Q(N819), .DIN1(N741), .DIN2(N764), .DIN3(N813));
nnd2s1 U327 (.Q(N822), .DIN1(N744), .DIN2(N812));
nor2s1 U328 (.Q(N825), .DIN1(N806), .DIN2(N807));
nor2s1 U329 (.Q(N826), .DIN1(N335), .DIN2(N808));
nor2s1 U330 (.Q(N827), .DIN1(N336), .DIN2(N809));
nor2s1 U331 (.Q(N828), .DIN1(N338), .DIN2(N810));
hi1s1 U332 (.Q(N829), .DIN(N811));
nor2s1 U333 (.Q(N830), .DIN1(N665), .DIN2(N815));
and2s1 U334 (.Q(N831), .DIN1(N665), .DIN2(N815));
nor2s1 U335 (.Q(N832), .DIN1(N673), .DIN2(N819));
and2s1 U336 (.Q(N833), .DIN1(N673), .DIN2(N819));
nor2s1 U337 (.Q(N834), .DIN1(N682), .DIN2(N822));
and2s1 U338 (.Q(N835), .DIN1(N682), .DIN2(N822));
and2s1 U339 (.Q(N836), .DIN1(N219), .DIN2(N825));
nnd3s1 U340 (.Q(N837), .DIN1(N826), .DIN2(N777), .DIN3(N704));
nnd4s1 U341 (.Q(N838), .DIN1(N827), .DIN2(N781), .DIN3(N712), .DIN4(N527));
nnd4s1 U342 (.Q(N839), .DIN1(N828), .DIN2(N785), .DIN3(N721), .DIN4(N528));
hi1s1 U343 (.Q(N840), .DIN(N829));
nnd2s1 U344 (.Q(N841), .DIN1(N815), .DIN2(N593));
nor2s1 U345 (.Q(N842), .DIN1(N830), .DIN2(N831));
nor2s1 U346 (.Q(N843), .DIN1(N832), .DIN2(N833));
nor2s1 U347 (.Q(N844), .DIN1(N834), .DIN2(N835));
nor2s1 U348 (.Q(N845), .DIN1(N334), .DIN2(N836));
hi1s1 U349 (.Q(N846), .DIN(N837));
hi1s1 U350 (.Q(N847), .DIN(N838));
hi1s1 U351 (.Q(N848), .DIN(N839));
and2s1 U352 (.Q(N849), .DIN1(N735), .DIN2(N841));
nb1s1 U353 (.Q(N850), .DIN(N840));
and2s1 U354 (.Q(N851), .DIN1(N219), .DIN2(N842));
and2s1 U355 (.Q(N852), .DIN1(N219), .DIN2(N843));
and2s1 U356 (.Q(N853), .DIN1(N219), .DIN2(N844));
nnd3s1 U357 (.Q(N854), .DIN1(N845), .DIN2(N772), .DIN3(N696));
hi1s1 U358 (.Q(N855), .DIN(N846));
hi1s1 U359 (.Q(N856), .DIN(N847));
hi1s1 U360 (.Q(N857), .DIN(N848));
hi1s1 U361 (.Q(N858), .DIN(N849));
nor2s1 U362 (.Q(N859), .DIN1(N417), .DIN2(N851));
nor2s1 U363 (.Q(N860), .DIN1(N332), .DIN2(N852));
nor2s1 U364 (.Q(N861), .DIN1(N333), .DIN2(N853));
hi1s1 U365 (.Q(N862), .DIN(N854));
nb1s1 U366 (.Q(N863), .DIN(N855));
nb1s1 U367 (.Q(N864), .DIN(N856));
nb1s1 U368 (.Q(N865), .DIN(N857));
nb1s1 U369 (.Q(N866), .DIN(N858));
nnd3s1 U370 (.Q(N867), .DIN1(N859), .DIN2(N769), .DIN3(N669));
nnd3s1 U371 (.Q(N868), .DIN1(N860), .DIN2(N770), .DIN3(N677));
nnd3s1 U372 (.Q(N869), .DIN1(N861), .DIN2(N771), .DIN3(N686));
hi1s1 U373 (.Q(N870), .DIN(N862));
hi1s1 U374 (.Q(N871), .DIN(N867));
hi1s1 U375 (.Q(N872), .DIN(N868));
hi1s1 U376 (.Q(N873), .DIN(N869));
nb1s1 U377 (.Q(N874), .DIN(N870));
hi1s1 U378 (.Q(N875), .DIN(N871));
hi1s1 U379 (.Q(N876), .DIN(N872));
hi1s1 U380 (.Q(N877), .DIN(N873));
nb1s1 U381 (.Q(N878), .DIN(N875));
nb1s1 U382 (.Q(N879), .DIN(N876));
nb1s1 U383 (.Q(N880), .DIN(N877));
endmodule
